`ifndef RAM_FAKE_REG_FILE_DEFINE
`define RAM_FAKE_REG_FILE_DEFINE

// temporary hardcoded values 
`define VX_MEM_BYTEEN_WIDTH     1
`define VX_MEM_ADDR_WIDTH       32
`define VX_MEM_DATA_WIDTH       32
`define VX_MEM_TAG_WIDTH        4     

`endif
