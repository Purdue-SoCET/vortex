`ifndef VORTEX_CTRL_SLAVE_DEFINE
`define VORTEX_CTRL_SLAVE_DEFINE

`define START_ADDR 32'b100001010 //read and write
`define STATUS_ADDR 32'b100001000 //read only


`endif
