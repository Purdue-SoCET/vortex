/*
    socet115 / zlagpaca@purdue.edu
    Zach Lagpacan

    module for faking memory with basic register file which can interface with Vortex memory interface
*/

`include "ram_fake_reg_file.vh"

module ram_fake_reg_file #(
    parameter WORD_W = 32
)(
    // seq
    input clk, reset,

    // Memory Request:
    // vortex outputs
    input logic                             mem_req_valid,
    input logic                             mem_req_rw,
    input logic [`VX_MEM_BYTEEN_WIDTH-1:0]  mem_req_byteen,    
    input logic [`VX_MEM_ADDR_WIDTH-1:0]    mem_req_addr,
    input logic [`VX_MEM_DATA_WIDTH-1:0]    mem_req_data,
    input logic [`VX_MEM_TAG_WIDTH-1:0]     mem_req_tag,
    // vortex inputs
    output logic                            mem_req_ready,

    // Memory response:
    // vortex inputs
    output logic                            mem_rsp_valid,        
    output logic [`VX_MEM_DATA_WIDTH-1:0]   mem_rsp_data,
    output logic [`VX_MEM_TAG_WIDTH-1:0]    mem_rsp_tag,
    // vortex outputs
    input logic                             mem_rsp_ready,

    // Status:
    // vortex outputs
    input logic                             busy,

    // tb:
    output logic                            tb_addr_out_of_bounds
);
    // register file instances
    
    // chunk 0
    logic wen_0_80000000;
    logic [9-1:0] wsel_0_80000000;
    logic [32-1:0] wdata_0_80000000;
    logic [9-1:0] rsel_0_80000000;
    logic [32-1:0] rdata_0_80000000;
    
    logic [32-1:0] reg_val_0_80000000 [512-1:0];
    logic [32-1:0] next_reg_val_0_80000000 [512-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_0_80000000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_0_80000000[0] <= 32'h6F008004;
            reg_val_0_80000000[1] <= 32'h732F2034;
            reg_val_0_80000000[2] <= 32'h930F8000;
            reg_val_0_80000000[3] <= 32'h6308FF03;
            reg_val_0_80000000[4] <= 32'h930F9000;
            reg_val_0_80000000[5] <= 32'h6304FF03;
            reg_val_0_80000000[6] <= 32'h930FB000;
            reg_val_0_80000000[7] <= 32'h6300FF03;
            reg_val_0_80000000[8] <= 32'h130F0000;
            reg_val_0_80000000[9] <= 32'h63040F00;
            reg_val_0_80000000[10] <= 32'h67000F00;
            reg_val_0_80000000[11] <= 32'h732F2034;
            reg_val_0_80000000[12] <= 32'h63540F00;
            reg_val_0_80000000[13] <= 32'h6F004000;
            reg_val_0_80000000[14] <= 32'h93E19153;
            reg_val_0_80000000[15] <= 32'h171F0000;
            reg_val_0_80000000[16] <= 32'h23223FFC;
            reg_val_0_80000000[17] <= 32'h6FF09FFF;
            reg_val_0_80000000[18] <= 32'h93000000;
            reg_val_0_80000000[19] <= 32'h13010000;
            reg_val_0_80000000[20] <= 32'h93010000;
            reg_val_0_80000000[21] <= 32'h13020000;
            reg_val_0_80000000[22] <= 32'h93020000;
            reg_val_0_80000000[23] <= 32'h13030000;
            reg_val_0_80000000[24] <= 32'h93030000;
            reg_val_0_80000000[25] <= 32'h13040000;
            reg_val_0_80000000[26] <= 32'h93040000;
            reg_val_0_80000000[27] <= 32'h13050000;
            reg_val_0_80000000[28] <= 32'h93050000;
            reg_val_0_80000000[29] <= 32'h13060000;
            reg_val_0_80000000[30] <= 32'h93060000;
            reg_val_0_80000000[31] <= 32'h13070000;
            reg_val_0_80000000[32] <= 32'h93070000;
            reg_val_0_80000000[33] <= 32'h13080000;
            reg_val_0_80000000[34] <= 32'h93080000;
            reg_val_0_80000000[35] <= 32'h13090000;
            reg_val_0_80000000[36] <= 32'h93090000;
            reg_val_0_80000000[37] <= 32'h130A0000;
            reg_val_0_80000000[38] <= 32'h930A0000;
            reg_val_0_80000000[39] <= 32'h130B0000;
            reg_val_0_80000000[40] <= 32'h930B0000;
            reg_val_0_80000000[41] <= 32'h130C0000;
            reg_val_0_80000000[42] <= 32'h930C0000;
            reg_val_0_80000000[43] <= 32'h130D0000;
            reg_val_0_80000000[44] <= 32'h930D0000;
            reg_val_0_80000000[45] <= 32'h130E0000;
            reg_val_0_80000000[46] <= 32'h930E0000;
            reg_val_0_80000000[47] <= 32'h130F0000;
            reg_val_0_80000000[48] <= 32'h930F0000;
            reg_val_0_80000000[49] <= 32'h732540F1;
            reg_val_0_80000000[50] <= 32'h63100500;
            reg_val_0_80000000[51] <= 32'h97020000;
            reg_val_0_80000000[52] <= 32'h93820201;
            reg_val_0_80000000[53] <= 32'h73905230;
            reg_val_0_80000000[54] <= 32'h73500018;
            reg_val_0_80000000[55] <= 32'h97020000;
            reg_val_0_80000000[56] <= 32'h93820202;
            reg_val_0_80000000[57] <= 32'h73905230;
            reg_val_0_80000000[58] <= 32'hB7020080;
            reg_val_0_80000000[59] <= 32'h9382F2FF;
            reg_val_0_80000000[60] <= 32'h7390023B;
            reg_val_0_80000000[61] <= 32'h9302F001;
            reg_val_0_80000000[62] <= 32'h7390023A;
            reg_val_0_80000000[63] <= 32'h73504030;
            reg_val_0_80000000[64] <= 32'h97020000;
            reg_val_0_80000000[65] <= 32'h93824201;
            reg_val_0_80000000[66] <= 32'h73905230;
            reg_val_0_80000000[67] <= 32'h73502030;
            reg_val_0_80000000[68] <= 32'h73503030;
            reg_val_0_80000000[69] <= 32'h93010000;
            reg_val_0_80000000[70] <= 32'h97020000;
            reg_val_0_80000000[71] <= 32'h9382C2EE;
            reg_val_0_80000000[72] <= 32'h73905230;
            reg_val_0_80000000[73] <= 32'h13051000;
            reg_val_0_80000000[74] <= 32'h1315F501;
            reg_val_0_80000000[75] <= 32'h634C0500;
            reg_val_0_80000000[76] <= 32'h0F00F00F;
            reg_val_0_80000000[77] <= 32'h93011000;
            reg_val_0_80000000[78] <= 32'h9308D005;
            reg_val_0_80000000[79] <= 32'h13050000;
            reg_val_0_80000000[80] <= 32'h73000000;
            reg_val_0_80000000[81] <= 32'h93020000;
            reg_val_0_80000000[82] <= 32'h638A0200;
            reg_val_0_80000000[83] <= 32'h73905210;
            reg_val_0_80000000[84] <= 32'hB7B20000;
            reg_val_0_80000000[85] <= 32'h93829210;
            reg_val_0_80000000[86] <= 32'h73902230;
            reg_val_0_80000000[87] <= 32'h73500030;
            reg_val_0_80000000[88] <= 32'h37250000;
            reg_val_0_80000000[89] <= 32'h73200530;
            reg_val_0_80000000[90] <= 32'h73503000;
            reg_val_0_80000000[91] <= 32'h97020000;
            reg_val_0_80000000[92] <= 32'h93824201;
            reg_val_0_80000000[93] <= 32'h73901234;
            reg_val_0_80000000[94] <= 32'h732540F1;
            reg_val_0_80000000[95] <= 32'h73002030;
            reg_val_0_80000000[96] <= 32'h93012000;
            reg_val_0_80000000[97] <= 32'h17250000;
            reg_val_0_80000000[98] <= 32'h1305C5E7;
            reg_val_0_80000000[99] <= 32'h07300500;
            reg_val_0_80000000[100] <= 32'h87308500;
            reg_val_0_80000000[101] <= 32'h07310501;
            reg_val_0_80000000[102] <= 32'h83268501;
            reg_val_0_80000000[103] <= 32'h0323C501;
            reg_val_0_80000000[104] <= 32'hD3711002;
            reg_val_0_80000000[105] <= 32'h27303500;
            reg_val_0_80000000[106] <= 32'h83234500;
            reg_val_0_80000000[107] <= 32'h03250500;
            reg_val_0_80000000[108] <= 32'hF3151000;
            reg_val_0_80000000[109] <= 32'h13060000;
            reg_val_0_80000000[110] <= 32'h631AD526;
            reg_val_0_80000000[111] <= 32'h63187326;
            reg_val_0_80000000[112] <= 32'h6396C526;
            reg_val_0_80000000[113] <= 32'h93013000;
            reg_val_0_80000000[114] <= 32'h17250000;
            reg_val_0_80000000[115] <= 32'h130585E5;
            reg_val_0_80000000[116] <= 32'h07300500;
            reg_val_0_80000000[117] <= 32'h87308500;
            reg_val_0_80000000[118] <= 32'h07310501;
            reg_val_0_80000000[119] <= 32'h83268501;
            reg_val_0_80000000[120] <= 32'h0323C501;
            reg_val_0_80000000[121] <= 32'hD3711002;
            reg_val_0_80000000[122] <= 32'h27303500;
            reg_val_0_80000000[123] <= 32'h83234500;
            reg_val_0_80000000[124] <= 32'h03250500;
            reg_val_0_80000000[125] <= 32'hF3151000;
            reg_val_0_80000000[126] <= 32'h13061000;
            reg_val_0_80000000[127] <= 32'h6318D522;
            reg_val_0_80000000[128] <= 32'h63167322;
            reg_val_0_80000000[129] <= 32'h6394C522;
            reg_val_0_80000000[130] <= 32'h93014000;
            reg_val_0_80000000[131] <= 32'h17250000;
            reg_val_0_80000000[132] <= 32'h130545E3;
            reg_val_0_80000000[133] <= 32'h07300500;
            reg_val_0_80000000[134] <= 32'h87308500;
            reg_val_0_80000000[135] <= 32'h07310501;
            reg_val_0_80000000[136] <= 32'h83268501;
            reg_val_0_80000000[137] <= 32'h0323C501;
            reg_val_0_80000000[138] <= 32'hD3711002;
            reg_val_0_80000000[139] <= 32'h27303500;
            reg_val_0_80000000[140] <= 32'h83234500;
            reg_val_0_80000000[141] <= 32'h03250500;
            reg_val_0_80000000[142] <= 32'hF3151000;
            reg_val_0_80000000[143] <= 32'h13061000;
            reg_val_0_80000000[144] <= 32'h6316D51E;
            reg_val_0_80000000[145] <= 32'h6314731E;
            reg_val_0_80000000[146] <= 32'h6392C51E;
            reg_val_0_80000000[147] <= 32'h93015000;
            reg_val_0_80000000[148] <= 32'h17250000;
            reg_val_0_80000000[149] <= 32'h130505E1;
            reg_val_0_80000000[150] <= 32'h07300500;
            reg_val_0_80000000[151] <= 32'h87308500;
            reg_val_0_80000000[152] <= 32'h07310501;
            reg_val_0_80000000[153] <= 32'h83268501;
            reg_val_0_80000000[154] <= 32'h0323C501;
            reg_val_0_80000000[155] <= 32'hD371100A;
            reg_val_0_80000000[156] <= 32'h27303500;
            reg_val_0_80000000[157] <= 32'h83234500;
            reg_val_0_80000000[158] <= 32'h03250500;
            reg_val_0_80000000[159] <= 32'hF3151000;
            reg_val_0_80000000[160] <= 32'h13060000;
            reg_val_0_80000000[161] <= 32'h6314D51A;
            reg_val_0_80000000[162] <= 32'h6312731A;
            reg_val_0_80000000[163] <= 32'h6390C51A;
            reg_val_0_80000000[164] <= 32'h93016000;
            reg_val_0_80000000[165] <= 32'h17250000;
            reg_val_0_80000000[166] <= 32'h1305C5DE;
            reg_val_0_80000000[167] <= 32'h07300500;
            reg_val_0_80000000[168] <= 32'h87308500;
            reg_val_0_80000000[169] <= 32'h07310501;
            reg_val_0_80000000[170] <= 32'h83268501;
            reg_val_0_80000000[171] <= 32'h0323C501;
            reg_val_0_80000000[172] <= 32'hD371100A;
            reg_val_0_80000000[173] <= 32'h27303500;
            reg_val_0_80000000[174] <= 32'h83234500;
            reg_val_0_80000000[175] <= 32'h03250500;
            reg_val_0_80000000[176] <= 32'hF3151000;
            reg_val_0_80000000[177] <= 32'h13061000;
            reg_val_0_80000000[178] <= 32'h6312D516;
            reg_val_0_80000000[179] <= 32'h63107316;
            reg_val_0_80000000[180] <= 32'h639EC514;
            reg_val_0_80000000[181] <= 32'h93017000;
            reg_val_0_80000000[182] <= 32'h17250000;
            reg_val_0_80000000[183] <= 32'h130585DC;
            reg_val_0_80000000[184] <= 32'h07300500;
            reg_val_0_80000000[185] <= 32'h87308500;
            reg_val_0_80000000[186] <= 32'h07310501;
            reg_val_0_80000000[187] <= 32'h83268501;
            reg_val_0_80000000[188] <= 32'h0323C501;
            reg_val_0_80000000[189] <= 32'hD371100A;
            reg_val_0_80000000[190] <= 32'h27303500;
            reg_val_0_80000000[191] <= 32'h83234500;
            reg_val_0_80000000[192] <= 32'h03250500;
            reg_val_0_80000000[193] <= 32'hF3151000;
            reg_val_0_80000000[194] <= 32'h13061000;
            reg_val_0_80000000[195] <= 32'h6310D512;
            reg_val_0_80000000[196] <= 32'h631E7310;
            reg_val_0_80000000[197] <= 32'h639CC510;
            reg_val_0_80000000[198] <= 32'h93018000;
            reg_val_0_80000000[199] <= 32'h17250000;
            reg_val_0_80000000[200] <= 32'h130545DA;
            reg_val_0_80000000[201] <= 32'h07300500;
            reg_val_0_80000000[202] <= 32'h87308500;
            reg_val_0_80000000[203] <= 32'h07310501;
            reg_val_0_80000000[204] <= 32'h83268501;
            reg_val_0_80000000[205] <= 32'h0323C501;
            reg_val_0_80000000[206] <= 32'hD3711012;
            reg_val_0_80000000[207] <= 32'h27303500;
            reg_val_0_80000000[208] <= 32'h83234500;
            reg_val_0_80000000[209] <= 32'h03250500;
            reg_val_0_80000000[210] <= 32'hF3151000;
            reg_val_0_80000000[211] <= 32'h13060000;
            reg_val_0_80000000[212] <= 32'h631ED50C;
            reg_val_0_80000000[213] <= 32'h631C730C;
            reg_val_0_80000000[214] <= 32'h639AC50C;
            reg_val_0_80000000[215] <= 32'h93019000;
            reg_val_0_80000000[216] <= 32'h17250000;
            reg_val_0_80000000[217] <= 32'h130505D8;
            reg_val_0_80000000[218] <= 32'h07300500;
            reg_val_0_80000000[219] <= 32'h87308500;
            reg_val_0_80000000[220] <= 32'h07310501;
            reg_val_0_80000000[221] <= 32'h83268501;
            reg_val_0_80000000[222] <= 32'h0323C501;
            reg_val_0_80000000[223] <= 32'hD3711012;
            reg_val_0_80000000[224] <= 32'h27303500;
            reg_val_0_80000000[225] <= 32'h83234500;
            reg_val_0_80000000[226] <= 32'h03250500;
            reg_val_0_80000000[227] <= 32'hF3151000;
            reg_val_0_80000000[228] <= 32'h13061000;
            reg_val_0_80000000[229] <= 32'h631CD508;
            reg_val_0_80000000[230] <= 32'h631A7308;
            reg_val_0_80000000[231] <= 32'h6398C508;
            reg_val_0_80000000[232] <= 32'h9301A000;
            reg_val_0_80000000[233] <= 32'h17250000;
            reg_val_0_80000000[234] <= 32'h1305C5D5;
            reg_val_0_80000000[235] <= 32'h07300500;
            reg_val_0_80000000[236] <= 32'h87308500;
            reg_val_0_80000000[237] <= 32'h07310501;
            reg_val_0_80000000[238] <= 32'h83268501;
            reg_val_0_80000000[239] <= 32'h0323C501;
            reg_val_0_80000000[240] <= 32'hD3711012;
            reg_val_0_80000000[241] <= 32'h27303500;
            reg_val_0_80000000[242] <= 32'h83234500;
            reg_val_0_80000000[243] <= 32'h03250500;
            reg_val_0_80000000[244] <= 32'hF3151000;
            reg_val_0_80000000[245] <= 32'h13061000;
            reg_val_0_80000000[246] <= 32'h631AD504;
            reg_val_0_80000000[247] <= 32'h63187304;
            reg_val_0_80000000[248] <= 32'h6396C504;
            reg_val_0_80000000[249] <= 32'h9301B000;
            reg_val_0_80000000[250] <= 32'h17250000;
            reg_val_0_80000000[251] <= 32'h130585D3;
            reg_val_0_80000000[252] <= 32'h07300500;
            reg_val_0_80000000[253] <= 32'h87308500;
            reg_val_0_80000000[254] <= 32'h07310501;
            reg_val_0_80000000[255] <= 32'h83268501;
            reg_val_0_80000000[256] <= 32'h0323C501;
            reg_val_0_80000000[257] <= 32'hD371100A;
            reg_val_0_80000000[258] <= 32'h27303500;
            reg_val_0_80000000[259] <= 32'h83234500;
            reg_val_0_80000000[260] <= 32'h03250500;
            reg_val_0_80000000[261] <= 32'hF3151000;
            reg_val_0_80000000[262] <= 32'h13060001;
            reg_val_0_80000000[263] <= 32'h6318D500;
            reg_val_0_80000000[264] <= 32'h63167300;
            reg_val_0_80000000[265] <= 32'h6394C500;
            reg_val_0_80000000[266] <= 32'h63103002;
            reg_val_0_80000000[267] <= 32'h0F00F00F;
            reg_val_0_80000000[268] <= 32'h63800100;
            reg_val_0_80000000[269] <= 32'h93911100;
            reg_val_0_80000000[270] <= 32'h93E11100;
            reg_val_0_80000000[271] <= 32'h9308D005;
            reg_val_0_80000000[272] <= 32'h13850100;
            reg_val_0_80000000[273] <= 32'h73000000;
            reg_val_0_80000000[274] <= 32'h0F00F00F;
            reg_val_0_80000000[275] <= 32'h93011000;
            reg_val_0_80000000[276] <= 32'h9308D005;
            reg_val_0_80000000[277] <= 32'h13050000;
            reg_val_0_80000000[278] <= 32'h73000000;
            reg_val_0_80000000[279] <= 32'h731000C0;
            reg_val_0_80000000[280] <= 32'h00000000;
            reg_val_0_80000000[281] <= 32'h00000000;
            reg_val_0_80000000[282] <= 32'h00000000;
            reg_val_0_80000000[283] <= 32'h00000000;
            reg_val_0_80000000[284] <= 32'h00000000;
            reg_val_0_80000000[285] <= 32'h00000000;
            reg_val_0_80000000[286] <= 32'h00000000;
            // fill-in reset values:
            reg_val_0_80000000[287] <= 32'h00000000;
            reg_val_0_80000000[288] <= 32'h00000000;
            reg_val_0_80000000[289] <= 32'h00000000;
            reg_val_0_80000000[290] <= 32'h00000000;
            reg_val_0_80000000[291] <= 32'h00000000;
            reg_val_0_80000000[292] <= 32'h00000000;
            reg_val_0_80000000[293] <= 32'h00000000;
            reg_val_0_80000000[294] <= 32'h00000000;
            reg_val_0_80000000[295] <= 32'h00000000;
            reg_val_0_80000000[296] <= 32'h00000000;
            reg_val_0_80000000[297] <= 32'h00000000;
            reg_val_0_80000000[298] <= 32'h00000000;
            reg_val_0_80000000[299] <= 32'h00000000;
            reg_val_0_80000000[300] <= 32'h00000000;
            reg_val_0_80000000[301] <= 32'h00000000;
            reg_val_0_80000000[302] <= 32'h00000000;
            reg_val_0_80000000[303] <= 32'h00000000;
            reg_val_0_80000000[304] <= 32'h00000000;
            reg_val_0_80000000[305] <= 32'h00000000;
            reg_val_0_80000000[306] <= 32'h00000000;
            reg_val_0_80000000[307] <= 32'h00000000;
            reg_val_0_80000000[308] <= 32'h00000000;
            reg_val_0_80000000[309] <= 32'h00000000;
            reg_val_0_80000000[310] <= 32'h00000000;
            reg_val_0_80000000[311] <= 32'h00000000;
            reg_val_0_80000000[312] <= 32'h00000000;
            reg_val_0_80000000[313] <= 32'h00000000;
            reg_val_0_80000000[314] <= 32'h00000000;
            reg_val_0_80000000[315] <= 32'h00000000;
            reg_val_0_80000000[316] <= 32'h00000000;
            reg_val_0_80000000[317] <= 32'h00000000;
            reg_val_0_80000000[318] <= 32'h00000000;
            reg_val_0_80000000[319] <= 32'h00000000;
            reg_val_0_80000000[320] <= 32'h00000000;
            reg_val_0_80000000[321] <= 32'h00000000;
            reg_val_0_80000000[322] <= 32'h00000000;
            reg_val_0_80000000[323] <= 32'h00000000;
            reg_val_0_80000000[324] <= 32'h00000000;
            reg_val_0_80000000[325] <= 32'h00000000;
            reg_val_0_80000000[326] <= 32'h00000000;
            reg_val_0_80000000[327] <= 32'h00000000;
            reg_val_0_80000000[328] <= 32'h00000000;
            reg_val_0_80000000[329] <= 32'h00000000;
            reg_val_0_80000000[330] <= 32'h00000000;
            reg_val_0_80000000[331] <= 32'h00000000;
            reg_val_0_80000000[332] <= 32'h00000000;
            reg_val_0_80000000[333] <= 32'h00000000;
            reg_val_0_80000000[334] <= 32'h00000000;
            reg_val_0_80000000[335] <= 32'h00000000;
            reg_val_0_80000000[336] <= 32'h00000000;
            reg_val_0_80000000[337] <= 32'h00000000;
            reg_val_0_80000000[338] <= 32'h00000000;
            reg_val_0_80000000[339] <= 32'h00000000;
            reg_val_0_80000000[340] <= 32'h00000000;
            reg_val_0_80000000[341] <= 32'h00000000;
            reg_val_0_80000000[342] <= 32'h00000000;
            reg_val_0_80000000[343] <= 32'h00000000;
            reg_val_0_80000000[344] <= 32'h00000000;
            reg_val_0_80000000[345] <= 32'h00000000;
            reg_val_0_80000000[346] <= 32'h00000000;
            reg_val_0_80000000[347] <= 32'h00000000;
            reg_val_0_80000000[348] <= 32'h00000000;
            reg_val_0_80000000[349] <= 32'h00000000;
            reg_val_0_80000000[350] <= 32'h00000000;
            reg_val_0_80000000[351] <= 32'h00000000;
            reg_val_0_80000000[352] <= 32'h00000000;
            reg_val_0_80000000[353] <= 32'h00000000;
            reg_val_0_80000000[354] <= 32'h00000000;
            reg_val_0_80000000[355] <= 32'h00000000;
            reg_val_0_80000000[356] <= 32'h00000000;
            reg_val_0_80000000[357] <= 32'h00000000;
            reg_val_0_80000000[358] <= 32'h00000000;
            reg_val_0_80000000[359] <= 32'h00000000;
            reg_val_0_80000000[360] <= 32'h00000000;
            reg_val_0_80000000[361] <= 32'h00000000;
            reg_val_0_80000000[362] <= 32'h00000000;
            reg_val_0_80000000[363] <= 32'h00000000;
            reg_val_0_80000000[364] <= 32'h00000000;
            reg_val_0_80000000[365] <= 32'h00000000;
            reg_val_0_80000000[366] <= 32'h00000000;
            reg_val_0_80000000[367] <= 32'h00000000;
            reg_val_0_80000000[368] <= 32'h00000000;
            reg_val_0_80000000[369] <= 32'h00000000;
            reg_val_0_80000000[370] <= 32'h00000000;
            reg_val_0_80000000[371] <= 32'h00000000;
            reg_val_0_80000000[372] <= 32'h00000000;
            reg_val_0_80000000[373] <= 32'h00000000;
            reg_val_0_80000000[374] <= 32'h00000000;
            reg_val_0_80000000[375] <= 32'h00000000;
            reg_val_0_80000000[376] <= 32'h00000000;
            reg_val_0_80000000[377] <= 32'h00000000;
            reg_val_0_80000000[378] <= 32'h00000000;
            reg_val_0_80000000[379] <= 32'h00000000;
            reg_val_0_80000000[380] <= 32'h00000000;
            reg_val_0_80000000[381] <= 32'h00000000;
            reg_val_0_80000000[382] <= 32'h00000000;
            reg_val_0_80000000[383] <= 32'h00000000;
            reg_val_0_80000000[384] <= 32'h00000000;
            reg_val_0_80000000[385] <= 32'h00000000;
            reg_val_0_80000000[386] <= 32'h00000000;
            reg_val_0_80000000[387] <= 32'h00000000;
            reg_val_0_80000000[388] <= 32'h00000000;
            reg_val_0_80000000[389] <= 32'h00000000;
            reg_val_0_80000000[390] <= 32'h00000000;
            reg_val_0_80000000[391] <= 32'h00000000;
            reg_val_0_80000000[392] <= 32'h00000000;
            reg_val_0_80000000[393] <= 32'h00000000;
            reg_val_0_80000000[394] <= 32'h00000000;
            reg_val_0_80000000[395] <= 32'h00000000;
            reg_val_0_80000000[396] <= 32'h00000000;
            reg_val_0_80000000[397] <= 32'h00000000;
            reg_val_0_80000000[398] <= 32'h00000000;
            reg_val_0_80000000[399] <= 32'h00000000;
            reg_val_0_80000000[400] <= 32'h00000000;
            reg_val_0_80000000[401] <= 32'h00000000;
            reg_val_0_80000000[402] <= 32'h00000000;
            reg_val_0_80000000[403] <= 32'h00000000;
            reg_val_0_80000000[404] <= 32'h00000000;
            reg_val_0_80000000[405] <= 32'h00000000;
            reg_val_0_80000000[406] <= 32'h00000000;
            reg_val_0_80000000[407] <= 32'h00000000;
            reg_val_0_80000000[408] <= 32'h00000000;
            reg_val_0_80000000[409] <= 32'h00000000;
            reg_val_0_80000000[410] <= 32'h00000000;
            reg_val_0_80000000[411] <= 32'h00000000;
            reg_val_0_80000000[412] <= 32'h00000000;
            reg_val_0_80000000[413] <= 32'h00000000;
            reg_val_0_80000000[414] <= 32'h00000000;
            reg_val_0_80000000[415] <= 32'h00000000;
            reg_val_0_80000000[416] <= 32'h00000000;
            reg_val_0_80000000[417] <= 32'h00000000;
            reg_val_0_80000000[418] <= 32'h00000000;
            reg_val_0_80000000[419] <= 32'h00000000;
            reg_val_0_80000000[420] <= 32'h00000000;
            reg_val_0_80000000[421] <= 32'h00000000;
            reg_val_0_80000000[422] <= 32'h00000000;
            reg_val_0_80000000[423] <= 32'h00000000;
            reg_val_0_80000000[424] <= 32'h00000000;
            reg_val_0_80000000[425] <= 32'h00000000;
            reg_val_0_80000000[426] <= 32'h00000000;
            reg_val_0_80000000[427] <= 32'h00000000;
            reg_val_0_80000000[428] <= 32'h00000000;
            reg_val_0_80000000[429] <= 32'h00000000;
            reg_val_0_80000000[430] <= 32'h00000000;
            reg_val_0_80000000[431] <= 32'h00000000;
            reg_val_0_80000000[432] <= 32'h00000000;
            reg_val_0_80000000[433] <= 32'h00000000;
            reg_val_0_80000000[434] <= 32'h00000000;
            reg_val_0_80000000[435] <= 32'h00000000;
            reg_val_0_80000000[436] <= 32'h00000000;
            reg_val_0_80000000[437] <= 32'h00000000;
            reg_val_0_80000000[438] <= 32'h00000000;
            reg_val_0_80000000[439] <= 32'h00000000;
            reg_val_0_80000000[440] <= 32'h00000000;
            reg_val_0_80000000[441] <= 32'h00000000;
            reg_val_0_80000000[442] <= 32'h00000000;
            reg_val_0_80000000[443] <= 32'h00000000;
            reg_val_0_80000000[444] <= 32'h00000000;
            reg_val_0_80000000[445] <= 32'h00000000;
            reg_val_0_80000000[446] <= 32'h00000000;
            reg_val_0_80000000[447] <= 32'h00000000;
            reg_val_0_80000000[448] <= 32'h00000000;
            reg_val_0_80000000[449] <= 32'h00000000;
            reg_val_0_80000000[450] <= 32'h00000000;
            reg_val_0_80000000[451] <= 32'h00000000;
            reg_val_0_80000000[452] <= 32'h00000000;
            reg_val_0_80000000[453] <= 32'h00000000;
            reg_val_0_80000000[454] <= 32'h00000000;
            reg_val_0_80000000[455] <= 32'h00000000;
            reg_val_0_80000000[456] <= 32'h00000000;
            reg_val_0_80000000[457] <= 32'h00000000;
            reg_val_0_80000000[458] <= 32'h00000000;
            reg_val_0_80000000[459] <= 32'h00000000;
            reg_val_0_80000000[460] <= 32'h00000000;
            reg_val_0_80000000[461] <= 32'h00000000;
            reg_val_0_80000000[462] <= 32'h00000000;
            reg_val_0_80000000[463] <= 32'h00000000;
            reg_val_0_80000000[464] <= 32'h00000000;
            reg_val_0_80000000[465] <= 32'h00000000;
            reg_val_0_80000000[466] <= 32'h00000000;
            reg_val_0_80000000[467] <= 32'h00000000;
            reg_val_0_80000000[468] <= 32'h00000000;
            reg_val_0_80000000[469] <= 32'h00000000;
            reg_val_0_80000000[470] <= 32'h00000000;
            reg_val_0_80000000[471] <= 32'h00000000;
            reg_val_0_80000000[472] <= 32'h00000000;
            reg_val_0_80000000[473] <= 32'h00000000;
            reg_val_0_80000000[474] <= 32'h00000000;
            reg_val_0_80000000[475] <= 32'h00000000;
            reg_val_0_80000000[476] <= 32'h00000000;
            reg_val_0_80000000[477] <= 32'h00000000;
            reg_val_0_80000000[478] <= 32'h00000000;
            reg_val_0_80000000[479] <= 32'h00000000;
            reg_val_0_80000000[480] <= 32'h00000000;
            reg_val_0_80000000[481] <= 32'h00000000;
            reg_val_0_80000000[482] <= 32'h00000000;
            reg_val_0_80000000[483] <= 32'h00000000;
            reg_val_0_80000000[484] <= 32'h00000000;
            reg_val_0_80000000[485] <= 32'h00000000;
            reg_val_0_80000000[486] <= 32'h00000000;
            reg_val_0_80000000[487] <= 32'h00000000;
            reg_val_0_80000000[488] <= 32'h00000000;
            reg_val_0_80000000[489] <= 32'h00000000;
            reg_val_0_80000000[490] <= 32'h00000000;
            reg_val_0_80000000[491] <= 32'h00000000;
            reg_val_0_80000000[492] <= 32'h00000000;
            reg_val_0_80000000[493] <= 32'h00000000;
            reg_val_0_80000000[494] <= 32'h00000000;
            reg_val_0_80000000[495] <= 32'h00000000;
            reg_val_0_80000000[496] <= 32'h00000000;
            reg_val_0_80000000[497] <= 32'h00000000;
            reg_val_0_80000000[498] <= 32'h00000000;
            reg_val_0_80000000[499] <= 32'h00000000;
            reg_val_0_80000000[500] <= 32'h00000000;
            reg_val_0_80000000[501] <= 32'h00000000;
            reg_val_0_80000000[502] <= 32'h00000000;
            reg_val_0_80000000[503] <= 32'h00000000;
            reg_val_0_80000000[504] <= 32'h00000000;
            reg_val_0_80000000[505] <= 32'h00000000;
            reg_val_0_80000000[506] <= 32'h00000000;
            reg_val_0_80000000[507] <= 32'h00000000;
            reg_val_0_80000000[508] <= 32'h00000000;
            reg_val_0_80000000[509] <= 32'h00000000;
            reg_val_0_80000000[510] <= 32'h00000000;
            reg_val_0_80000000[511] <= 32'h00000000;
        end
        else
        begin
            reg_val_0_80000000 = next_reg_val_0_80000000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_0_80000000
        // hold reg val by default
        for (int i = 0; i < 512; i++)
        begin
            next_reg_val_0_80000000[i] = reg_val_0_80000000[i];
        end
        // update reg val if wen
        if (wen_0_80000000)
        begin
            next_reg_val_0_80000000[wsel_0_80000000] = wdata_0_80000000;
        end
    end
    
    always_comb begin : READ_LOGIC_0_80000000
        // read val at rsel
        rdata_0_80000000 = reg_val_0_80000000[rsel_0_80000000];
    end
    
    // chunk 1
    logic wen_1_80001000;
    logic [5-1:0] wsel_1_80001000;
    logic [32-1:0] wdata_1_80001000;
    logic [5-1:0] rsel_1_80001000;
    logic [32-1:0] rdata_1_80001000;
    
    logic [32-1:0] reg_val_1_80001000 [32-1:0];
    logic [32-1:0] next_reg_val_1_80001000 [32-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_1_80001000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_1_80001000[0] <= 32'h00000000;
            reg_val_1_80001000[1] <= 32'h00000000;
            reg_val_1_80001000[2] <= 32'h00000000;
            reg_val_1_80001000[3] <= 32'h00000000;
            reg_val_1_80001000[4] <= 32'h00000000;
            reg_val_1_80001000[5] <= 32'h00000000;
            reg_val_1_80001000[6] <= 32'h00000000;
            reg_val_1_80001000[7] <= 32'h00000000;
            reg_val_1_80001000[8] <= 32'h00000000;
            reg_val_1_80001000[9] <= 32'h00000000;
            reg_val_1_80001000[10] <= 32'h00000000;
            reg_val_1_80001000[11] <= 32'h00000000;
            reg_val_1_80001000[12] <= 32'h00000000;
            reg_val_1_80001000[13] <= 32'h00000000;
            reg_val_1_80001000[14] <= 32'h00000000;
            reg_val_1_80001000[15] <= 32'h00000000;
            reg_val_1_80001000[16] <= 32'h00000000;
            reg_val_1_80001000[17] <= 32'h00000000;
            // fill-in reset values:
            reg_val_1_80001000[18] <= 32'h00000000;
            reg_val_1_80001000[19] <= 32'h00000000;
            reg_val_1_80001000[20] <= 32'h00000000;
            reg_val_1_80001000[21] <= 32'h00000000;
            reg_val_1_80001000[22] <= 32'h00000000;
            reg_val_1_80001000[23] <= 32'h00000000;
            reg_val_1_80001000[24] <= 32'h00000000;
            reg_val_1_80001000[25] <= 32'h00000000;
            reg_val_1_80001000[26] <= 32'h00000000;
            reg_val_1_80001000[27] <= 32'h00000000;
            reg_val_1_80001000[28] <= 32'h00000000;
            reg_val_1_80001000[29] <= 32'h00000000;
            reg_val_1_80001000[30] <= 32'h00000000;
            reg_val_1_80001000[31] <= 32'h00000000;
        end
        else
        begin
            reg_val_1_80001000 = next_reg_val_1_80001000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_1_80001000
        // hold reg val by default
        for (int i = 0; i < 32; i++)
        begin
            next_reg_val_1_80001000[i] = reg_val_1_80001000[i];
        end
        // update reg val if wen
        if (wen_1_80001000)
        begin
            next_reg_val_1_80001000[wsel_1_80001000] = wdata_1_80001000;
        end
    end
    
    always_comb begin : READ_LOGIC_1_80001000
        // read val at rsel
        rdata_1_80001000 = reg_val_1_80001000[rsel_1_80001000];
    end
    
    // chunk 2
    logic wen_2_80002000;
    logic [7-1:0] wsel_2_80002000;
    logic [32-1:0] wdata_2_80002000;
    logic [7-1:0] rsel_2_80002000;
    logic [32-1:0] rdata_2_80002000;
    
    logic [32-1:0] reg_val_2_80002000 [128-1:0];
    logic [32-1:0] next_reg_val_2_80002000 [128-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_2_80002000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_2_80002000[0] <= 32'h00000000;
            reg_val_2_80002000[1] <= 32'h00000440;
            reg_val_2_80002000[2] <= 32'h00000000;
            reg_val_2_80002000[3] <= 32'h0000F03F;
            reg_val_2_80002000[4] <= 32'h00000000;
            reg_val_2_80002000[5] <= 32'h00000000;
            reg_val_2_80002000[6] <= 32'h00000000;
            reg_val_2_80002000[7] <= 32'h00000C40;
            reg_val_2_80002000[8] <= 32'h66666666;
            reg_val_2_80002000[9] <= 32'h664C93C0;
            reg_val_2_80002000[10] <= 32'h9A999999;
            reg_val_2_80002000[11] <= 32'h9999F13F;
            reg_val_2_80002000[12] <= 32'h00000000;
            reg_val_2_80002000[13] <= 32'h00000000;
            reg_val_2_80002000[14] <= 32'h00000000;
            reg_val_2_80002000[15] <= 32'h004893C0;
            reg_val_2_80002000[16] <= 32'hF1D4C853;
            reg_val_2_80002000[17] <= 32'hFB210940;
            reg_val_2_80002000[18] <= 32'h3A8C30E2;
            reg_val_2_80002000[19] <= 32'h8E79453E;
            reg_val_2_80002000[20] <= 32'h00000000;
            reg_val_2_80002000[21] <= 32'h00000000;
            reg_val_2_80002000[22] <= 32'hDF6D2055;
            reg_val_2_80002000[23] <= 32'hFB210940;
            reg_val_2_80002000[24] <= 32'h00000000;
            reg_val_2_80002000[25] <= 32'h00000440;
            reg_val_2_80002000[26] <= 32'h00000000;
            reg_val_2_80002000[27] <= 32'h0000F03F;
            reg_val_2_80002000[28] <= 32'h00000000;
            reg_val_2_80002000[29] <= 32'h00000000;
            reg_val_2_80002000[30] <= 32'h00000000;
            reg_val_2_80002000[31] <= 32'h0000F83F;
            reg_val_2_80002000[32] <= 32'h66666666;
            reg_val_2_80002000[33] <= 32'h664C93C0;
            reg_val_2_80002000[34] <= 32'h9A999999;
            reg_val_2_80002000[35] <= 32'h9999F1BF;
            reg_val_2_80002000[36] <= 32'h00000000;
            reg_val_2_80002000[37] <= 32'h00000000;
            reg_val_2_80002000[38] <= 32'h00000000;
            reg_val_2_80002000[39] <= 32'h004893C0;
            reg_val_2_80002000[40] <= 32'hF1D4C853;
            reg_val_2_80002000[41] <= 32'hFB210940;
            reg_val_2_80002000[42] <= 32'h3A8C30E2;
            reg_val_2_80002000[43] <= 32'h8E79453E;
            reg_val_2_80002000[44] <= 32'h00000000;
            reg_val_2_80002000[45] <= 32'h00000000;
            reg_val_2_80002000[46] <= 32'h033C7152;
            reg_val_2_80002000[47] <= 32'hFB210940;
            reg_val_2_80002000[48] <= 32'h00000000;
            reg_val_2_80002000[49] <= 32'h00000440;
            reg_val_2_80002000[50] <= 32'h00000000;
            reg_val_2_80002000[51] <= 32'h0000F03F;
            reg_val_2_80002000[52] <= 32'h00000000;
            reg_val_2_80002000[53] <= 32'h00000000;
            reg_val_2_80002000[54] <= 32'h00000000;
            reg_val_2_80002000[55] <= 32'h00000440;
            reg_val_2_80002000[56] <= 32'h66666666;
            reg_val_2_80002000[57] <= 32'h664C93C0;
            reg_val_2_80002000[58] <= 32'h9A999999;
            reg_val_2_80002000[59] <= 32'h9999F1BF;
            reg_val_2_80002000[60] <= 32'h00000000;
            reg_val_2_80002000[61] <= 32'h00000000;
            reg_val_2_80002000[62] <= 32'h3D0AD7A3;
            reg_val_2_80002000[63] <= 32'h703A9540;
            reg_val_2_80002000[64] <= 32'hF1D4C853;
            reg_val_2_80002000[65] <= 32'hFB210940;
            reg_val_2_80002000[66] <= 32'h3A8C30E2;
            reg_val_2_80002000[67] <= 32'h8E79453E;
            reg_val_2_80002000[68] <= 32'h00000000;
            reg_val_2_80002000[69] <= 32'h00000000;
            reg_val_2_80002000[70] <= 32'h09FFC1A5;
            reg_val_2_80002000[71] <= 32'hC5DD603E;
            reg_val_2_80002000[72] <= 32'h00000000;
            reg_val_2_80002000[73] <= 32'h0000F07F;
            reg_val_2_80002000[74] <= 32'h00000000;
            reg_val_2_80002000[75] <= 32'h0000F07F;
            reg_val_2_80002000[76] <= 32'h00000000;
            reg_val_2_80002000[77] <= 32'h00000000;
            reg_val_2_80002000[78] <= 32'h00000000;
            reg_val_2_80002000[79] <= 32'h0000F87F;
            // fill-in reset values:
            reg_val_2_80002000[80] <= 32'h00000000;
            reg_val_2_80002000[81] <= 32'h00000000;
            reg_val_2_80002000[82] <= 32'h00000000;
            reg_val_2_80002000[83] <= 32'h00000000;
            reg_val_2_80002000[84] <= 32'h00000000;
            reg_val_2_80002000[85] <= 32'h00000000;
            reg_val_2_80002000[86] <= 32'h00000000;
            reg_val_2_80002000[87] <= 32'h00000000;
            reg_val_2_80002000[88] <= 32'h00000000;
            reg_val_2_80002000[89] <= 32'h00000000;
            reg_val_2_80002000[90] <= 32'h00000000;
            reg_val_2_80002000[91] <= 32'h00000000;
            reg_val_2_80002000[92] <= 32'h00000000;
            reg_val_2_80002000[93] <= 32'h00000000;
            reg_val_2_80002000[94] <= 32'h00000000;
            reg_val_2_80002000[95] <= 32'h00000000;
            reg_val_2_80002000[96] <= 32'h00000000;
            reg_val_2_80002000[97] <= 32'h00000000;
            reg_val_2_80002000[98] <= 32'h00000000;
            reg_val_2_80002000[99] <= 32'h00000000;
            reg_val_2_80002000[100] <= 32'h00000000;
            reg_val_2_80002000[101] <= 32'h00000000;
            reg_val_2_80002000[102] <= 32'h00000000;
            reg_val_2_80002000[103] <= 32'h00000000;
            reg_val_2_80002000[104] <= 32'h00000000;
            reg_val_2_80002000[105] <= 32'h00000000;
            reg_val_2_80002000[106] <= 32'h00000000;
            reg_val_2_80002000[107] <= 32'h00000000;
            reg_val_2_80002000[108] <= 32'h00000000;
            reg_val_2_80002000[109] <= 32'h00000000;
            reg_val_2_80002000[110] <= 32'h00000000;
            reg_val_2_80002000[111] <= 32'h00000000;
            reg_val_2_80002000[112] <= 32'h00000000;
            reg_val_2_80002000[113] <= 32'h00000000;
            reg_val_2_80002000[114] <= 32'h00000000;
            reg_val_2_80002000[115] <= 32'h00000000;
            reg_val_2_80002000[116] <= 32'h00000000;
            reg_val_2_80002000[117] <= 32'h00000000;
            reg_val_2_80002000[118] <= 32'h00000000;
            reg_val_2_80002000[119] <= 32'h00000000;
            reg_val_2_80002000[120] <= 32'h00000000;
            reg_val_2_80002000[121] <= 32'h00000000;
            reg_val_2_80002000[122] <= 32'h00000000;
            reg_val_2_80002000[123] <= 32'h00000000;
            reg_val_2_80002000[124] <= 32'h00000000;
            reg_val_2_80002000[125] <= 32'h00000000;
            reg_val_2_80002000[126] <= 32'h00000000;
            reg_val_2_80002000[127] <= 32'h00000000;
        end
        else
        begin
            reg_val_2_80002000 = next_reg_val_2_80002000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_2_80002000
        // hold reg val by default
        for (int i = 0; i < 128; i++)
        begin
            next_reg_val_2_80002000[i] = reg_val_2_80002000[i];
        end
        // update reg val if wen
        if (wen_2_80002000)
        begin
            next_reg_val_2_80002000[wsel_2_80002000] = wdata_2_80002000;
        end
    end
    
    always_comb begin : READ_LOGIC_2_80002000
        // read val at rsel
        rdata_2_80002000 = reg_val_2_80002000[rsel_2_80002000];
    end
    
    // need reg file/chunk selection signal
    logic [2-1:0] chunk_sel;

    // addr hashing logic
    always_comb begin : ADDR_HASHING_LOGIC
        
        // bad address assertion:
        assert (
            (32'h80000000 <= mem_req_addr && mem_req_addr <= 32'h8000011f) ||
            (32'h80001000 <= mem_req_addr && mem_req_addr <= 32'h80001012) ||
            (32'h80002000 <= mem_req_addr && mem_req_addr <= 32'h80002050)
        ) else begin
            $display("mem request at address not available in chunk");
        end
        
        // bit = 1 branch
        if (mem_req_addr[WORD_W - 19] == 1'b1)
        begin
            // select chunk @ 0x80002000
            chunk_sel = 2;
        end
        // bit = 0 branch
        else if (mem_req_addr[WORD_W - 19] == 1'b0)
        begin
            if (mem_req_addr[WORD_W - 20] == 1'b0)
            begin
                // select chunk @ 0x80000000
                chunk_sel = 0;
            end
            else if (mem_req_addr[WORD_W - 20] == 1'b1)
            begin
                // select chunk @ 0x80001000
                chunk_sel = 1;
            end
        end
        else
        begin
            $display("error: got to else in high-level branch");
        end
        
        // hardwired outputs:
        // hardwiring for chunk 0
        wsel_0_80000000 = mem_req_addr[9-1 +2 : 0 +2];
        wdata_0_80000000 = mem_req_data[9-1 +2 : 0 +2];
        rsel_0_80000000 = mem_req_addr[9-1 +2 : 0 +2];
        // hardwiring for chunk 1
        wsel_1_80001000 = mem_req_addr[5-1 +2 : 0 +2];
        wdata_1_80001000 = mem_req_data[5-1 +2 : 0 +2];
        rsel_1_80001000 = mem_req_addr[5-1 +2 : 0 +2];
        // hardwiring for chunk 2
        wsel_2_80002000 = mem_req_addr[7-1 +2 : 0 +2];
        wdata_2_80002000 = mem_req_data[7-1 +2 : 0 +2];
        rsel_2_80002000 = mem_req_addr[7-1 +2 : 0 +2];
        
        // default outputs:
        mem_rsp_data = '0;
        tb_addr_out_of_bounds = 1'b0;
        // chunk wen's:
        wen_0_80000000 = 1'b0;
        wen_1_80001000 = 1'b0;
        wen_2_80002000 = 1'b0;
        
        // case for routing to diff reg file chunks
        casez (chunk_sel)
        
            // select chunk 0 @ 0x80000000
            0:
            begin
                // write routing
                wen_0_80000000 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_0_80000000;
            end
        
            // select chunk 1 @ 0x80001000
            1:
            begin
                // write routing
                wen_1_80001000 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_1_80001000;
            end
        
            // select chunk 2 @ 0x80002000
            2:
            begin
                // write routing
                wen_2_80002000 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_2_80002000;
            end
        
            // shouldn't get here
            default:
            begin
                mem_rsp_data = '0;
                tb_addr_out_of_bounds = 1'b1;
            end
        endcase
    end

    // other combinational logic for memory interface
    always_comb begin : OTHER_MEM_COMB_LOGIC

        mem_req_ready = 1'b1;           // always ready for request
        mem_rsp_valid = mem_req_valid;  // read ready immediately
        mem_rsp_tag = mem_req_tag;      // match req immediately
    end

    // NOTES:
    // don't know what to do with: 
        // mem_req_byteeen
        // busy

endmodule
