/*
    socet115 / zlagpaca@purdue.edu
    Zach Lagpacan

    module for on-chip RAM fake register file with AFTx07 AHB slave interface (at generic bus interface) 
    and Vortex memory interface 

    assumptions:
        AHB only references word addresses
*/

//////////////////////////////////////
// LOADED IN "hex_files/double.hex" //
//////////////////////////////////////

// temporary include to have defined vals
`include "Vortex_mem_slave.vh"

// include for Vortex widths
`include "../include/VX_define.vh"

module Vortex_mem_slave #(
    /////////////////
    // parameters: //
    /////////////////

    // parameter VORTEX_START_PC_ADDR = 32'h80000000,
    parameter VORTEX_MEM_SLAVE_AHB_BASE_ADDR = 32'hF000_0000,
    // parameter LOCAL_MEM_SIZE = 12
	parameter LOCAL_MEM_SIZE = 15
)(
    /////////////////
    // Sequential: //
    /////////////////
    input clk, nRST,

    ///////////////////////
    // Memory Interface: //
    ///////////////////////

    // Memory Request:
    // vortex outputs
    input logic                             mem_req_valid,
    input logic                             mem_req_rw,
    input logic [`VX_MEM_BYTEEN_WIDTH-1:0]  mem_req_byteen, // 64 (512 / 8)
    input logic [`VX_MEM_ADDR_WIDTH-1:0]    mem_req_addr,   // 26
    input logic [`VX_MEM_DATA_WIDTH-1:0]    mem_req_data,   // 512
    input logic [`VX_MEM_TAG_WIDTH-1:0]     mem_req_tag,    // 56 (55 for SM disabled)
    // vortex inputs
    output logic                            mem_req_ready,

    // Memory response:
    // vortex inputs
    output logic                            mem_rsp_valid,        
    output logic [`VX_MEM_DATA_WIDTH-1:0]   mem_rsp_data,   // 512
    output logic [`VX_MEM_TAG_WIDTH-1:0]    mem_rsp_tag,    // 56 (55 for SM disabled)
    // vortex outputs
    input logic                             mem_rsp_ready,

    // Status:
    // vortex outputs
    input logic                             busy,

    //////////////////////////////////
    // Generic Bus Interface (AHB): //
    //////////////////////////////////

    bus_protocol_if.peripheral_vital        bpif
        // // Vital signals
        // logic wen; // request is a data write
        // logic ren; // request is a data read
        // logic request_stall; // High when protocol should insert wait states in transaction
        // logic [ADDR_WIDTH-1 : 0] addr; // *offset* address of request TODO: Is this good for general use?
        // logic error; // Indicate error condition to bus
        // logic [(DATA_WIDTH/8)-1 : 0] strobe; // byte enable for writes
        // logic [DATA_WIDTH-1 : 0] wdata, rdata; // data lines -- from perspective of bus master. rdata should be data read from peripheral.

        // modport peripheral_vital (
        //     input wen, ren, addr, wdata, strobe,
        //     output rdata, error, request_stall
        // );
);

    ///////////////////////
    // internal signals: //
    ///////////////////////

    // bad address signals
    logic Vortex_bad_address;
    // logic AHB_bad_address;

    // buffered Vortex memory interface signals
    logic                           next_mem_rsp_valid;
    logic [`VX_MEM_DATA_WIDTH-1:0]  next_mem_rsp_data;
    logic [`VX_MEM_TAG_WIDTH-1:0]   next_mem_rsp_tag;

    // reg file signals (bytewise, packed)
    // logic [2**14-1:0][7:0] reg_file;
    // logic [2**14-1:0][7:0] next_reg_file;
    logic [2**LOCAL_MEM_SIZE-1:0][7:0] reg_file;
    logic [2**LOCAL_MEM_SIZE-1:0][7:0] next_reg_file;

    ////////////////
    // registers: //
    ////////////////

    // output buffer registers
    always_ff @ (posedge clk, negedge nRST) begin : VORTEX_MEM_INTERFACE_OUTPUT_BUFFER_FF_LOGIC
        if (~nRST)
        begin
            mem_rsp_valid <= 1'b0;
            mem_rsp_data <= 512'd0;
            mem_rsp_tag <= 26'd0;
        end
        else
        begin
            mem_rsp_valid <= next_mem_rsp_valid;
            mem_rsp_data <= next_mem_rsp_data;
            mem_rsp_tag <= next_mem_rsp_tag;
        end
    end

    // reg file instance
    always_ff @ (posedge clk, negedge nRST) begin : REG_FILE_FF_LOGIC
        if (~nRST)
        begin
            reg_file[0] <= 8'h73;
            reg_file[1] <= 8'h25;
            reg_file[2] <= 8'h10;
            reg_file[3] <= 8'hFC;
            reg_file[4] <= 8'h97;
            reg_file[5] <= 8'h05;
            reg_file[6] <= 8'h00;
            reg_file[7] <= 8'h00;
            reg_file[8] <= 8'h93;
            reg_file[9] <= 8'h85;
            reg_file[10] <= 8'h45;
            reg_file[11] <= 8'h1C;
            reg_file[12] <= 8'h6B;
            reg_file[13] <= 8'h10;
            reg_file[14] <= 8'hB5;
            reg_file[15] <= 8'h00;
            reg_file[16] <= 8'hEF;
            reg_file[17] <= 8'h00;
            reg_file[18] <= 8'h80;
            reg_file[19] <= 8'h1B;
            reg_file[20] <= 8'h13;
            reg_file[21] <= 8'h05;
            reg_file[22] <= 8'h10;
            reg_file[23] <= 8'h00;
            reg_file[24] <= 8'h6B;
            reg_file[25] <= 8'h00;
            reg_file[26] <= 8'h05;
            reg_file[27] <= 8'h00;
            reg_file[28] <= 8'h73;
            reg_file[29] <= 8'h25;
            reg_file[30] <= 8'h10;
            reg_file[31] <= 8'hFC;
            reg_file[32] <= 8'h97;
            reg_file[33] <= 8'h05;
            reg_file[34] <= 8'h00;
            reg_file[35] <= 8'h00;
            reg_file[36] <= 8'h93;
            reg_file[37] <= 8'h85;
            reg_file[38] <= 8'h85;
            reg_file[39] <= 8'h24;
            reg_file[40] <= 8'h6B;
            reg_file[41] <= 8'h10;
            reg_file[42] <= 8'hB5;
            reg_file[43] <= 8'h00;
            reg_file[44] <= 8'hEF;
            reg_file[45] <= 8'h00;
            reg_file[46] <= 8'hC0;
            reg_file[47] <= 8'h23;
            reg_file[48] <= 8'h13;
            reg_file[49] <= 8'h05;
            reg_file[50] <= 8'h10;
            reg_file[51] <= 8'h00;
            reg_file[52] <= 8'h6B;
            reg_file[53] <= 8'h00;
            reg_file[54] <= 8'h05;
            reg_file[55] <= 8'h00;
            reg_file[56] <= 8'h17;
            reg_file[57] <= 8'h55;
            reg_file[58] <= 8'h00;
            reg_file[59] <= 8'h00;
            reg_file[60] <= 8'h13;
            reg_file[61] <= 8'h05;
            reg_file[62] <= 8'h45;
            reg_file[63] <= 8'hCD;
            reg_file[64] <= 8'h17;
            reg_file[65] <= 8'h56;
            reg_file[66] <= 8'h00;
            reg_file[67] <= 8'h00;
            reg_file[68] <= 8'h13;
            reg_file[69] <= 8'h06;
            reg_file[70] <= 8'h06;
            reg_file[71] <= 8'hD8;
            reg_file[72] <= 8'h33;
            reg_file[73] <= 8'h06;
            reg_file[74] <= 8'hA6;
            reg_file[75] <= 8'h40;
            reg_file[76] <= 8'h93;
            reg_file[77] <= 8'h05;
            reg_file[78] <= 8'h00;
            reg_file[79] <= 8'h00;
            reg_file[80] <= 8'hEF;
            reg_file[81] <= 8'h30;
            reg_file[82] <= 8'h00;
            reg_file[83] <= 8'h35;
            reg_file[84] <= 8'h17;
            reg_file[85] <= 8'h05;
            reg_file[86] <= 8'h00;
            reg_file[87] <= 8'h00;
            reg_file[88] <= 8'h13;
            reg_file[89] <= 8'h05;
            reg_file[90] <= 8'h45;
            reg_file[91] <= 8'h30;
            reg_file[92] <= 8'hEF;
            reg_file[93] <= 8'h30;
            reg_file[94] <= 8'h00;
            reg_file[95] <= 8'h1E;
            reg_file[96] <= 8'hEF;
            reg_file[97] <= 8'h00;
            reg_file[98] <= 8'h40;
            reg_file[99] <= 8'h26;
            reg_file[100] <= 8'hEF;
            reg_file[101] <= 8'h00;
            reg_file[102] <= 8'h80;
            reg_file[103] <= 8'h00;
            reg_file[104] <= 8'h6F;
            reg_file[105] <= 8'h30;
            reg_file[106] <= 8'h80;
            reg_file[107] <= 8'h1E;
            reg_file[108] <= 8'h13;
            reg_file[109] <= 8'h01;
            reg_file[110] <= 8'h01;
            reg_file[111] <= 8'hFE;
            reg_file[112] <= 8'h97;
            reg_file[113] <= 8'h57;
            reg_file[114] <= 8'h00;
            reg_file[115] <= 8'h00;
            reg_file[116] <= 8'h93;
            reg_file[117] <= 8'h87;
            reg_file[118] <= 8'h87;
            reg_file[119] <= 8'hC8;
            reg_file[120] <= 8'h23;
            reg_file[121] <= 8'h28;
            reg_file[122] <= 8'h21;
            reg_file[123] <= 8'h01;
            reg_file[124] <= 8'h23;
            reg_file[125] <= 8'h26;
            reg_file[126] <= 8'h31;
            reg_file[127] <= 8'h01;
            reg_file[128] <= 8'h03;
            reg_file[129] <= 8'hA9;
            reg_file[130] <= 8'h07;
            reg_file[131] <= 8'h00;
            reg_file[132] <= 8'h83;
            reg_file[133] <= 8'hA9;
            reg_file[134] <= 8'h47;
            reg_file[135] <= 8'h00;
            reg_file[136] <= 8'h97;
            reg_file[137] <= 8'h57;
            reg_file[138] <= 8'h00;
            reg_file[139] <= 8'h00;
            reg_file[140] <= 8'h93;
            reg_file[141] <= 8'h87;
            reg_file[142] <= 8'h87;
            reg_file[143] <= 8'hC7;
            reg_file[144] <= 8'h23;
            reg_file[145] <= 8'h2C;
            reg_file[146] <= 8'h81;
            reg_file[147] <= 8'h00;
            reg_file[148] <= 8'h23;
            reg_file[149] <= 8'h2A;
            reg_file[150] <= 8'h91;
            reg_file[151] <= 8'h00;
            reg_file[152] <= 8'h03;
            reg_file[153] <= 8'hA4;
            reg_file[154] <= 8'h07;
            reg_file[155] <= 8'h00;
            reg_file[156] <= 8'h83;
            reg_file[157] <= 8'hA4;
            reg_file[158] <= 8'h47;
            reg_file[159] <= 8'h00;
            reg_file[160] <= 8'h13;
            reg_file[161] <= 8'h05;
            reg_file[162] <= 8'h09;
            reg_file[163] <= 8'h00;
            reg_file[164] <= 8'h13;
            reg_file[165] <= 8'h06;
            reg_file[166] <= 8'h04;
            reg_file[167] <= 8'h00;
            reg_file[168] <= 8'h93;
            reg_file[169] <= 8'h86;
            reg_file[170] <= 8'h04;
            reg_file[171] <= 8'h00;
            reg_file[172] <= 8'h93;
            reg_file[173] <= 8'h85;
            reg_file[174] <= 8'h09;
            reg_file[175] <= 8'h00;
            reg_file[176] <= 8'h23;
            reg_file[177] <= 8'h2E;
            reg_file[178] <= 8'h11;
            reg_file[179] <= 8'h00;
            reg_file[180] <= 8'hEF;
            reg_file[181] <= 8'h00;
            reg_file[182] <= 8'hD0;
            reg_file[183] <= 8'h1F;
            reg_file[184] <= 8'h97;
            reg_file[185] <= 8'h57;
            reg_file[186] <= 8'h00;
            reg_file[187] <= 8'h00;
            reg_file[188] <= 8'h93;
            reg_file[189] <= 8'h87;
            reg_file[190] <= 8'h07;
            reg_file[191] <= 8'hC8;
            reg_file[192] <= 8'h13;
            reg_file[193] <= 8'h06;
            reg_file[194] <= 8'h04;
            reg_file[195] <= 8'h00;
            reg_file[196] <= 8'h93;
            reg_file[197] <= 8'h86;
            reg_file[198] <= 8'h04;
            reg_file[199] <= 8'h00;
            reg_file[200] <= 8'h23;
            reg_file[201] <= 8'hA0;
            reg_file[202] <= 8'hA7;
            reg_file[203] <= 8'h00;
            reg_file[204] <= 8'h23;
            reg_file[205] <= 8'hA2;
            reg_file[206] <= 8'hB7;
            reg_file[207] <= 8'h00;
            reg_file[208] <= 8'h13;
            reg_file[209] <= 8'h05;
            reg_file[210] <= 8'h09;
            reg_file[211] <= 8'h00;
            reg_file[212] <= 8'h93;
            reg_file[213] <= 8'h85;
            reg_file[214] <= 8'h09;
            reg_file[215] <= 8'h00;
            reg_file[216] <= 8'hEF;
            reg_file[217] <= 8'h20;
            reg_file[218] <= 8'hC0;
            reg_file[219] <= 8'h59;
            reg_file[220] <= 8'h97;
            reg_file[221] <= 8'h57;
            reg_file[222] <= 8'h00;
            reg_file[223] <= 8'h00;
            reg_file[224] <= 8'h93;
            reg_file[225] <= 8'h87;
            reg_file[226] <= 8'h47;
            reg_file[227] <= 8'hC5;
            reg_file[228] <= 8'h13;
            reg_file[229] <= 8'h06;
            reg_file[230] <= 8'h09;
            reg_file[231] <= 8'h00;
            reg_file[232] <= 8'h93;
            reg_file[233] <= 8'h86;
            reg_file[234] <= 8'h09;
            reg_file[235] <= 8'h00;
            reg_file[236] <= 8'h23;
            reg_file[237] <= 8'hA0;
            reg_file[238] <= 8'hA7;
            reg_file[239] <= 8'h00;
            reg_file[240] <= 8'h23;
            reg_file[241] <= 8'hA2;
            reg_file[242] <= 8'hB7;
            reg_file[243] <= 8'h00;
            reg_file[244] <= 8'h13;
            reg_file[245] <= 8'h05;
            reg_file[246] <= 8'h04;
            reg_file[247] <= 8'h00;
            reg_file[248] <= 8'h93;
            reg_file[249] <= 8'h85;
            reg_file[250] <= 8'h04;
            reg_file[251] <= 8'h00;
            reg_file[252] <= 8'hEF;
            reg_file[253] <= 8'h20;
            reg_file[254] <= 8'h80;
            reg_file[255] <= 8'h57;
            reg_file[256] <= 8'h97;
            reg_file[257] <= 8'h57;
            reg_file[258] <= 8'h00;
            reg_file[259] <= 8'h00;
            reg_file[260] <= 8'h93;
            reg_file[261] <= 8'h87;
            reg_file[262] <= 8'h87;
            reg_file[263] <= 8'hC1;
            reg_file[264] <= 8'h13;
            reg_file[265] <= 8'h06;
            reg_file[266] <= 8'h04;
            reg_file[267] <= 8'h00;
            reg_file[268] <= 8'h93;
            reg_file[269] <= 8'h86;
            reg_file[270] <= 8'h04;
            reg_file[271] <= 8'h00;
            reg_file[272] <= 8'h23;
            reg_file[273] <= 8'hA0;
            reg_file[274] <= 8'hA7;
            reg_file[275] <= 8'h00;
            reg_file[276] <= 8'h23;
            reg_file[277] <= 8'hA2;
            reg_file[278] <= 8'hB7;
            reg_file[279] <= 8'h00;
            reg_file[280] <= 8'h13;
            reg_file[281] <= 8'h05;
            reg_file[282] <= 8'h09;
            reg_file[283] <= 8'h00;
            reg_file[284] <= 8'h93;
            reg_file[285] <= 8'h85;
            reg_file[286] <= 8'h09;
            reg_file[287] <= 8'h00;
            reg_file[288] <= 8'hEF;
            reg_file[289] <= 8'h10;
            reg_file[290] <= 8'hD0;
            reg_file[291] <= 8'h5A;
            reg_file[292] <= 8'h97;
            reg_file[293] <= 8'h57;
            reg_file[294] <= 8'h00;
            reg_file[295] <= 8'h00;
            reg_file[296] <= 8'h93;
            reg_file[297] <= 8'h87;
            reg_file[298] <= 8'h47;
            reg_file[299] <= 8'hC0;
            reg_file[300] <= 8'h13;
            reg_file[301] <= 8'h06;
            reg_file[302] <= 8'h04;
            reg_file[303] <= 8'h00;
            reg_file[304] <= 8'h93;
            reg_file[305] <= 8'h86;
            reg_file[306] <= 8'h04;
            reg_file[307] <= 8'h00;
            reg_file[308] <= 8'h23;
            reg_file[309] <= 8'hA0;
            reg_file[310] <= 8'hA7;
            reg_file[311] <= 8'h00;
            reg_file[312] <= 8'h23;
            reg_file[313] <= 8'hA2;
            reg_file[314] <= 8'hB7;
            reg_file[315] <= 8'h00;
            reg_file[316] <= 8'h13;
            reg_file[317] <= 8'h05;
            reg_file[318] <= 8'h09;
            reg_file[319] <= 8'h00;
            reg_file[320] <= 8'h93;
            reg_file[321] <= 8'h85;
            reg_file[322] <= 8'h09;
            reg_file[323] <= 8'h00;
            reg_file[324] <= 8'hEF;
            reg_file[325] <= 8'h10;
            reg_file[326] <= 8'h80;
            reg_file[327] <= 8'h4C;
            reg_file[328] <= 8'h97;
            reg_file[329] <= 8'h57;
            reg_file[330] <= 8'h00;
            reg_file[331] <= 8'h00;
            reg_file[332] <= 8'h93;
            reg_file[333] <= 8'h87;
            reg_file[334] <= 8'h87;
            reg_file[335] <= 8'hBC;
            reg_file[336] <= 8'h23;
            reg_file[337] <= 8'hA0;
            reg_file[338] <= 8'hA7;
            reg_file[339] <= 8'h00;
            reg_file[340] <= 8'h23;
            reg_file[341] <= 8'hA2;
            reg_file[342] <= 8'hB7;
            reg_file[343] <= 8'h00;
            reg_file[344] <= 8'h13;
            reg_file[345] <= 8'h06;
            reg_file[346] <= 8'h09;
            reg_file[347] <= 8'h00;
            reg_file[348] <= 8'h93;
            reg_file[349] <= 8'h86;
            reg_file[350] <= 8'h09;
            reg_file[351] <= 8'h00;
            reg_file[352] <= 8'h13;
            reg_file[353] <= 8'h05;
            reg_file[354] <= 8'h04;
            reg_file[355] <= 8'h00;
            reg_file[356] <= 8'h93;
            reg_file[357] <= 8'h85;
            reg_file[358] <= 8'h04;
            reg_file[359] <= 8'h00;
            reg_file[360] <= 8'hEF;
            reg_file[361] <= 8'h10;
            reg_file[362] <= 8'h40;
            reg_file[363] <= 8'h4A;
            reg_file[364] <= 8'h97;
            reg_file[365] <= 8'h57;
            reg_file[366] <= 8'h00;
            reg_file[367] <= 8'h00;
            reg_file[368] <= 8'h93;
            reg_file[369] <= 8'h87;
            reg_file[370] <= 8'h47;
            reg_file[371] <= 8'hBB;
            reg_file[372] <= 8'h23;
            reg_file[373] <= 8'hA0;
            reg_file[374] <= 8'hA7;
            reg_file[375] <= 8'h00;
            reg_file[376] <= 8'h23;
            reg_file[377] <= 8'hA2;
            reg_file[378] <= 8'hB7;
            reg_file[379] <= 8'h00;
            reg_file[380] <= 8'h93;
            reg_file[381] <= 8'h07;
            reg_file[382] <= 8'hF0;
            reg_file[383] <= 8'hFF;
            reg_file[384] <= 8'h6B;
            reg_file[385] <= 8'h80;
            reg_file[386] <= 8'h07;
            reg_file[387] <= 8'h00;
            reg_file[388] <= 8'h83;
            reg_file[389] <= 8'h20;
            reg_file[390] <= 8'hC1;
            reg_file[391] <= 8'h01;
            reg_file[392] <= 8'h03;
            reg_file[393] <= 8'h24;
            reg_file[394] <= 8'h81;
            reg_file[395] <= 8'h01;
            reg_file[396] <= 8'h83;
            reg_file[397] <= 8'h24;
            reg_file[398] <= 8'h41;
            reg_file[399] <= 8'h01;
            reg_file[400] <= 8'h03;
            reg_file[401] <= 8'h29;
            reg_file[402] <= 8'h01;
            reg_file[403] <= 8'h01;
            reg_file[404] <= 8'h83;
            reg_file[405] <= 8'h29;
            reg_file[406] <= 8'hC1;
            reg_file[407] <= 8'h00;
            reg_file[408] <= 8'h13;
            reg_file[409] <= 8'h05;
            reg_file[410] <= 8'h10;
            reg_file[411] <= 8'h00;
            reg_file[412] <= 8'h13;
            reg_file[413] <= 8'h01;
            reg_file[414] <= 8'h01;
            reg_file[415] <= 8'h02;
            reg_file[416] <= 8'h67;
            reg_file[417] <= 8'h80;
            reg_file[418] <= 8'h00;
            reg_file[419] <= 8'h00;
            reg_file[420] <= 8'h93;
            reg_file[421] <= 8'h07;
            reg_file[422] <= 8'h00;
            reg_file[423] <= 8'h00;
            reg_file[424] <= 8'h63;
            reg_file[425] <= 8'h88;
            reg_file[426] <= 8'h07;
            reg_file[427] <= 8'h00;
            reg_file[428] <= 8'h37;
            reg_file[429] <= 8'h05;
            reg_file[430] <= 8'h00;
            reg_file[431] <= 8'h80;
            reg_file[432] <= 8'h13;
            reg_file[433] <= 8'h05;
            reg_file[434] <= 8'h85;
            reg_file[435] <= 8'h35;
            reg_file[436] <= 8'h6F;
            reg_file[437] <= 8'h30;
            reg_file[438] <= 8'h80;
            reg_file[439] <= 8'h08;
            reg_file[440] <= 8'h67;
            reg_file[441] <= 8'h80;
            reg_file[442] <= 8'h00;
            reg_file[443] <= 8'h00;
            reg_file[444] <= 8'h93;
            reg_file[445] <= 8'h01;
            reg_file[446] <= 8'h04;
            reg_file[447] <= 8'h00;
            reg_file[448] <= 8'h13;
            reg_file[449] <= 8'h05;
            reg_file[450] <= 8'h00;
            reg_file[451] <= 8'h00;
            reg_file[452] <= 8'h6B;
            reg_file[453] <= 8'h00;
            reg_file[454] <= 8'h05;
            reg_file[455] <= 8'h00;
            reg_file[456] <= 8'h13;
            reg_file[457] <= 8'h05;
            reg_file[458] <= 8'hF0;
            reg_file[459] <= 8'hFF;
            reg_file[460] <= 8'h6B;
            reg_file[461] <= 8'h00;
            reg_file[462] <= 8'h05;
            reg_file[463] <= 8'h00;
            reg_file[464] <= 8'h97;
            reg_file[465] <= 8'h51;
            reg_file[466] <= 8'h00;
            reg_file[467] <= 8'h00;
            reg_file[468] <= 8'h93;
            reg_file[469] <= 8'h81;
            reg_file[470] <= 8'h01;
            reg_file[471] <= 8'hEF;
            reg_file[472] <= 8'h37;
            reg_file[473] <= 8'h01;
            reg_file[474] <= 8'h00;
            reg_file[475] <= 8'hFF;
            reg_file[476] <= 8'h73;
            reg_file[477] <= 8'h25;
            reg_file[478] <= 8'h10;
            reg_file[479] <= 8'hCC;
            reg_file[480] <= 8'h93;
            reg_file[481] <= 8'h15;
            reg_file[482] <= 8'hA5;
            reg_file[483] <= 8'h00;
            reg_file[484] <= 8'h33;
            reg_file[485] <= 8'h01;
            reg_file[486] <= 8'hB1;
            reg_file[487] <= 8'h40;
            reg_file[488] <= 8'h93;
            reg_file[489] <= 8'h05;
            reg_file[490] <= 8'h00;
            reg_file[491] <= 8'h00;
            reg_file[492] <= 8'h33;
            reg_file[493] <= 8'h05;
            reg_file[494] <= 8'hB5;
            reg_file[495] <= 8'h02;
            reg_file[496] <= 8'h17;
            reg_file[497] <= 8'h52;
            reg_file[498] <= 8'h00;
            reg_file[499] <= 8'h00;
            reg_file[500] <= 8'h13;
            reg_file[501] <= 8'h02;
            reg_file[502] <= 8'hF2;
            reg_file[503] <= 8'hC0;
            reg_file[504] <= 8'h33;
            reg_file[505] <= 8'h02;
            reg_file[506] <= 8'hA2;
            reg_file[507] <= 8'h00;
            reg_file[508] <= 8'h13;
            reg_file[509] <= 8'h72;
            reg_file[510] <= 8'h02;
            reg_file[511] <= 8'hFC;
            reg_file[512] <= 8'hF3;
            reg_file[513] <= 8'h26;
            reg_file[514] <= 8'h30;
            reg_file[515] <= 8'hCC;
            reg_file[516] <= 8'h63;
            reg_file[517] <= 8'h86;
            reg_file[518] <= 8'h06;
            reg_file[519] <= 8'h00;
            reg_file[520] <= 8'h13;
            reg_file[521] <= 8'h05;
            reg_file[522] <= 8'h00;
            reg_file[523] <= 8'h00;
            reg_file[524] <= 8'h6B;
            reg_file[525] <= 8'h00;
            reg_file[526] <= 8'h05;
            reg_file[527] <= 8'h00;
            reg_file[528] <= 8'h67;
            reg_file[529] <= 8'h80;
            reg_file[530] <= 8'h00;
            reg_file[531] <= 8'h00;
            reg_file[532] <= 8'h13;
            reg_file[533] <= 8'h05;
            reg_file[534] <= 8'hF0;
            reg_file[535] <= 8'hFF;
            reg_file[536] <= 8'h67;
            reg_file[537] <= 8'h80;
            reg_file[538] <= 8'h00;
            reg_file[539] <= 8'h00;
            reg_file[540] <= 8'h13;
            reg_file[541] <= 8'h05;
            reg_file[542] <= 8'hF0;
            reg_file[543] <= 8'hFF;
            reg_file[544] <= 8'h67;
            reg_file[545] <= 8'h80;
            reg_file[546] <= 8'h00;
            reg_file[547] <= 8'h00;
            reg_file[548] <= 8'h13;
            reg_file[549] <= 8'h05;
            reg_file[550] <= 8'h00;
            reg_file[551] <= 8'h00;
            reg_file[552] <= 8'h67;
            reg_file[553] <= 8'h80;
            reg_file[554] <= 8'h00;
            reg_file[555] <= 8'h00;
            reg_file[556] <= 8'h13;
            reg_file[557] <= 8'h05;
            reg_file[558] <= 8'h00;
            reg_file[559] <= 8'h00;
            reg_file[560] <= 8'h67;
            reg_file[561] <= 8'h80;
            reg_file[562] <= 8'h00;
            reg_file[563] <= 8'h00;
            reg_file[564] <= 8'h13;
            reg_file[565] <= 8'h05;
            reg_file[566] <= 8'hF0;
            reg_file[567] <= 8'hFF;
            reg_file[568] <= 8'h67;
            reg_file[569] <= 8'h80;
            reg_file[570] <= 8'h00;
            reg_file[571] <= 8'h00;
            reg_file[572] <= 8'h13;
            reg_file[573] <= 8'h05;
            reg_file[574] <= 8'hF0;
            reg_file[575] <= 8'hFF;
            reg_file[576] <= 8'h67;
            reg_file[577] <= 8'h80;
            reg_file[578] <= 8'h00;
            reg_file[579] <= 8'h00;
            reg_file[580] <= 8'h73;
            reg_file[581] <= 8'h00;
            reg_file[582] <= 8'h10;
            reg_file[583] <= 8'h00;
            reg_file[584] <= 8'h13;
            reg_file[585] <= 8'h05;
            reg_file[586] <= 8'h00;
            reg_file[587] <= 8'h00;
            reg_file[588] <= 8'h67;
            reg_file[589] <= 8'h80;
            reg_file[590] <= 8'h00;
            reg_file[591] <= 8'h00;
            reg_file[592] <= 8'h13;
            reg_file[593] <= 8'h05;
            reg_file[594] <= 8'h06;
            reg_file[595] <= 8'h00;
            reg_file[596] <= 8'h67;
            reg_file[597] <= 8'h80;
            reg_file[598] <= 8'h00;
            reg_file[599] <= 8'h00;
            reg_file[600] <= 8'h13;
            reg_file[601] <= 8'h05;
            reg_file[602] <= 8'hF0;
            reg_file[603] <= 8'hFF;
            reg_file[604] <= 8'h67;
            reg_file[605] <= 8'h80;
            reg_file[606] <= 8'h00;
            reg_file[607] <= 8'h00;
            reg_file[608] <= 8'h73;
            reg_file[609] <= 8'h25;
            reg_file[610] <= 8'h40;
            reg_file[611] <= 8'hF1;
            reg_file[612] <= 8'h67;
            reg_file[613] <= 8'h80;
            reg_file[614] <= 8'h00;
            reg_file[615] <= 8'h00;
            reg_file[616] <= 8'h13;
            reg_file[617] <= 8'h01;
            reg_file[618] <= 8'h01;
            reg_file[619] <= 8'hFF;
            reg_file[620] <= 8'h23;
            reg_file[621] <= 8'h26;
            reg_file[622] <= 8'h11;
            reg_file[623] <= 8'h00;
            reg_file[624] <= 8'h23;
            reg_file[625] <= 8'h24;
            reg_file[626] <= 8'h81;
            reg_file[627] <= 8'h00;
            reg_file[628] <= 8'h93;
            reg_file[629] <= 8'h07;
            reg_file[630] <= 8'hF0;
            reg_file[631] <= 8'hFF;
            reg_file[632] <= 8'h6B;
            reg_file[633] <= 8'h80;
            reg_file[634] <= 8'h07;
            reg_file[635] <= 8'h00;
            reg_file[636] <= 8'h13;
            reg_file[637] <= 8'h06;
            reg_file[638] <= 8'h00;
            reg_file[639] <= 8'h00;
            reg_file[640] <= 8'h13;
            reg_file[641] <= 8'h05;
            reg_file[642] <= 8'h02;
            reg_file[643] <= 8'h00;
            reg_file[644] <= 8'h97;
            reg_file[645] <= 8'h45;
            reg_file[646] <= 8'h00;
            reg_file[647] <= 8'h00;
            reg_file[648] <= 8'h93;
            reg_file[649] <= 8'h85;
            reg_file[650] <= 8'h45;
            reg_file[651] <= 8'h63;
            reg_file[652] <= 8'h13;
            reg_file[653] <= 8'h04;
            reg_file[654] <= 8'h02;
            reg_file[655] <= 8'h00;
            reg_file[656] <= 8'hEF;
            reg_file[657] <= 8'h20;
            reg_file[658] <= 8'h50;
            reg_file[659] <= 8'h7F;
            reg_file[660] <= 8'h13;
            reg_file[661] <= 8'h05;
            reg_file[662] <= 8'h00;
            reg_file[663] <= 8'h00;
            reg_file[664] <= 8'h13;
            reg_file[665] <= 8'h06;
            reg_file[666] <= 8'h00;
            reg_file[667] <= 8'h00;
            reg_file[668] <= 8'h93;
            reg_file[669] <= 8'h05;
            reg_file[670] <= 8'h00;
            reg_file[671] <= 8'h00;
            reg_file[672] <= 8'h33;
            reg_file[673] <= 8'h05;
            reg_file[674] <= 8'hA4;
            reg_file[675] <= 8'h00;
            reg_file[676] <= 8'hEF;
            reg_file[677] <= 8'h30;
            reg_file[678] <= 8'hC0;
            reg_file[679] <= 8'h0F;
            reg_file[680] <= 8'hF3;
            reg_file[681] <= 8'h27;
            reg_file[682] <= 8'h30;
            reg_file[683] <= 8'hCC;
            reg_file[684] <= 8'h93;
            reg_file[685] <= 8'hB7;
            reg_file[686] <= 8'h17;
            reg_file[687] <= 8'h00;
            reg_file[688] <= 8'h6B;
            reg_file[689] <= 8'h80;
            reg_file[690] <= 8'h07;
            reg_file[691] <= 8'h00;
            reg_file[692] <= 8'h83;
            reg_file[693] <= 8'h20;
            reg_file[694] <= 8'hC1;
            reg_file[695] <= 8'h00;
            reg_file[696] <= 8'h03;
            reg_file[697] <= 8'h24;
            reg_file[698] <= 8'h81;
            reg_file[699] <= 8'h00;
            reg_file[700] <= 8'h13;
            reg_file[701] <= 8'h01;
            reg_file[702] <= 8'h01;
            reg_file[703] <= 8'h01;
            reg_file[704] <= 8'h67;
            reg_file[705] <= 8'h80;
            reg_file[706] <= 8'h00;
            reg_file[707] <= 8'h00;
            reg_file[708] <= 8'h13;
            reg_file[709] <= 8'h01;
            reg_file[710] <= 8'h01;
            reg_file[711] <= 8'hFF;
            reg_file[712] <= 8'h23;
            reg_file[713] <= 8'h24;
            reg_file[714] <= 8'h81;
            reg_file[715] <= 8'h00;
            reg_file[716] <= 8'h23;
            reg_file[717] <= 8'h20;
            reg_file[718] <= 8'h21;
            reg_file[719] <= 8'h01;
            reg_file[720] <= 8'h17;
            reg_file[721] <= 8'h44;
            reg_file[722] <= 8'h00;
            reg_file[723] <= 8'h00;
            reg_file[724] <= 8'h13;
            reg_file[725] <= 8'h04;
            reg_file[726] <= 8'h84;
            reg_file[727] <= 8'h5E;
            reg_file[728] <= 8'h17;
            reg_file[729] <= 8'h49;
            reg_file[730] <= 8'h00;
            reg_file[731] <= 8'h00;
            reg_file[732] <= 8'h13;
            reg_file[733] <= 8'h09;
            reg_file[734] <= 8'h09;
            reg_file[735] <= 8'h5E;
            reg_file[736] <= 8'h33;
            reg_file[737] <= 8'h09;
            reg_file[738] <= 8'h89;
            reg_file[739] <= 8'h40;
            reg_file[740] <= 8'h23;
            reg_file[741] <= 8'h26;
            reg_file[742] <= 8'h11;
            reg_file[743] <= 8'h00;
            reg_file[744] <= 8'h23;
            reg_file[745] <= 8'h22;
            reg_file[746] <= 8'h91;
            reg_file[747] <= 8'h00;
            reg_file[748] <= 8'h13;
            reg_file[749] <= 8'h59;
            reg_file[750] <= 8'h29;
            reg_file[751] <= 8'h40;
            reg_file[752] <= 8'h63;
            reg_file[753] <= 8'h0E;
            reg_file[754] <= 8'h09;
            reg_file[755] <= 8'h00;
            reg_file[756] <= 8'h93;
            reg_file[757] <= 8'h04;
            reg_file[758] <= 8'h00;
            reg_file[759] <= 8'h00;
            reg_file[760] <= 8'h83;
            reg_file[761] <= 8'h27;
            reg_file[762] <= 8'h04;
            reg_file[763] <= 8'h00;
            reg_file[764] <= 8'h93;
            reg_file[765] <= 8'h84;
            reg_file[766] <= 8'h14;
            reg_file[767] <= 8'h00;
            reg_file[768] <= 8'h13;
            reg_file[769] <= 8'h04;
            reg_file[770] <= 8'h44;
            reg_file[771] <= 8'h00;
            reg_file[772] <= 8'hE7;
            reg_file[773] <= 8'h80;
            reg_file[774] <= 8'h07;
            reg_file[775] <= 8'h00;
            reg_file[776] <= 8'hE3;
            reg_file[777] <= 8'h18;
            reg_file[778] <= 8'h99;
            reg_file[779] <= 8'hFE;
            reg_file[780] <= 8'h17;
            reg_file[781] <= 8'h44;
            reg_file[782] <= 8'h00;
            reg_file[783] <= 8'h00;
            reg_file[784] <= 8'h13;
            reg_file[785] <= 8'h04;
            reg_file[786] <= 8'hC4;
            reg_file[787] <= 8'h5A;
            reg_file[788] <= 8'h17;
            reg_file[789] <= 8'h49;
            reg_file[790] <= 8'h00;
            reg_file[791] <= 8'h00;
            reg_file[792] <= 8'h13;
            reg_file[793] <= 8'h09;
            reg_file[794] <= 8'h89;
            reg_file[795] <= 8'h5A;
            reg_file[796] <= 8'h33;
            reg_file[797] <= 8'h09;
            reg_file[798] <= 8'h89;
            reg_file[799] <= 8'h40;
            reg_file[800] <= 8'h13;
            reg_file[801] <= 8'h59;
            reg_file[802] <= 8'h29;
            reg_file[803] <= 8'h40;
            reg_file[804] <= 8'h63;
            reg_file[805] <= 8'h0E;
            reg_file[806] <= 8'h09;
            reg_file[807] <= 8'h00;
            reg_file[808] <= 8'h93;
            reg_file[809] <= 8'h04;
            reg_file[810] <= 8'h00;
            reg_file[811] <= 8'h00;
            reg_file[812] <= 8'h83;
            reg_file[813] <= 8'h27;
            reg_file[814] <= 8'h04;
            reg_file[815] <= 8'h00;
            reg_file[816] <= 8'h93;
            reg_file[817] <= 8'h84;
            reg_file[818] <= 8'h14;
            reg_file[819] <= 8'h00;
            reg_file[820] <= 8'h13;
            reg_file[821] <= 8'h04;
            reg_file[822] <= 8'h44;
            reg_file[823] <= 8'h00;
            reg_file[824] <= 8'hE7;
            reg_file[825] <= 8'h80;
            reg_file[826] <= 8'h07;
            reg_file[827] <= 8'h00;
            reg_file[828] <= 8'hE3;
            reg_file[829] <= 8'h18;
            reg_file[830] <= 8'h99;
            reg_file[831] <= 8'hFE;
            reg_file[832] <= 8'h83;
            reg_file[833] <= 8'h20;
            reg_file[834] <= 8'hC1;
            reg_file[835] <= 8'h00;
            reg_file[836] <= 8'h03;
            reg_file[837] <= 8'h24;
            reg_file[838] <= 8'h81;
            reg_file[839] <= 8'h00;
            reg_file[840] <= 8'h83;
            reg_file[841] <= 8'h24;
            reg_file[842] <= 8'h41;
            reg_file[843] <= 8'h00;
            reg_file[844] <= 8'h03;
            reg_file[845] <= 8'h29;
            reg_file[846] <= 8'h01;
            reg_file[847] <= 8'h00;
            reg_file[848] <= 8'h13;
            reg_file[849] <= 8'h01;
            reg_file[850] <= 8'h01;
            reg_file[851] <= 8'h01;
            reg_file[852] <= 8'h67;
            reg_file[853] <= 8'h80;
            reg_file[854] <= 8'h00;
            reg_file[855] <= 8'h00;
            reg_file[856] <= 8'h13;
            reg_file[857] <= 8'h01;
            reg_file[858] <= 8'h01;
            reg_file[859] <= 8'hFF;
            reg_file[860] <= 8'h23;
            reg_file[861] <= 8'h24;
            reg_file[862] <= 8'h81;
            reg_file[863] <= 8'h00;
            reg_file[864] <= 8'h97;
            reg_file[865] <= 8'h47;
            reg_file[866] <= 8'h00;
            reg_file[867] <= 8'h00;
            reg_file[868] <= 8'h93;
            reg_file[869] <= 8'h87;
            reg_file[870] <= 8'hC7;
            reg_file[871] <= 8'h55;
            reg_file[872] <= 8'h17;
            reg_file[873] <= 8'h44;
            reg_file[874] <= 8'h00;
            reg_file[875] <= 8'h00;
            reg_file[876] <= 8'h13;
            reg_file[877] <= 8'h04;
            reg_file[878] <= 8'h44;
            reg_file[879] <= 8'h55;
            reg_file[880] <= 8'hB3;
            reg_file[881] <= 8'h87;
            reg_file[882] <= 8'h87;
            reg_file[883] <= 8'h40;
            reg_file[884] <= 8'h23;
            reg_file[885] <= 8'h22;
            reg_file[886] <= 8'h91;
            reg_file[887] <= 8'h00;
            reg_file[888] <= 8'h23;
            reg_file[889] <= 8'h26;
            reg_file[890] <= 8'h11;
            reg_file[891] <= 8'h00;
            reg_file[892] <= 8'h93;
            reg_file[893] <= 8'hD4;
            reg_file[894] <= 8'h27;
            reg_file[895] <= 8'h40;
            reg_file[896] <= 8'h63;
            reg_file[897] <= 8'h80;
            reg_file[898] <= 8'h04;
            reg_file[899] <= 8'h02;
            reg_file[900] <= 8'h93;
            reg_file[901] <= 8'h87;
            reg_file[902] <= 8'hC7;
            reg_file[903] <= 8'hFF;
            reg_file[904] <= 8'h33;
            reg_file[905] <= 8'h84;
            reg_file[906] <= 8'h87;
            reg_file[907] <= 8'h00;
            reg_file[908] <= 8'h83;
            reg_file[909] <= 8'h27;
            reg_file[910] <= 8'h04;
            reg_file[911] <= 8'h00;
            reg_file[912] <= 8'h93;
            reg_file[913] <= 8'h84;
            reg_file[914] <= 8'hF4;
            reg_file[915] <= 8'hFF;
            reg_file[916] <= 8'h13;
            reg_file[917] <= 8'h04;
            reg_file[918] <= 8'hC4;
            reg_file[919] <= 8'hFF;
            reg_file[920] <= 8'hE7;
            reg_file[921] <= 8'h80;
            reg_file[922] <= 8'h07;
            reg_file[923] <= 8'h00;
            reg_file[924] <= 8'hE3;
            reg_file[925] <= 8'h98;
            reg_file[926] <= 8'h04;
            reg_file[927] <= 8'hFE;
            reg_file[928] <= 8'h83;
            reg_file[929] <= 8'h20;
            reg_file[930] <= 8'hC1;
            reg_file[931] <= 8'h00;
            reg_file[932] <= 8'h03;
            reg_file[933] <= 8'h24;
            reg_file[934] <= 8'h81;
            reg_file[935] <= 8'h00;
            reg_file[936] <= 8'h83;
            reg_file[937] <= 8'h24;
            reg_file[938] <= 8'h41;
            reg_file[939] <= 8'h00;
            reg_file[940] <= 8'h13;
            reg_file[941] <= 8'h01;
            reg_file[942] <= 8'h01;
            reg_file[943] <= 8'h01;
            reg_file[944] <= 8'h67;
            reg_file[945] <= 8'h80;
            reg_file[946] <= 8'h00;
            reg_file[947] <= 8'h00;
            reg_file[948] <= 8'h13;
            reg_file[949] <= 8'h01;
            reg_file[950] <= 8'h01;
            reg_file[951] <= 8'hFF;
            reg_file[952] <= 8'h23;
            reg_file[953] <= 8'h26;
            reg_file[954] <= 8'h11;
            reg_file[955] <= 8'h00;
            reg_file[956] <= 8'h23;
            reg_file[957] <= 8'h24;
            reg_file[958] <= 8'h81;
            reg_file[959] <= 8'h00;
            reg_file[960] <= 8'h23;
            reg_file[961] <= 8'h22;
            reg_file[962] <= 8'h91;
            reg_file[963] <= 8'h00;
            reg_file[964] <= 8'h23;
            reg_file[965] <= 8'h20;
            reg_file[966] <= 8'h21;
            reg_file[967] <= 8'h01;
            reg_file[968] <= 8'hF3;
            reg_file[969] <= 8'h27;
            reg_file[970] <= 8'h50;
            reg_file[971] <= 8'hCC;
            reg_file[972] <= 8'h73;
            reg_file[973] <= 8'h27;
            reg_file[974] <= 8'h30;
            reg_file[975] <= 8'hCC;
            reg_file[976] <= 8'hF3;
            reg_file[977] <= 8'h26;
            reg_file[978] <= 8'h00;
            reg_file[979] <= 8'hCC;
            reg_file[980] <= 8'hF3;
            reg_file[981] <= 8'h25;
            reg_file[982] <= 8'h00;
            reg_file[983] <= 8'hFC;
            reg_file[984] <= 8'h13;
            reg_file[985] <= 8'h96;
            reg_file[986] <= 8'h27;
            reg_file[987] <= 8'h00;
            reg_file[988] <= 8'h97;
            reg_file[989] <= 8'h57;
            reg_file[990] <= 8'h00;
            reg_file[991] <= 8'h00;
            reg_file[992] <= 8'h93;
            reg_file[993] <= 8'h87;
            reg_file[994] <= 8'h47;
            reg_file[995] <= 8'h96;
            reg_file[996] <= 8'hB3;
            reg_file[997] <= 8'h87;
            reg_file[998] <= 8'hC7;
            reg_file[999] <= 8'h00;
            reg_file[1000] <= 8'h83;
            reg_file[1001] <= 8'hA4;
            reg_file[1002] <= 8'h07;
            reg_file[1003] <= 8'h00;
            reg_file[1004] <= 8'h03;
            reg_file[1005] <= 8'hA4;
            reg_file[1006] <= 8'h04;
            reg_file[1007] <= 8'h01;
            reg_file[1008] <= 8'h03;
            reg_file[1009] <= 8'hA6;
            reg_file[1010] <= 8'hC4;
            reg_file[1011] <= 8'h00;
            reg_file[1012] <= 8'h33;
            reg_file[1013] <= 8'h29;
            reg_file[1014] <= 8'h87;
            reg_file[1015] <= 8'h00;
            reg_file[1016] <= 8'h93;
            reg_file[1017] <= 8'h07;
            reg_file[1018] <= 8'h04;
            reg_file[1019] <= 8'h00;
            reg_file[1020] <= 8'h33;
            reg_file[1021] <= 8'h09;
            reg_file[1022] <= 8'hC9;
            reg_file[1023] <= 8'h00;
            reg_file[1024] <= 8'h33;
            reg_file[1025] <= 8'h04;
            reg_file[1026] <= 8'hE6;
            reg_file[1027] <= 8'h02;
            reg_file[1028] <= 8'h63;
            reg_file[1029] <= 8'h54;
            reg_file[1030] <= 8'hF7;
            reg_file[1031] <= 8'h00;
            reg_file[1032] <= 8'h93;
            reg_file[1033] <= 8'h07;
            reg_file[1034] <= 8'h07;
            reg_file[1035] <= 8'h00;
            reg_file[1036] <= 8'h33;
            reg_file[1037] <= 8'h04;
            reg_file[1038] <= 8'hF4;
            reg_file[1039] <= 8'h00;
            reg_file[1040] <= 8'h03;
            reg_file[1041] <= 8'hA7;
            reg_file[1042] <= 8'h84;
            reg_file[1043] <= 8'h00;
            reg_file[1044] <= 8'h33;
            reg_file[1045] <= 8'h04;
            reg_file[1046] <= 8'hB4;
            reg_file[1047] <= 8'h02;
            reg_file[1048] <= 8'hB3;
            reg_file[1049] <= 8'h07;
            reg_file[1050] <= 8'hD9;
            reg_file[1051] <= 8'h02;
            reg_file[1052] <= 8'h33;
            reg_file[1053] <= 8'h04;
            reg_file[1054] <= 8'hE4;
            reg_file[1055] <= 8'h00;
            reg_file[1056] <= 8'h33;
            reg_file[1057] <= 8'h04;
            reg_file[1058] <= 8'hF4;
            reg_file[1059] <= 8'h00;
            reg_file[1060] <= 8'h33;
            reg_file[1061] <= 8'h09;
            reg_file[1062] <= 8'h89;
            reg_file[1063] <= 8'h00;
            reg_file[1064] <= 8'h63;
            reg_file[1065] <= 8'h5E;
            reg_file[1066] <= 8'h24;
            reg_file[1067] <= 8'h01;
            reg_file[1068] <= 8'h83;
            reg_file[1069] <= 8'hA7;
            reg_file[1070] <= 8'h04;
            reg_file[1071] <= 8'h00;
            reg_file[1072] <= 8'h83;
            reg_file[1073] <= 8'hA5;
            reg_file[1074] <= 8'h44;
            reg_file[1075] <= 8'h00;
            reg_file[1076] <= 8'h13;
            reg_file[1077] <= 8'h05;
            reg_file[1078] <= 8'h04;
            reg_file[1079] <= 8'h00;
            reg_file[1080] <= 8'h13;
            reg_file[1081] <= 8'h04;
            reg_file[1082] <= 8'h14;
            reg_file[1083] <= 8'h00;
            reg_file[1084] <= 8'hE7;
            reg_file[1085] <= 8'h80;
            reg_file[1086] <= 8'h07;
            reg_file[1087] <= 8'h00;
            reg_file[1088] <= 8'hE3;
            reg_file[1089] <= 8'h16;
            reg_file[1090] <= 8'h89;
            reg_file[1091] <= 8'hFE;
            reg_file[1092] <= 8'h03;
            reg_file[1093] <= 8'hA7;
            reg_file[1094] <= 8'h44;
            reg_file[1095] <= 8'h01;
            reg_file[1096] <= 8'h93;
            reg_file[1097] <= 8'h07;
            reg_file[1098] <= 8'h00;
            reg_file[1099] <= 8'h00;
            reg_file[1100] <= 8'h6B;
            reg_file[1101] <= 8'hC0;
            reg_file[1102] <= 8'hE7;
            reg_file[1103] <= 8'h00;
            reg_file[1104] <= 8'h83;
            reg_file[1105] <= 8'h20;
            reg_file[1106] <= 8'hC1;
            reg_file[1107] <= 8'h00;
            reg_file[1108] <= 8'h03;
            reg_file[1109] <= 8'h24;
            reg_file[1110] <= 8'h81;
            reg_file[1111] <= 8'h00;
            reg_file[1112] <= 8'h83;
            reg_file[1113] <= 8'h24;
            reg_file[1114] <= 8'h41;
            reg_file[1115] <= 8'h00;
            reg_file[1116] <= 8'h03;
            reg_file[1117] <= 8'h29;
            reg_file[1118] <= 8'h01;
            reg_file[1119] <= 8'h00;
            reg_file[1120] <= 8'h13;
            reg_file[1121] <= 8'h01;
            reg_file[1122] <= 8'h01;
            reg_file[1123] <= 8'h01;
            reg_file[1124] <= 8'h67;
            reg_file[1125] <= 8'h80;
            reg_file[1126] <= 8'h00;
            reg_file[1127] <= 8'h00;
            reg_file[1128] <= 8'hF3;
            reg_file[1129] <= 8'h27;
            reg_file[1130] <= 8'h50;
            reg_file[1131] <= 8'hCC;
            reg_file[1132] <= 8'h73;
            reg_file[1133] <= 8'h25;
            reg_file[1134] <= 8'h20;
            reg_file[1135] <= 8'hCC;
            reg_file[1136] <= 8'h13;
            reg_file[1137] <= 8'h97;
            reg_file[1138] <= 8'h27;
            reg_file[1139] <= 8'h00;
            reg_file[1140] <= 8'h97;
            reg_file[1141] <= 8'h57;
            reg_file[1142] <= 8'h00;
            reg_file[1143] <= 8'h00;
            reg_file[1144] <= 8'h93;
            reg_file[1145] <= 8'h87;
            reg_file[1146] <= 8'hC7;
            reg_file[1147] <= 8'h8C;
            reg_file[1148] <= 8'hB3;
            reg_file[1149] <= 8'h87;
            reg_file[1150] <= 8'hE7;
            reg_file[1151] <= 8'h00;
            reg_file[1152] <= 8'h83;
            reg_file[1153] <= 8'hA7;
            reg_file[1154] <= 8'h07;
            reg_file[1155] <= 8'h00;
            reg_file[1156] <= 8'h03;
            reg_file[1157] <= 8'hA7;
            reg_file[1158] <= 8'h87;
            reg_file[1159] <= 8'h00;
            reg_file[1160] <= 8'h03;
            reg_file[1161] <= 8'hA3;
            reg_file[1162] <= 8'h07;
            reg_file[1163] <= 8'h00;
            reg_file[1164] <= 8'h83;
            reg_file[1165] <= 8'hA5;
            reg_file[1166] <= 8'h47;
            reg_file[1167] <= 8'h00;
            reg_file[1168] <= 8'h33;
            reg_file[1169] <= 8'h05;
            reg_file[1170] <= 8'hE5;
            reg_file[1171] <= 8'h00;
            reg_file[1172] <= 8'h67;
            reg_file[1173] <= 8'h00;
            reg_file[1174] <= 8'h03;
            reg_file[1175] <= 8'h00;
            reg_file[1176] <= 8'h13;
            reg_file[1177] <= 8'h01;
            reg_file[1178] <= 8'h01;
            reg_file[1179] <= 8'hFF;
            reg_file[1180] <= 8'h23;
            reg_file[1181] <= 8'h26;
            reg_file[1182] <= 8'h11;
            reg_file[1183] <= 8'h00;
            reg_file[1184] <= 8'h93;
            reg_file[1185] <= 8'h07;
            reg_file[1186] <= 8'hF0;
            reg_file[1187] <= 8'hFF;
            reg_file[1188] <= 8'h6B;
            reg_file[1189] <= 8'h80;
            reg_file[1190] <= 8'h07;
            reg_file[1191] <= 8'h00;
            reg_file[1192] <= 8'hEF;
            reg_file[1193] <= 8'hF0;
            reg_file[1194] <= 8'hDF;
            reg_file[1195] <= 8'hF0;
            reg_file[1196] <= 8'hF3;
            reg_file[1197] <= 8'h27;
            reg_file[1198] <= 8'h30;
            reg_file[1199] <= 8'hCC;
            reg_file[1200] <= 8'h93;
            reg_file[1201] <= 8'hB7;
            reg_file[1202] <= 8'h17;
            reg_file[1203] <= 8'h00;
            reg_file[1204] <= 8'h6B;
            reg_file[1205] <= 8'h80;
            reg_file[1206] <= 8'h07;
            reg_file[1207] <= 8'h00;
            reg_file[1208] <= 8'h83;
            reg_file[1209] <= 8'h20;
            reg_file[1210] <= 8'hC1;
            reg_file[1211] <= 8'h00;
            reg_file[1212] <= 8'h13;
            reg_file[1213] <= 8'h01;
            reg_file[1214] <= 8'h01;
            reg_file[1215] <= 8'h01;
            reg_file[1216] <= 8'h67;
            reg_file[1217] <= 8'h80;
            reg_file[1218] <= 8'h00;
            reg_file[1219] <= 8'h00;
            reg_file[1220] <= 8'h13;
            reg_file[1221] <= 8'h01;
            reg_file[1222] <= 8'h01;
            reg_file[1223] <= 8'hFE;
            reg_file[1224] <= 8'h23;
            reg_file[1225] <= 8'h2E;
            reg_file[1226] <= 8'h11;
            reg_file[1227] <= 8'h00;
            reg_file[1228] <= 8'h23;
            reg_file[1229] <= 8'h2C;
            reg_file[1230] <= 8'h81;
            reg_file[1231] <= 8'h00;
            reg_file[1232] <= 8'h23;
            reg_file[1233] <= 8'h2A;
            reg_file[1234] <= 8'h91;
            reg_file[1235] <= 8'h00;
            reg_file[1236] <= 8'h23;
            reg_file[1237] <= 8'h28;
            reg_file[1238] <= 8'h21;
            reg_file[1239] <= 8'h01;
            reg_file[1240] <= 8'h23;
            reg_file[1241] <= 8'h26;
            reg_file[1242] <= 8'h31;
            reg_file[1243] <= 8'h01;
            reg_file[1244] <= 8'h23;
            reg_file[1245] <= 8'h24;
            reg_file[1246] <= 8'h41;
            reg_file[1247] <= 8'h01;
            reg_file[1248] <= 8'hF3;
            reg_file[1249] <= 8'h27;
            reg_file[1250] <= 8'h50;
            reg_file[1251] <= 8'hCC;
            reg_file[1252] <= 8'h73;
            reg_file[1253] <= 8'h27;
            reg_file[1254] <= 8'h30;
            reg_file[1255] <= 8'hCC;
            reg_file[1256] <= 8'hF3;
            reg_file[1257] <= 8'h26;
            reg_file[1258] <= 8'h00;
            reg_file[1259] <= 8'hCC;
            reg_file[1260] <= 8'h73;
            reg_file[1261] <= 8'h25;
            reg_file[1262] <= 8'h00;
            reg_file[1263] <= 8'hFC;
            reg_file[1264] <= 8'h13;
            reg_file[1265] <= 8'h96;
            reg_file[1266] <= 8'h27;
            reg_file[1267] <= 8'h00;
            reg_file[1268] <= 8'h97;
            reg_file[1269] <= 8'h57;
            reg_file[1270] <= 8'h00;
            reg_file[1271] <= 8'h00;
            reg_file[1272] <= 8'h93;
            reg_file[1273] <= 8'h87;
            reg_file[1274] <= 8'hC7;
            reg_file[1275] <= 8'h84;
            reg_file[1276] <= 8'hB3;
            reg_file[1277] <= 8'h87;
            reg_file[1278] <= 8'hC7;
            reg_file[1279] <= 8'h00;
            reg_file[1280] <= 8'h03;
            reg_file[1281] <= 8'hA4;
            reg_file[1282] <= 8'h07;
            reg_file[1283] <= 8'h00;
            reg_file[1284] <= 8'h83;
            reg_file[1285] <= 8'h24;
            reg_file[1286] <= 8'h44;
            reg_file[1287] <= 8'h01;
            reg_file[1288] <= 8'h03;
            reg_file[1289] <= 8'h26;
            reg_file[1290] <= 8'h04;
            reg_file[1291] <= 8'h01;
            reg_file[1292] <= 8'h33;
            reg_file[1293] <= 8'h2A;
            reg_file[1294] <= 8'h97;
            reg_file[1295] <= 8'h00;
            reg_file[1296] <= 8'h93;
            reg_file[1297] <= 8'h87;
            reg_file[1298] <= 8'h04;
            reg_file[1299] <= 8'h00;
            reg_file[1300] <= 8'h33;
            reg_file[1301] <= 8'h0A;
            reg_file[1302] <= 8'hCA;
            reg_file[1303] <= 8'h00;
            reg_file[1304] <= 8'hB3;
            reg_file[1305] <= 8'h04;
            reg_file[1306] <= 8'hE6;
            reg_file[1307] <= 8'h02;
            reg_file[1308] <= 8'h63;
            reg_file[1309] <= 8'h54;
            reg_file[1310] <= 8'hF7;
            reg_file[1311] <= 8'h00;
            reg_file[1312] <= 8'h93;
            reg_file[1313] <= 8'h07;
            reg_file[1314] <= 8'h07;
            reg_file[1315] <= 8'h00;
            reg_file[1316] <= 8'hB3;
            reg_file[1317] <= 8'h84;
            reg_file[1318] <= 8'hF4;
            reg_file[1319] <= 8'h00;
            reg_file[1320] <= 8'h83;
            reg_file[1321] <= 8'h25;
            reg_file[1322] <= 8'h04;
            reg_file[1323] <= 8'h00;
            reg_file[1324] <= 8'h03;
            reg_file[1325] <= 8'h27;
            reg_file[1326] <= 8'hC4;
            reg_file[1327] <= 8'h00;
            reg_file[1328] <= 8'h03;
            reg_file[1329] <= 8'hA9;
            reg_file[1330] <= 8'h05;
            reg_file[1331] <= 8'h00;
            reg_file[1332] <= 8'h83;
            reg_file[1333] <= 8'hA9;
            reg_file[1334] <= 8'h45;
            reg_file[1335] <= 8'h00;
            reg_file[1336] <= 8'hB3;
            reg_file[1337] <= 8'h84;
            reg_file[1338] <= 8'hA4;
            reg_file[1339] <= 8'h02;
            reg_file[1340] <= 8'hB3;
            reg_file[1341] <= 8'h07;
            reg_file[1342] <= 8'hDA;
            reg_file[1343] <= 8'h02;
            reg_file[1344] <= 8'hB3;
            reg_file[1345] <= 8'h84;
            reg_file[1346] <= 8'hE4;
            reg_file[1347] <= 8'h00;
            reg_file[1348] <= 8'hB3;
            reg_file[1349] <= 8'h84;
            reg_file[1350] <= 8'hF4;
            reg_file[1351] <= 8'h00;
            reg_file[1352] <= 8'h33;
            reg_file[1353] <= 8'h0A;
            reg_file[1354] <= 8'h9A;
            reg_file[1355] <= 8'h00;
            reg_file[1356] <= 8'hB3;
            reg_file[1357] <= 8'h09;
            reg_file[1358] <= 8'h39;
            reg_file[1359] <= 8'h03;
            reg_file[1360] <= 8'h63;
            reg_file[1361] <= 8'hC0;
            reg_file[1362] <= 8'h44;
            reg_file[1363] <= 8'h07;
            reg_file[1364] <= 8'h6F;
            reg_file[1365] <= 8'h00;
            reg_file[1366] <= 8'h00;
            reg_file[1367] <= 8'h08;
            reg_file[1368] <= 8'h03;
            reg_file[1369] <= 8'h47;
            reg_file[1370] <= 8'hE4;
            reg_file[1371] <= 8'h01;
            reg_file[1372] <= 8'h83;
            reg_file[1373] <= 8'h46;
            reg_file[1374] <= 8'hD4;
            reg_file[1375] <= 8'h01;
            reg_file[1376] <= 8'h33;
            reg_file[1377] <= 8'hD7;
            reg_file[1378] <= 8'hE4;
            reg_file[1379] <= 8'h40;
            reg_file[1380] <= 8'hB3;
            reg_file[1381] <= 8'h07;
            reg_file[1382] <= 8'h37;
            reg_file[1383] <= 8'h03;
            reg_file[1384] <= 8'hB3;
            reg_file[1385] <= 8'h87;
            reg_file[1386] <= 8'hF4;
            reg_file[1387] <= 8'h40;
            reg_file[1388] <= 8'h63;
            reg_file[1389] <= 8'h80;
            reg_file[1390] <= 8'h06;
            reg_file[1391] <= 8'h06;
            reg_file[1392] <= 8'h83;
            reg_file[1393] <= 8'h46;
            reg_file[1394] <= 8'hF4;
            reg_file[1395] <= 8'h01;
            reg_file[1396] <= 8'hB3;
            reg_file[1397] <= 8'hD6;
            reg_file[1398] <= 8'hD7;
            reg_file[1399] <= 8'h40;
            reg_file[1400] <= 8'hB3;
            reg_file[1401] <= 8'h88;
            reg_file[1402] <= 8'h26;
            reg_file[1403] <= 8'h03;
            reg_file[1404] <= 8'h03;
            reg_file[1405] <= 8'hAE;
            reg_file[1406] <= 8'h45;
            reg_file[1407] <= 8'h01;
            reg_file[1408] <= 8'h03;
            reg_file[1409] <= 8'hA3;
            reg_file[1410] <= 8'h05;
            reg_file[1411] <= 8'h01;
            reg_file[1412] <= 8'h03;
            reg_file[1413] <= 8'hA6;
            reg_file[1414] <= 8'hC5;
            reg_file[1415] <= 8'h00;
            reg_file[1416] <= 8'h03;
            reg_file[1417] <= 8'h28;
            reg_file[1418] <= 8'h44;
            reg_file[1419] <= 8'h00;
            reg_file[1420] <= 8'h03;
            reg_file[1421] <= 8'h25;
            reg_file[1422] <= 8'h84;
            reg_file[1423] <= 8'h00;
            reg_file[1424] <= 8'h93;
            reg_file[1425] <= 8'h84;
            reg_file[1426] <= 8'h14;
            reg_file[1427] <= 8'h00;
            reg_file[1428] <= 8'h33;
            reg_file[1429] <= 8'h07;
            reg_file[1430] <= 8'hC7;
            reg_file[1431] <= 8'h01;
            reg_file[1432] <= 8'hB3;
            reg_file[1433] <= 8'h86;
            reg_file[1434] <= 8'h66;
            reg_file[1435] <= 8'h00;
            reg_file[1436] <= 8'hB3;
            reg_file[1437] <= 8'h87;
            reg_file[1438] <= 8'h17;
            reg_file[1439] <= 8'h41;
            reg_file[1440] <= 8'h33;
            reg_file[1441] <= 8'h86;
            reg_file[1442] <= 8'hC7;
            reg_file[1443] <= 8'h00;
            reg_file[1444] <= 8'hE7;
            reg_file[1445] <= 8'h00;
            reg_file[1446] <= 8'h08;
            reg_file[1447] <= 8'h00;
            reg_file[1448] <= 8'h63;
            reg_file[1449] <= 8'h06;
            reg_file[1450] <= 8'h9A;
            reg_file[1451] <= 8'h02;
            reg_file[1452] <= 8'h83;
            reg_file[1453] <= 8'h25;
            reg_file[1454] <= 8'h04;
            reg_file[1455] <= 8'h00;
            reg_file[1456] <= 8'h83;
            reg_file[1457] <= 8'h47;
            reg_file[1458] <= 8'hC4;
            reg_file[1459] <= 8'h01;
            reg_file[1460] <= 8'hE3;
            reg_file[1461] <= 8'h92;
            reg_file[1462] <= 8'h07;
            reg_file[1463] <= 8'hFA;
            reg_file[1464] <= 8'h33;
            reg_file[1465] <= 8'hC7;
            reg_file[1466] <= 8'h34;
            reg_file[1467] <= 8'h03;
            reg_file[1468] <= 8'h83;
            reg_file[1469] <= 8'h46;
            reg_file[1470] <= 8'hD4;
            reg_file[1471] <= 8'h01;
            reg_file[1472] <= 8'hB3;
            reg_file[1473] <= 8'h07;
            reg_file[1474] <= 8'h37;
            reg_file[1475] <= 8'h03;
            reg_file[1476] <= 8'hB3;
            reg_file[1477] <= 8'h87;
            reg_file[1478] <= 8'hF4;
            reg_file[1479] <= 8'h40;
            reg_file[1480] <= 8'hE3;
            reg_file[1481] <= 8'h94;
            reg_file[1482] <= 8'h06;
            reg_file[1483] <= 8'hFA;
            reg_file[1484] <= 8'hB3;
            reg_file[1485] <= 8'hC6;
            reg_file[1486] <= 8'h27;
            reg_file[1487] <= 8'h03;
            reg_file[1488] <= 8'h6F;
            reg_file[1489] <= 8'hF0;
            reg_file[1490] <= 8'h9F;
            reg_file[1491] <= 8'hFA;
            reg_file[1492] <= 8'h03;
            reg_file[1493] <= 8'h27;
            reg_file[1494] <= 8'h84;
            reg_file[1495] <= 8'h01;
            reg_file[1496] <= 8'h93;
            reg_file[1497] <= 8'h07;
            reg_file[1498] <= 8'h00;
            reg_file[1499] <= 8'h00;
            reg_file[1500] <= 8'h6B;
            reg_file[1501] <= 8'hC0;
            reg_file[1502] <= 8'hE7;
            reg_file[1503] <= 8'h00;
            reg_file[1504] <= 8'h83;
            reg_file[1505] <= 8'h20;
            reg_file[1506] <= 8'hC1;
            reg_file[1507] <= 8'h01;
            reg_file[1508] <= 8'h03;
            reg_file[1509] <= 8'h24;
            reg_file[1510] <= 8'h81;
            reg_file[1511] <= 8'h01;
            reg_file[1512] <= 8'h83;
            reg_file[1513] <= 8'h24;
            reg_file[1514] <= 8'h41;
            reg_file[1515] <= 8'h01;
            reg_file[1516] <= 8'h03;
            reg_file[1517] <= 8'h29;
            reg_file[1518] <= 8'h01;
            reg_file[1519] <= 8'h01;
            reg_file[1520] <= 8'h83;
            reg_file[1521] <= 8'h29;
            reg_file[1522] <= 8'hC1;
            reg_file[1523] <= 8'h00;
            reg_file[1524] <= 8'h03;
            reg_file[1525] <= 8'h2A;
            reg_file[1526] <= 8'h81;
            reg_file[1527] <= 8'h00;
            reg_file[1528] <= 8'h13;
            reg_file[1529] <= 8'h01;
            reg_file[1530] <= 8'h01;
            reg_file[1531] <= 8'h02;
            reg_file[1532] <= 8'h67;
            reg_file[1533] <= 8'h80;
            reg_file[1534] <= 8'h00;
            reg_file[1535] <= 8'h00;
            reg_file[1536] <= 8'h73;
            reg_file[1537] <= 8'h27;
            reg_file[1538] <= 8'h50;
            reg_file[1539] <= 8'hCC;
            reg_file[1540] <= 8'hF3;
            reg_file[1541] <= 8'h27;
            reg_file[1542] <= 8'h20;
            reg_file[1543] <= 8'hCC;
            reg_file[1544] <= 8'h93;
            reg_file[1545] <= 8'h16;
            reg_file[1546] <= 8'h27;
            reg_file[1547] <= 8'h00;
            reg_file[1548] <= 8'h17;
            reg_file[1549] <= 8'h47;
            reg_file[1550] <= 8'h00;
            reg_file[1551] <= 8'h00;
            reg_file[1552] <= 8'h13;
            reg_file[1553] <= 8'h07;
            reg_file[1554] <= 8'h47;
            reg_file[1555] <= 8'h73;
            reg_file[1556] <= 8'h33;
            reg_file[1557] <= 8'h07;
            reg_file[1558] <= 8'hD7;
            reg_file[1559] <= 8'h00;
            reg_file[1560] <= 8'h03;
            reg_file[1561] <= 8'h25;
            reg_file[1562] <= 8'h07;
            reg_file[1563] <= 8'h00;
            reg_file[1564] <= 8'h83;
            reg_file[1565] <= 8'h25;
            reg_file[1566] <= 8'h05;
            reg_file[1567] <= 8'h00;
            reg_file[1568] <= 8'h83;
            reg_file[1569] <= 8'h26;
            reg_file[1570] <= 8'hC5;
            reg_file[1571] <= 8'h00;
            reg_file[1572] <= 8'h03;
            reg_file[1573] <= 8'h47;
            reg_file[1574] <= 8'hC5;
            reg_file[1575] <= 8'h01;
            reg_file[1576] <= 8'h83;
            reg_file[1577] <= 8'hA8;
            reg_file[1578] <= 8'h05;
            reg_file[1579] <= 8'h00;
            reg_file[1580] <= 8'h03;
            reg_file[1581] <= 8'hA6;
            reg_file[1582] <= 8'h45;
            reg_file[1583] <= 8'h00;
            reg_file[1584] <= 8'hB3;
            reg_file[1585] <= 8'h87;
            reg_file[1586] <= 8'hD7;
            reg_file[1587] <= 8'h00;
            reg_file[1588] <= 8'h33;
            reg_file[1589] <= 8'h86;
            reg_file[1590] <= 8'hC8;
            reg_file[1591] <= 8'h02;
            reg_file[1592] <= 8'h63;
            reg_file[1593] <= 8'h08;
            reg_file[1594] <= 8'h07;
            reg_file[1595] <= 8'h04;
            reg_file[1596] <= 8'h03;
            reg_file[1597] <= 8'h47;
            reg_file[1598] <= 8'hE5;
            reg_file[1599] <= 8'h01;
            reg_file[1600] <= 8'h83;
            reg_file[1601] <= 8'h46;
            reg_file[1602] <= 8'hD5;
            reg_file[1603] <= 8'h01;
            reg_file[1604] <= 8'h33;
            reg_file[1605] <= 8'hD7;
            reg_file[1606] <= 8'hE7;
            reg_file[1607] <= 8'h40;
            reg_file[1608] <= 8'h33;
            reg_file[1609] <= 8'h06;
            reg_file[1610] <= 8'hC7;
            reg_file[1611] <= 8'h02;
            reg_file[1612] <= 8'hB3;
            reg_file[1613] <= 8'h87;
            reg_file[1614] <= 8'hC7;
            reg_file[1615] <= 8'h40;
            reg_file[1616] <= 8'h63;
            reg_file[1617] <= 8'h86;
            reg_file[1618] <= 8'h06;
            reg_file[1619] <= 8'h04;
            reg_file[1620] <= 8'h83;
            reg_file[1621] <= 8'h46;
            reg_file[1622] <= 8'hF5;
            reg_file[1623] <= 8'h01;
            reg_file[1624] <= 8'h33;
            reg_file[1625] <= 8'hD8;
            reg_file[1626] <= 8'hD7;
            reg_file[1627] <= 8'h40;
            reg_file[1628] <= 8'h83;
            reg_file[1629] <= 8'hA6;
            reg_file[1630] <= 8'h05;
            reg_file[1631] <= 8'h01;
            reg_file[1632] <= 8'h03;
            reg_file[1633] <= 8'hAE;
            reg_file[1634] <= 8'h45;
            reg_file[1635] <= 8'h01;
            reg_file[1636] <= 8'h03;
            reg_file[1637] <= 8'hA6;
            reg_file[1638] <= 8'hC5;
            reg_file[1639] <= 8'h00;
            reg_file[1640] <= 8'hB3;
            reg_file[1641] <= 8'h06;
            reg_file[1642] <= 8'hD8;
            reg_file[1643] <= 8'h00;
            reg_file[1644] <= 8'h33;
            reg_file[1645] <= 8'h08;
            reg_file[1646] <= 8'h18;
            reg_file[1647] <= 8'h03;
            reg_file[1648] <= 8'h03;
            reg_file[1649] <= 8'h23;
            reg_file[1650] <= 8'h45;
            reg_file[1651] <= 8'h00;
            reg_file[1652] <= 8'h03;
            reg_file[1653] <= 8'h25;
            reg_file[1654] <= 8'h85;
            reg_file[1655] <= 8'h00;
            reg_file[1656] <= 8'h33;
            reg_file[1657] <= 8'h07;
            reg_file[1658] <= 8'hC7;
            reg_file[1659] <= 8'h01;
            reg_file[1660] <= 8'hB3;
            reg_file[1661] <= 8'h87;
            reg_file[1662] <= 8'h07;
            reg_file[1663] <= 8'h41;
            reg_file[1664] <= 8'h33;
            reg_file[1665] <= 8'h86;
            reg_file[1666] <= 8'hC7;
            reg_file[1667] <= 8'h00;
            reg_file[1668] <= 8'h67;
            reg_file[1669] <= 8'h00;
            reg_file[1670] <= 8'h03;
            reg_file[1671] <= 8'h00;
            reg_file[1672] <= 8'h33;
            reg_file[1673] <= 8'hC7;
            reg_file[1674] <= 8'hC7;
            reg_file[1675] <= 8'h02;
            reg_file[1676] <= 8'h83;
            reg_file[1677] <= 8'h46;
            reg_file[1678] <= 8'hD5;
            reg_file[1679] <= 8'h01;
            reg_file[1680] <= 8'h33;
            reg_file[1681] <= 8'h06;
            reg_file[1682] <= 8'hC7;
            reg_file[1683] <= 8'h02;
            reg_file[1684] <= 8'hB3;
            reg_file[1685] <= 8'h87;
            reg_file[1686] <= 8'hC7;
            reg_file[1687] <= 8'h40;
            reg_file[1688] <= 8'hE3;
            reg_file[1689] <= 8'h9E;
            reg_file[1690] <= 8'h06;
            reg_file[1691] <= 8'hFA;
            reg_file[1692] <= 8'h33;
            reg_file[1693] <= 8'hC8;
            reg_file[1694] <= 8'h17;
            reg_file[1695] <= 8'h03;
            reg_file[1696] <= 8'h6F;
            reg_file[1697] <= 8'hF0;
            reg_file[1698] <= 8'hDF;
            reg_file[1699] <= 8'hFB;
            reg_file[1700] <= 8'h13;
            reg_file[1701] <= 8'h01;
            reg_file[1702] <= 8'h01;
            reg_file[1703] <= 8'hFF;
            reg_file[1704] <= 8'h23;
            reg_file[1705] <= 8'h26;
            reg_file[1706] <= 8'h11;
            reg_file[1707] <= 8'h00;
            reg_file[1708] <= 8'h93;
            reg_file[1709] <= 8'h07;
            reg_file[1710] <= 8'hF0;
            reg_file[1711] <= 8'hFF;
            reg_file[1712] <= 8'h6B;
            reg_file[1713] <= 8'h80;
            reg_file[1714] <= 8'h07;
            reg_file[1715] <= 8'h00;
            reg_file[1716] <= 8'hEF;
            reg_file[1717] <= 8'hF0;
            reg_file[1718] <= 8'h1F;
            reg_file[1719] <= 8'hE1;
            reg_file[1720] <= 8'hF3;
            reg_file[1721] <= 8'h27;
            reg_file[1722] <= 8'h30;
            reg_file[1723] <= 8'hCC;
            reg_file[1724] <= 8'h93;
            reg_file[1725] <= 8'hB7;
            reg_file[1726] <= 8'h17;
            reg_file[1727] <= 8'h00;
            reg_file[1728] <= 8'h6B;
            reg_file[1729] <= 8'h80;
            reg_file[1730] <= 8'h07;
            reg_file[1731] <= 8'h00;
            reg_file[1732] <= 8'h83;
            reg_file[1733] <= 8'h20;
            reg_file[1734] <= 8'hC1;
            reg_file[1735] <= 8'h00;
            reg_file[1736] <= 8'h13;
            reg_file[1737] <= 8'h01;
            reg_file[1738] <= 8'h01;
            reg_file[1739] <= 8'h01;
            reg_file[1740] <= 8'h67;
            reg_file[1741] <= 8'h80;
            reg_file[1742] <= 8'h00;
            reg_file[1743] <= 8'h00;
            reg_file[1744] <= 8'h13;
            reg_file[1745] <= 8'h01;
            reg_file[1746] <= 8'h01;
            reg_file[1747] <= 8'hFD;
            reg_file[1748] <= 8'h23;
            reg_file[1749] <= 8'h26;
            reg_file[1750] <= 8'h11;
            reg_file[1751] <= 8'h02;
            reg_file[1752] <= 8'h23;
            reg_file[1753] <= 8'h24;
            reg_file[1754] <= 8'h81;
            reg_file[1755] <= 8'h02;
            reg_file[1756] <= 8'h23;
            reg_file[1757] <= 8'h22;
            reg_file[1758] <= 8'h91;
            reg_file[1759] <= 8'h02;
            reg_file[1760] <= 8'h23;
            reg_file[1761] <= 8'h20;
            reg_file[1762] <= 8'h21;
            reg_file[1763] <= 8'h03;
            reg_file[1764] <= 8'hF3;
            reg_file[1765] <= 8'h26;
            reg_file[1766] <= 8'h20;
            reg_file[1767] <= 8'hFC;
            reg_file[1768] <= 8'hF3;
            reg_file[1769] <= 8'h28;
            reg_file[1770] <= 8'h10;
            reg_file[1771] <= 8'hFC;
            reg_file[1772] <= 8'hF3;
            reg_file[1773] <= 8'h24;
            reg_file[1774] <= 8'h00;
            reg_file[1775] <= 8'hFC;
            reg_file[1776] <= 8'hF3;
            reg_file[1777] <= 8'h27;
            reg_file[1778] <= 8'h50;
            reg_file[1779] <= 8'hCC;
            reg_file[1780] <= 8'h13;
            reg_file[1781] <= 8'h07;
            reg_file[1782] <= 8'hF0;
            reg_file[1783] <= 8'h01;
            reg_file[1784] <= 8'h63;
            reg_file[1785] <= 8'h48;
            reg_file[1786] <= 8'hF7;
            reg_file[1787] <= 8'h08;
            reg_file[1788] <= 8'h33;
            reg_file[1789] <= 8'h88;
            reg_file[1790] <= 8'h14;
            reg_file[1791] <= 8'h03;
            reg_file[1792] <= 8'h13;
            reg_file[1793] <= 8'h07;
            reg_file[1794] <= 8'h10;
            reg_file[1795] <= 8'h00;
            reg_file[1796] <= 8'h63;
            reg_file[1797] <= 8'h54;
            reg_file[1798] <= 8'hA8;
            reg_file[1799] <= 8'h00;
            reg_file[1800] <= 8'h33;
            reg_file[1801] <= 8'h47;
            reg_file[1802] <= 8'h05;
            reg_file[1803] <= 8'h03;
            reg_file[1804] <= 8'h63;
            reg_file[1805] <= 8'hCA;
            reg_file[1806] <= 8'hE6;
            reg_file[1807] <= 8'h08;
            reg_file[1808] <= 8'h63;
            reg_file[1809] <= 8'hDC;
            reg_file[1810] <= 8'hE7;
            reg_file[1811] <= 8'h06;
            reg_file[1812] <= 8'h93;
            reg_file[1813] <= 8'h86;
            reg_file[1814] <= 8'hF6;
            reg_file[1815] <= 8'hFF;
            reg_file[1816] <= 8'h33;
            reg_file[1817] <= 8'h43;
            reg_file[1818] <= 8'hE5;
            reg_file[1819] <= 8'h02;
            reg_file[1820] <= 8'h13;
            reg_file[1821] <= 8'h08;
            reg_file[1822] <= 8'h03;
            reg_file[1823] <= 8'h00;
            reg_file[1824] <= 8'h63;
            reg_file[1825] <= 8'h96;
            reg_file[1826] <= 8'hF6;
            reg_file[1827] <= 8'h00;
            reg_file[1828] <= 8'h33;
            reg_file[1829] <= 8'h65;
            reg_file[1830] <= 8'hE5;
            reg_file[1831] <= 8'h02;
            reg_file[1832] <= 8'h33;
            reg_file[1833] <= 8'h08;
            reg_file[1834] <= 8'h65;
            reg_file[1835] <= 8'h00;
            reg_file[1836] <= 8'h33;
            reg_file[1837] <= 8'h49;
            reg_file[1838] <= 8'h98;
            reg_file[1839] <= 8'h02;
            reg_file[1840] <= 8'h33;
            reg_file[1841] <= 8'h64;
            reg_file[1842] <= 8'h98;
            reg_file[1843] <= 8'h02;
            reg_file[1844] <= 8'h63;
            reg_file[1845] <= 8'h4C;
            reg_file[1846] <= 8'h19;
            reg_file[1847] <= 8'h07;
            reg_file[1848] <= 8'h13;
            reg_file[1849] <= 8'h05;
            reg_file[1850] <= 8'h10;
            reg_file[1851] <= 8'h00;
            reg_file[1852] <= 8'hB3;
            reg_file[1853] <= 8'h46;
            reg_file[1854] <= 8'h19;
            reg_file[1855] <= 8'h03;
            reg_file[1856] <= 8'h63;
            reg_file[1857] <= 8'h86;
            reg_file[1858] <= 8'h06;
            reg_file[1859] <= 8'h00;
            reg_file[1860] <= 8'h13;
            reg_file[1861] <= 8'h85;
            reg_file[1862] <= 8'h06;
            reg_file[1863] <= 8'h00;
            reg_file[1864] <= 8'hB3;
            reg_file[1865] <= 8'h66;
            reg_file[1866] <= 8'h19;
            reg_file[1867] <= 8'h03;
            reg_file[1868] <= 8'h17;
            reg_file[1869] <= 8'h47;
            reg_file[1870] <= 8'h00;
            reg_file[1871] <= 8'h00;
            reg_file[1872] <= 8'h13;
            reg_file[1873] <= 8'h07;
            reg_file[1874] <= 8'h47;
            reg_file[1875] <= 8'h5F;
            reg_file[1876] <= 8'h23;
            reg_file[1877] <= 8'h24;
            reg_file[1878] <= 8'hB1;
            reg_file[1879] <= 8'h00;
            reg_file[1880] <= 8'h23;
            reg_file[1881] <= 8'h26;
            reg_file[1882] <= 8'hC1;
            reg_file[1883] <= 8'h00;
            reg_file[1884] <= 8'h23;
            reg_file[1885] <= 8'h2A;
            reg_file[1886] <= 8'hA1;
            reg_file[1887] <= 8'h00;
            reg_file[1888] <= 8'h23;
            reg_file[1889] <= 8'h2C;
            reg_file[1890] <= 8'hD1;
            reg_file[1891] <= 8'h00;
            reg_file[1892] <= 8'h23;
            reg_file[1893] <= 8'h2E;
            reg_file[1894] <= 8'h01;
            reg_file[1895] <= 8'h00;
            reg_file[1896] <= 8'h33;
            reg_file[1897] <= 8'h03;
            reg_file[1898] <= 8'hF3;
            reg_file[1899] <= 8'h02;
            reg_file[1900] <= 8'h93;
            reg_file[1901] <= 8'h97;
            reg_file[1902] <= 8'h27;
            reg_file[1903] <= 8'h00;
            reg_file[1904] <= 8'hB3;
            reg_file[1905] <= 8'h07;
            reg_file[1906] <= 8'hF7;
            reg_file[1907] <= 8'h00;
            reg_file[1908] <= 8'h13;
            reg_file[1909] <= 8'h07;
            reg_file[1910] <= 8'h81;
            reg_file[1911] <= 8'h00;
            reg_file[1912] <= 8'h23;
            reg_file[1913] <= 8'hA0;
            reg_file[1914] <= 8'hE7;
            reg_file[1915] <= 8'h00;
            reg_file[1916] <= 8'h23;
            reg_file[1917] <= 8'h28;
            reg_file[1918] <= 8'h61;
            reg_file[1919] <= 8'h00;
            reg_file[1920] <= 8'h63;
            reg_file[1921] <= 8'h4C;
            reg_file[1922] <= 8'h20;
            reg_file[1923] <= 8'h03;
            reg_file[1924] <= 8'h63;
            reg_file[1925] <= 8'h16;
            reg_file[1926] <= 8'h04;
            reg_file[1927] <= 8'h06;
            reg_file[1928] <= 8'h83;
            reg_file[1929] <= 8'h20;
            reg_file[1930] <= 8'hC1;
            reg_file[1931] <= 8'h02;
            reg_file[1932] <= 8'h03;
            reg_file[1933] <= 8'h24;
            reg_file[1934] <= 8'h81;
            reg_file[1935] <= 8'h02;
            reg_file[1936] <= 8'h83;
            reg_file[1937] <= 8'h24;
            reg_file[1938] <= 8'h41;
            reg_file[1939] <= 8'h02;
            reg_file[1940] <= 8'h03;
            reg_file[1941] <= 8'h29;
            reg_file[1942] <= 8'h01;
            reg_file[1943] <= 8'h02;
            reg_file[1944] <= 8'h13;
            reg_file[1945] <= 8'h01;
            reg_file[1946] <= 8'h01;
            reg_file[1947] <= 8'h03;
            reg_file[1948] <= 8'h67;
            reg_file[1949] <= 8'h80;
            reg_file[1950] <= 8'h00;
            reg_file[1951] <= 8'h00;
            reg_file[1952] <= 8'h13;
            reg_file[1953] <= 8'h87;
            reg_file[1954] <= 8'h06;
            reg_file[1955] <= 8'h00;
            reg_file[1956] <= 8'hE3;
            reg_file[1957] <= 8'hC8;
            reg_file[1958] <= 8'hE7;
            reg_file[1959] <= 8'hF6;
            reg_file[1960] <= 8'h6F;
            reg_file[1961] <= 8'hF0;
            reg_file[1962] <= 8'h1F;
            reg_file[1963] <= 8'hFE;
            reg_file[1964] <= 8'h93;
            reg_file[1965] <= 8'h06;
            reg_file[1966] <= 8'h00;
            reg_file[1967] <= 8'h00;
            reg_file[1968] <= 8'h13;
            reg_file[1969] <= 8'h05;
            reg_file[1970] <= 8'h10;
            reg_file[1971] <= 8'h00;
            reg_file[1972] <= 8'h6F;
            reg_file[1973] <= 8'hF0;
            reg_file[1974] <= 8'h9F;
            reg_file[1975] <= 8'hF9;
            reg_file[1976] <= 8'h93;
            reg_file[1977] <= 8'h07;
            reg_file[1978] <= 8'h09;
            reg_file[1979] <= 8'h00;
            reg_file[1980] <= 8'h63;
            reg_file[1981] <= 8'hD4;
            reg_file[1982] <= 8'h28;
            reg_file[1983] <= 8'h01;
            reg_file[1984] <= 8'h93;
            reg_file[1985] <= 8'h87;
            reg_file[1986] <= 8'h08;
            reg_file[1987] <= 8'h00;
            reg_file[1988] <= 8'h23;
            reg_file[1989] <= 8'h2E;
            reg_file[1990] <= 8'hF1;
            reg_file[1991] <= 8'h00;
            reg_file[1992] <= 8'h17;
            reg_file[1993] <= 8'h07;
            reg_file[1994] <= 8'h00;
            reg_file[1995] <= 8'h00;
            reg_file[1996] <= 8'h13;
            reg_file[1997] <= 8'h07;
            reg_file[1998] <= 8'h07;
            reg_file[1999] <= 8'hCD;
            reg_file[2000] <= 8'h6B;
            reg_file[2001] <= 8'h90;
            reg_file[2002] <= 8'hE7;
            reg_file[2003] <= 8'h00;
            reg_file[2004] <= 8'h93;
            reg_file[2005] <= 8'h07;
            reg_file[2006] <= 8'hF0;
            reg_file[2007] <= 8'hFF;
            reg_file[2008] <= 8'h6B;
            reg_file[2009] <= 8'h80;
            reg_file[2010] <= 8'h07;
            reg_file[2011] <= 8'h00;
            reg_file[2012] <= 8'hEF;
            reg_file[2013] <= 8'hF0;
            reg_file[2014] <= 8'h9F;
            reg_file[2015] <= 8'hBD;
            reg_file[2016] <= 8'hF3;
            reg_file[2017] <= 8'h27;
            reg_file[2018] <= 8'h30;
            reg_file[2019] <= 8'hCC;
            reg_file[2020] <= 8'h93;
            reg_file[2021] <= 8'hB7;
            reg_file[2022] <= 8'h17;
            reg_file[2023] <= 8'h00;
            reg_file[2024] <= 8'h6B;
            reg_file[2025] <= 8'h80;
            reg_file[2026] <= 8'h07;
            reg_file[2027] <= 8'h00;
            reg_file[2028] <= 8'hE3;
            reg_file[2029] <= 8'h0E;
            reg_file[2030] <= 8'h04;
            reg_file[2031] <= 8'hF8;
            reg_file[2032] <= 8'hB3;
            reg_file[2033] <= 8'h04;
            reg_file[2034] <= 8'h99;
            reg_file[2035] <= 8'h02;
            reg_file[2036] <= 8'h13;
            reg_file[2037] <= 8'h09;
            reg_file[2038] <= 8'h10;
            reg_file[2039] <= 8'h00;
            reg_file[2040] <= 8'h33;
            reg_file[2041] <= 8'h18;
            reg_file[2042] <= 8'h89;
            reg_file[2043] <= 8'h00;
            reg_file[2044] <= 8'h13;
            reg_file[2045] <= 8'h08;
            reg_file[2046] <= 8'hF8;
            reg_file[2047] <= 8'hFF;
            reg_file[2048] <= 8'h23;
            reg_file[2049] <= 8'h28;
            reg_file[2050] <= 8'h91;
            reg_file[2051] <= 8'h00;
            reg_file[2052] <= 8'h6B;
            reg_file[2053] <= 8'h00;
            reg_file[2054] <= 8'h08;
            reg_file[2055] <= 8'h00;
            reg_file[2056] <= 8'hEF;
            reg_file[2057] <= 8'hF0;
            reg_file[2058] <= 8'h1F;
            reg_file[2059] <= 8'hC6;
            reg_file[2060] <= 8'h6B;
            reg_file[2061] <= 8'h00;
            reg_file[2062] <= 8'h09;
            reg_file[2063] <= 8'h00;
            reg_file[2064] <= 8'h83;
            reg_file[2065] <= 8'h20;
            reg_file[2066] <= 8'hC1;
            reg_file[2067] <= 8'h02;
            reg_file[2068] <= 8'h03;
            reg_file[2069] <= 8'h24;
            reg_file[2070] <= 8'h81;
            reg_file[2071] <= 8'h02;
            reg_file[2072] <= 8'h83;
            reg_file[2073] <= 8'h24;
            reg_file[2074] <= 8'h41;
            reg_file[2075] <= 8'h02;
            reg_file[2076] <= 8'h03;
            reg_file[2077] <= 8'h29;
            reg_file[2078] <= 8'h01;
            reg_file[2079] <= 8'h02;
            reg_file[2080] <= 8'h13;
            reg_file[2081] <= 8'h01;
            reg_file[2082] <= 8'h01;
            reg_file[2083] <= 8'h03;
            reg_file[2084] <= 8'h67;
            reg_file[2085] <= 8'h80;
            reg_file[2086] <= 8'h00;
            reg_file[2087] <= 8'h00;
            reg_file[2088] <= 8'h13;
            reg_file[2089] <= 8'h01;
            reg_file[2090] <= 8'h01;
            reg_file[2091] <= 8'hFD;
            reg_file[2092] <= 8'h23;
            reg_file[2093] <= 8'h26;
            reg_file[2094] <= 8'h11;
            reg_file[2095] <= 8'h02;
            reg_file[2096] <= 8'h23;
            reg_file[2097] <= 8'h24;
            reg_file[2098] <= 8'h81;
            reg_file[2099] <= 8'h02;
            reg_file[2100] <= 8'h23;
            reg_file[2101] <= 8'h22;
            reg_file[2102] <= 8'h91;
            reg_file[2103] <= 8'h02;
            reg_file[2104] <= 8'h23;
            reg_file[2105] <= 8'h20;
            reg_file[2106] <= 8'h21;
            reg_file[2107] <= 8'h03;
            reg_file[2108] <= 8'hF3;
            reg_file[2109] <= 8'h28;
            reg_file[2110] <= 8'h20;
            reg_file[2111] <= 8'hFC;
            reg_file[2112] <= 8'h73;
            reg_file[2113] <= 8'h23;
            reg_file[2114] <= 8'h10;
            reg_file[2115] <= 8'hFC;
            reg_file[2116] <= 8'hF3;
            reg_file[2117] <= 8'h24;
            reg_file[2118] <= 8'h00;
            reg_file[2119] <= 8'hFC;
            reg_file[2120] <= 8'hF3;
            reg_file[2121] <= 8'h27;
            reg_file[2122] <= 8'h50;
            reg_file[2123] <= 8'hCC;
            reg_file[2124] <= 8'h13;
            reg_file[2125] <= 8'h07;
            reg_file[2126] <= 8'hF0;
            reg_file[2127] <= 8'h01;
            reg_file[2128] <= 8'h63;
            reg_file[2129] <= 8'h46;
            reg_file[2130] <= 8'hF7;
            reg_file[2131] <= 8'h0E;
            reg_file[2132] <= 8'h03;
            reg_file[2133] <= 8'h2E;
            reg_file[2134] <= 8'h05;
            reg_file[2135] <= 8'h00;
            reg_file[2136] <= 8'h83;
            reg_file[2137] <= 8'h26;
            reg_file[2138] <= 8'h45;
            reg_file[2139] <= 8'h00;
            reg_file[2140] <= 8'h03;
            reg_file[2141] <= 8'h28;
            reg_file[2142] <= 8'h85;
            reg_file[2143] <= 8'h00;
            reg_file[2144] <= 8'hB3;
            reg_file[2145] <= 8'h0E;
            reg_file[2146] <= 8'h93;
            reg_file[2147] <= 8'h02;
            reg_file[2148] <= 8'h13;
            reg_file[2149] <= 8'h07;
            reg_file[2150] <= 8'h10;
            reg_file[2151] <= 8'h00;
            reg_file[2152] <= 8'hB3;
            reg_file[2153] <= 8'h06;
            reg_file[2154] <= 8'hDE;
            reg_file[2155] <= 8'h02;
            reg_file[2156] <= 8'h33;
            reg_file[2157] <= 8'h88;
            reg_file[2158] <= 8'h06;
            reg_file[2159] <= 8'h03;
            reg_file[2160] <= 8'h63;
            reg_file[2161] <= 8'hD4;
            reg_file[2162] <= 8'h0E;
            reg_file[2163] <= 8'h01;
            reg_file[2164] <= 8'h33;
            reg_file[2165] <= 8'h47;
            reg_file[2166] <= 8'hD8;
            reg_file[2167] <= 8'h03;
            reg_file[2168] <= 8'h63;
            reg_file[2169] <= 8'hCE;
            reg_file[2170] <= 8'hE8;
            reg_file[2171] <= 8'h0C;
            reg_file[2172] <= 8'h63;
            reg_file[2173] <= 8'hD0;
            reg_file[2174] <= 8'hE7;
            reg_file[2175] <= 8'h0C;
            reg_file[2176] <= 8'h93;
            reg_file[2177] <= 8'h88;
            reg_file[2178] <= 8'hF8;
            reg_file[2179] <= 8'hFF;
            reg_file[2180] <= 8'h33;
            reg_file[2181] <= 8'h4F;
            reg_file[2182] <= 8'hE8;
            reg_file[2183] <= 8'h02;
            reg_file[2184] <= 8'h13;
            reg_file[2185] <= 8'h04;
            reg_file[2186] <= 8'h0F;
            reg_file[2187] <= 8'h00;
            reg_file[2188] <= 8'h63;
            reg_file[2189] <= 8'h96;
            reg_file[2190] <= 8'hF8;
            reg_file[2191] <= 8'h00;
            reg_file[2192] <= 8'h33;
            reg_file[2193] <= 8'h67;
            reg_file[2194] <= 8'hE8;
            reg_file[2195] <= 8'h02;
            reg_file[2196] <= 8'h33;
            reg_file[2197] <= 8'h04;
            reg_file[2198] <= 8'hE7;
            reg_file[2199] <= 8'h01;
            reg_file[2200] <= 8'h33;
            reg_file[2201] <= 8'h49;
            reg_file[2202] <= 8'h94;
            reg_file[2203] <= 8'h02;
            reg_file[2204] <= 8'h33;
            reg_file[2205] <= 8'h64;
            reg_file[2206] <= 8'h94;
            reg_file[2207] <= 8'h02;
            reg_file[2208] <= 8'h63;
            reg_file[2209] <= 8'h40;
            reg_file[2210] <= 8'h69;
            reg_file[2211] <= 8'h0C;
            reg_file[2212] <= 8'h93;
            reg_file[2213] <= 8'h02;
            reg_file[2214] <= 8'h10;
            reg_file[2215] <= 8'h00;
            reg_file[2216] <= 8'hB3;
            reg_file[2217] <= 8'h4F;
            reg_file[2218] <= 8'h69;
            reg_file[2219] <= 8'h02;
            reg_file[2220] <= 8'h63;
            reg_file[2221] <= 8'h86;
            reg_file[2222] <= 8'h0F;
            reg_file[2223] <= 8'h00;
            reg_file[2224] <= 8'h93;
            reg_file[2225] <= 8'h82;
            reg_file[2226] <= 8'h0F;
            reg_file[2227] <= 8'h00;
            reg_file[2228] <= 8'hB3;
            reg_file[2229] <= 8'h6F;
            reg_file[2230] <= 8'h69;
            reg_file[2231] <= 8'h02;
            reg_file[2232] <= 8'hD3;
            reg_file[2233] <= 8'hF7;
            reg_file[2234] <= 8'h06;
            reg_file[2235] <= 8'hD0;
            reg_file[2236] <= 8'h93;
            reg_file[2237] <= 8'h08;
            reg_file[2238] <= 8'hFE;
            reg_file[2239] <= 8'hFF;
            reg_file[2240] <= 8'h93;
            reg_file[2241] <= 8'h8E;
            reg_file[2242] <= 8'hF6;
            reg_file[2243] <= 8'hFF;
            reg_file[2244] <= 8'h53;
            reg_file[2245] <= 8'h88;
            reg_file[2246] <= 8'h07;
            reg_file[2247] <= 8'hE0;
            reg_file[2248] <= 8'hD3;
            reg_file[2249] <= 8'h77;
            reg_file[2250] <= 8'h0E;
            reg_file[2251] <= 8'hD0;
            reg_file[2252] <= 8'hB3;
            reg_file[2253] <= 8'hF6;
            reg_file[2254] <= 8'hDE;
            reg_file[2255] <= 8'h00;
            reg_file[2256] <= 8'h33;
            reg_file[2257] <= 8'hFE;
            reg_file[2258] <= 8'hC8;
            reg_file[2259] <= 8'h01;
            reg_file[2260] <= 8'h53;
            reg_file[2261] <= 8'h87;
            reg_file[2262] <= 8'h07;
            reg_file[2263] <= 8'hE0;
            reg_file[2264] <= 8'h13;
            reg_file[2265] <= 8'h58;
            reg_file[2266] <= 8'h78;
            reg_file[2267] <= 8'h41;
            reg_file[2268] <= 8'h97;
            reg_file[2269] <= 8'h48;
            reg_file[2270] <= 8'h00;
            reg_file[2271] <= 8'h00;
            reg_file[2272] <= 8'h93;
            reg_file[2273] <= 8'h88;
            reg_file[2274] <= 8'h48;
            reg_file[2275] <= 8'h46;
            reg_file[2276] <= 8'h13;
            reg_file[2277] <= 8'h57;
            reg_file[2278] <= 8'h77;
            reg_file[2279] <= 8'h41;
            reg_file[2280] <= 8'h93;
            reg_file[2281] <= 8'hB6;
            reg_file[2282] <= 8'h16;
            reg_file[2283] <= 8'h00;
            reg_file[2284] <= 8'h13;
            reg_file[2285] <= 8'h3E;
            reg_file[2286] <= 8'h1E;
            reg_file[2287] <= 8'h00;
            reg_file[2288] <= 8'h13;
            reg_file[2289] <= 8'h08;
            reg_file[2290] <= 8'h18;
            reg_file[2291] <= 8'hF8;
            reg_file[2292] <= 8'h13;
            reg_file[2293] <= 8'h07;
            reg_file[2294] <= 8'h17;
            reg_file[2295] <= 8'hF8;
            reg_file[2296] <= 8'h23;
            reg_file[2297] <= 8'h20;
            reg_file[2298] <= 8'hA1;
            reg_file[2299] <= 8'h00;
            reg_file[2300] <= 8'h23;
            reg_file[2301] <= 8'h22;
            reg_file[2302] <= 8'hB1;
            reg_file[2303] <= 8'h00;
            reg_file[2304] <= 8'h23;
            reg_file[2305] <= 8'h24;
            reg_file[2306] <= 8'hC1;
            reg_file[2307] <= 8'h00;
            reg_file[2308] <= 8'h23;
            reg_file[2309] <= 8'h28;
            reg_file[2310] <= 8'h51;
            reg_file[2311] <= 8'h00;
            reg_file[2312] <= 8'h23;
            reg_file[2313] <= 8'h2A;
            reg_file[2314] <= 8'hF1;
            reg_file[2315] <= 8'h01;
            reg_file[2316] <= 8'h23;
            reg_file[2317] <= 8'h2C;
            reg_file[2318] <= 8'h01;
            reg_file[2319] <= 8'h00;
            reg_file[2320] <= 8'h23;
            reg_file[2321] <= 8'h0E;
            reg_file[2322] <= 8'hD1;
            reg_file[2323] <= 8'h00;
            reg_file[2324] <= 8'hA3;
            reg_file[2325] <= 8'h0E;
            reg_file[2326] <= 8'hC1;
            reg_file[2327] <= 8'h01;
            reg_file[2328] <= 8'h23;
            reg_file[2329] <= 8'h0F;
            reg_file[2330] <= 8'h01;
            reg_file[2331] <= 8'h01;
            reg_file[2332] <= 8'hA3;
            reg_file[2333] <= 8'h0F;
            reg_file[2334] <= 8'hE1;
            reg_file[2335] <= 8'h00;
            reg_file[2336] <= 8'h33;
            reg_file[2337] <= 8'h0F;
            reg_file[2338] <= 8'hFF;
            reg_file[2339] <= 8'h02;
            reg_file[2340] <= 8'h93;
            reg_file[2341] <= 8'h97;
            reg_file[2342] <= 8'h27;
            reg_file[2343] <= 8'h00;
            reg_file[2344] <= 8'hB3;
            reg_file[2345] <= 8'h87;
            reg_file[2346] <= 8'hF8;
            reg_file[2347] <= 8'h00;
            reg_file[2348] <= 8'h23;
            reg_file[2349] <= 8'hA0;
            reg_file[2350] <= 8'h27;
            reg_file[2351] <= 8'h00;
            reg_file[2352] <= 8'h23;
            reg_file[2353] <= 8'h26;
            reg_file[2354] <= 8'hE1;
            reg_file[2355] <= 8'h01;
            reg_file[2356] <= 8'h63;
            reg_file[2357] <= 8'h4C;
            reg_file[2358] <= 8'h20;
            reg_file[2359] <= 8'h03;
            reg_file[2360] <= 8'h63;
            reg_file[2361] <= 8'h16;
            reg_file[2362] <= 8'h04;
            reg_file[2363] <= 8'h06;
            reg_file[2364] <= 8'h83;
            reg_file[2365] <= 8'h20;
            reg_file[2366] <= 8'hC1;
            reg_file[2367] <= 8'h02;
            reg_file[2368] <= 8'h03;
            reg_file[2369] <= 8'h24;
            reg_file[2370] <= 8'h81;
            reg_file[2371] <= 8'h02;
            reg_file[2372] <= 8'h83;
            reg_file[2373] <= 8'h24;
            reg_file[2374] <= 8'h41;
            reg_file[2375] <= 8'h02;
            reg_file[2376] <= 8'h03;
            reg_file[2377] <= 8'h29;
            reg_file[2378] <= 8'h01;
            reg_file[2379] <= 8'h02;
            reg_file[2380] <= 8'h13;
            reg_file[2381] <= 8'h01;
            reg_file[2382] <= 8'h01;
            reg_file[2383] <= 8'h03;
            reg_file[2384] <= 8'h67;
            reg_file[2385] <= 8'h80;
            reg_file[2386] <= 8'h00;
            reg_file[2387] <= 8'h00;
            reg_file[2388] <= 8'h13;
            reg_file[2389] <= 8'h87;
            reg_file[2390] <= 8'h08;
            reg_file[2391] <= 8'h00;
            reg_file[2392] <= 8'hE3;
            reg_file[2393] <= 8'hC4;
            reg_file[2394] <= 8'hE7;
            reg_file[2395] <= 8'hF2;
            reg_file[2396] <= 8'h6F;
            reg_file[2397] <= 8'hF0;
            reg_file[2398] <= 8'h1F;
            reg_file[2399] <= 8'hFE;
            reg_file[2400] <= 8'h93;
            reg_file[2401] <= 8'h0F;
            reg_file[2402] <= 8'h00;
            reg_file[2403] <= 8'h00;
            reg_file[2404] <= 8'h93;
            reg_file[2405] <= 8'h02;
            reg_file[2406] <= 8'h10;
            reg_file[2407] <= 8'h00;
            reg_file[2408] <= 8'h6F;
            reg_file[2409] <= 8'hF0;
            reg_file[2410] <= 8'h1F;
            reg_file[2411] <= 8'hF5;
            reg_file[2412] <= 8'h93;
            reg_file[2413] <= 8'h07;
            reg_file[2414] <= 8'h09;
            reg_file[2415] <= 8'h00;
            reg_file[2416] <= 8'h63;
            reg_file[2417] <= 8'h54;
            reg_file[2418] <= 8'h23;
            reg_file[2419] <= 8'h01;
            reg_file[2420] <= 8'h93;
            reg_file[2421] <= 8'h07;
            reg_file[2422] <= 8'h03;
            reg_file[2423] <= 8'h00;
            reg_file[2424] <= 8'h23;
            reg_file[2425] <= 8'h2C;
            reg_file[2426] <= 8'hF1;
            reg_file[2427] <= 8'h00;
            reg_file[2428] <= 8'h17;
            reg_file[2429] <= 8'h07;
            reg_file[2430] <= 8'h00;
            reg_file[2431] <= 8'h00;
            reg_file[2432] <= 8'h13;
            reg_file[2433] <= 8'h07;
            reg_file[2434] <= 8'h87;
            reg_file[2435] <= 8'hD2;
            reg_file[2436] <= 8'h6B;
            reg_file[2437] <= 8'h90;
            reg_file[2438] <= 8'hE7;
            reg_file[2439] <= 8'h00;
            reg_file[2440] <= 8'h93;
            reg_file[2441] <= 8'h07;
            reg_file[2442] <= 8'hF0;
            reg_file[2443] <= 8'hFF;
            reg_file[2444] <= 8'h6B;
            reg_file[2445] <= 8'h80;
            reg_file[2446] <= 8'h07;
            reg_file[2447] <= 8'h00;
            reg_file[2448] <= 8'hEF;
            reg_file[2449] <= 8'hF0;
            reg_file[2450] <= 8'h5F;
            reg_file[2451] <= 8'hB3;
            reg_file[2452] <= 8'hF3;
            reg_file[2453] <= 8'h27;
            reg_file[2454] <= 8'h30;
            reg_file[2455] <= 8'hCC;
            reg_file[2456] <= 8'h93;
            reg_file[2457] <= 8'hB7;
            reg_file[2458] <= 8'h17;
            reg_file[2459] <= 8'h00;
            reg_file[2460] <= 8'h6B;
            reg_file[2461] <= 8'h80;
            reg_file[2462] <= 8'h07;
            reg_file[2463] <= 8'h00;
            reg_file[2464] <= 8'hE3;
            reg_file[2465] <= 8'h0E;
            reg_file[2466] <= 8'h04;
            reg_file[2467] <= 8'hF8;
            reg_file[2468] <= 8'hB3;
            reg_file[2469] <= 8'h04;
            reg_file[2470] <= 8'h99;
            reg_file[2471] <= 8'h02;
            reg_file[2472] <= 8'h13;
            reg_file[2473] <= 8'h09;
            reg_file[2474] <= 8'h10;
            reg_file[2475] <= 8'h00;
            reg_file[2476] <= 8'h33;
            reg_file[2477] <= 8'h14;
            reg_file[2478] <= 8'h89;
            reg_file[2479] <= 8'h00;
            reg_file[2480] <= 8'h13;
            reg_file[2481] <= 8'h04;
            reg_file[2482] <= 8'hF4;
            reg_file[2483] <= 8'hFF;
            reg_file[2484] <= 8'h23;
            reg_file[2485] <= 8'h26;
            reg_file[2486] <= 8'h91;
            reg_file[2487] <= 8'h00;
            reg_file[2488] <= 8'h6B;
            reg_file[2489] <= 8'h00;
            reg_file[2490] <= 8'h04;
            reg_file[2491] <= 8'h00;
            reg_file[2492] <= 8'hEF;
            reg_file[2493] <= 8'hF0;
            reg_file[2494] <= 8'h5F;
            reg_file[2495] <= 8'hC4;
            reg_file[2496] <= 8'h6B;
            reg_file[2497] <= 8'h00;
            reg_file[2498] <= 8'h09;
            reg_file[2499] <= 8'h00;
            reg_file[2500] <= 8'h83;
            reg_file[2501] <= 8'h20;
            reg_file[2502] <= 8'hC1;
            reg_file[2503] <= 8'h02;
            reg_file[2504] <= 8'h03;
            reg_file[2505] <= 8'h24;
            reg_file[2506] <= 8'h81;
            reg_file[2507] <= 8'h02;
            reg_file[2508] <= 8'h83;
            reg_file[2509] <= 8'h24;
            reg_file[2510] <= 8'h41;
            reg_file[2511] <= 8'h02;
            reg_file[2512] <= 8'h03;
            reg_file[2513] <= 8'h29;
            reg_file[2514] <= 8'h01;
            reg_file[2515] <= 8'h02;
            reg_file[2516] <= 8'h13;
            reg_file[2517] <= 8'h01;
            reg_file[2518] <= 8'h01;
            reg_file[2519] <= 8'h03;
            reg_file[2520] <= 8'h67;
            reg_file[2521] <= 8'h80;
            reg_file[2522] <= 8'h00;
            reg_file[2523] <= 8'h00;
            reg_file[2524] <= 8'h13;
            reg_file[2525] <= 8'h01;
            reg_file[2526] <= 8'h81;
            reg_file[2527] <= 8'hFE;
            reg_file[2528] <= 8'h23;
            reg_file[2529] <= 8'h2A;
            reg_file[2530] <= 8'h11;
            reg_file[2531] <= 8'h00;
            reg_file[2532] <= 8'h23;
            reg_file[2533] <= 8'h28;
            reg_file[2534] <= 8'h41;
            reg_file[2535] <= 8'h01;
            reg_file[2536] <= 8'h23;
            reg_file[2537] <= 8'h26;
            reg_file[2538] <= 8'h31;
            reg_file[2539] <= 8'h01;
            reg_file[2540] <= 8'h23;
            reg_file[2541] <= 8'h24;
            reg_file[2542] <= 8'h21;
            reg_file[2543] <= 8'h01;
            reg_file[2544] <= 8'h23;
            reg_file[2545] <= 8'h22;
            reg_file[2546] <= 8'h91;
            reg_file[2547] <= 8'h00;
            reg_file[2548] <= 8'h23;
            reg_file[2549] <= 8'h20;
            reg_file[2550] <= 8'h81;
            reg_file[2551] <= 8'h00;
            reg_file[2552] <= 8'h13;
            reg_file[2553] <= 8'h0A;
            reg_file[2554] <= 8'h05;
            reg_file[2555] <= 8'h00;
            reg_file[2556] <= 8'h93;
            reg_file[2557] <= 8'h89;
            reg_file[2558] <= 8'h05;
            reg_file[2559] <= 8'h00;
            reg_file[2560] <= 8'h73;
            reg_file[2561] <= 8'h29;
            reg_file[2562] <= 8'h00;
            reg_file[2563] <= 8'hFC;
            reg_file[2564] <= 8'hF3;
            reg_file[2565] <= 8'h24;
            reg_file[2566] <= 8'h00;
            reg_file[2567] <= 8'hCC;
            reg_file[2568] <= 8'h13;
            reg_file[2569] <= 8'h04;
            reg_file[2570] <= 8'h00;
            reg_file[2571] <= 8'h00;
            reg_file[2572] <= 8'hB3;
            reg_file[2573] <= 8'h02;
            reg_file[2574] <= 8'h94;
            reg_file[2575] <= 8'h40;
            reg_file[2576] <= 8'h13;
            reg_file[2577] <= 8'hB3;
            reg_file[2578] <= 8'h12;
            reg_file[2579] <= 8'h00;
            reg_file[2580] <= 8'h6B;
            reg_file[2581] <= 8'h20;
            reg_file[2582] <= 8'h03;
            reg_file[2583] <= 8'h00;
            reg_file[2584] <= 8'h63;
            reg_file[2585] <= 8'h96;
            reg_file[2586] <= 8'h02;
            reg_file[2587] <= 8'h00;
            reg_file[2588] <= 8'h13;
            reg_file[2589] <= 8'h85;
            reg_file[2590] <= 8'h09;
            reg_file[2591] <= 8'h00;
            reg_file[2592] <= 8'hE7;
            reg_file[2593] <= 8'h00;
            reg_file[2594] <= 8'h0A;
            reg_file[2595] <= 8'h00;
            reg_file[2596] <= 8'h6B;
            reg_file[2597] <= 8'h30;
            reg_file[2598] <= 8'h00;
            reg_file[2599] <= 8'h00;
            reg_file[2600] <= 8'h13;
            reg_file[2601] <= 8'h04;
            reg_file[2602] <= 8'h14;
            reg_file[2603] <= 8'h00;
            reg_file[2604] <= 8'hE3;
            reg_file[2605] <= 8'h40;
            reg_file[2606] <= 8'h24;
            reg_file[2607] <= 8'hFF;
            reg_file[2608] <= 8'h83;
            reg_file[2609] <= 8'h20;
            reg_file[2610] <= 8'h41;
            reg_file[2611] <= 8'h01;
            reg_file[2612] <= 8'h03;
            reg_file[2613] <= 8'h2A;
            reg_file[2614] <= 8'h01;
            reg_file[2615] <= 8'h01;
            reg_file[2616] <= 8'h83;
            reg_file[2617] <= 8'h29;
            reg_file[2618] <= 8'hC1;
            reg_file[2619] <= 8'h00;
            reg_file[2620] <= 8'h03;
            reg_file[2621] <= 8'h29;
            reg_file[2622] <= 8'h81;
            reg_file[2623] <= 8'h00;
            reg_file[2624] <= 8'h83;
            reg_file[2625] <= 8'h24;
            reg_file[2626] <= 8'h41;
            reg_file[2627] <= 8'h00;
            reg_file[2628] <= 8'h03;
            reg_file[2629] <= 8'h24;
            reg_file[2630] <= 8'h01;
            reg_file[2631] <= 8'h00;
            reg_file[2632] <= 8'h13;
            reg_file[2633] <= 8'h01;
            reg_file[2634] <= 8'h81;
            reg_file[2635] <= 8'h01;
            reg_file[2636] <= 8'h67;
            reg_file[2637] <= 8'h80;
            reg_file[2638] <= 8'h00;
            reg_file[2639] <= 8'h00;
            reg_file[2640] <= 8'h13;
            reg_file[2641] <= 8'h05;
            reg_file[2642] <= 8'hF0;
            reg_file[2643] <= 8'hFF;
            reg_file[2644] <= 8'h67;
            reg_file[2645] <= 8'h80;
            reg_file[2646] <= 8'h00;
            reg_file[2647] <= 8'h00;
            reg_file[2648] <= 8'h13;
            reg_file[2649] <= 8'h05;
            reg_file[2650] <= 8'hF0;
            reg_file[2651] <= 8'hFF;
            reg_file[2652] <= 8'h67;
            reg_file[2653] <= 8'h80;
            reg_file[2654] <= 8'h00;
            reg_file[2655] <= 8'h00;
            reg_file[2656] <= 8'h13;
            reg_file[2657] <= 8'h05;
            reg_file[2658] <= 8'hF0;
            reg_file[2659] <= 8'hFF;
            reg_file[2660] <= 8'h67;
            reg_file[2661] <= 8'h80;
            reg_file[2662] <= 8'h00;
            reg_file[2663] <= 8'h00;
            reg_file[2664] <= 8'h13;
            reg_file[2665] <= 8'h05;
            reg_file[2666] <= 8'hF0;
            reg_file[2667] <= 8'hFF;
            reg_file[2668] <= 8'h67;
            reg_file[2669] <= 8'h80;
            reg_file[2670] <= 8'h00;
            reg_file[2671] <= 8'h00;
            reg_file[2672] <= 8'h13;
            reg_file[2673] <= 8'h05;
            reg_file[2674] <= 8'hF0;
            reg_file[2675] <= 8'hFF;
            reg_file[2676] <= 8'h67;
            reg_file[2677] <= 8'h80;
            reg_file[2678] <= 8'h00;
            reg_file[2679] <= 8'h00;
            reg_file[2680] <= 8'h13;
            reg_file[2681] <= 8'h05;
            reg_file[2682] <= 8'hF0;
            reg_file[2683] <= 8'hFF;
            reg_file[2684] <= 8'h67;
            reg_file[2685] <= 8'h80;
            reg_file[2686] <= 8'h00;
            reg_file[2687] <= 8'h00;
            reg_file[2688] <= 8'h13;
            reg_file[2689] <= 8'h05;
            reg_file[2690] <= 8'h00;
            reg_file[2691] <= 8'h00;
            reg_file[2692] <= 8'h67;
            reg_file[2693] <= 8'h80;
            reg_file[2694] <= 8'h00;
            reg_file[2695] <= 8'h00;
            reg_file[2696] <= 8'h13;
            reg_file[2697] <= 8'h05;
            reg_file[2698] <= 8'hF0;
            reg_file[2699] <= 8'hFF;
            reg_file[2700] <= 8'h67;
            reg_file[2701] <= 8'h80;
            reg_file[2702] <= 8'h00;
            reg_file[2703] <= 8'h00;
            reg_file[2704] <= 8'h13;
            reg_file[2705] <= 8'h05;
            reg_file[2706] <= 8'hF0;
            reg_file[2707] <= 8'hFF;
            reg_file[2708] <= 8'h67;
            reg_file[2709] <= 8'h80;
            reg_file[2710] <= 8'h00;
            reg_file[2711] <= 8'h00;
            reg_file[2712] <= 8'h13;
            reg_file[2713] <= 8'h05;
            reg_file[2714] <= 8'hF0;
            reg_file[2715] <= 8'hFF;
            reg_file[2716] <= 8'h67;
            reg_file[2717] <= 8'h80;
            reg_file[2718] <= 8'h00;
            reg_file[2719] <= 8'h00;
            reg_file[2720] <= 8'h13;
            reg_file[2721] <= 8'h05;
            reg_file[2722] <= 8'hF0;
            reg_file[2723] <= 8'hFF;
            reg_file[2724] <= 8'h67;
            reg_file[2725] <= 8'h80;
            reg_file[2726] <= 8'h00;
            reg_file[2727] <= 8'h00;
            reg_file[2728] <= 8'h13;
            reg_file[2729] <= 8'h05;
            reg_file[2730] <= 8'hF0;
            reg_file[2731] <= 8'hFF;
            reg_file[2732] <= 8'h67;
            reg_file[2733] <= 8'h80;
            reg_file[2734] <= 8'h00;
            reg_file[2735] <= 8'h00;
            reg_file[2736] <= 8'h13;
            reg_file[2737] <= 8'h01;
            reg_file[2738] <= 8'h01;
            reg_file[2739] <= 8'hFE;
            reg_file[2740] <= 8'h23;
            reg_file[2741] <= 8'h2E;
            reg_file[2742] <= 8'h11;
            reg_file[2743] <= 8'h00;
            reg_file[2744] <= 8'h23;
            reg_file[2745] <= 8'h2C;
            reg_file[2746] <= 8'h81;
            reg_file[2747] <= 8'h00;
            reg_file[2748] <= 8'h23;
            reg_file[2749] <= 8'h2A;
            reg_file[2750] <= 8'h91;
            reg_file[2751] <= 8'h00;
            reg_file[2752] <= 8'h23;
            reg_file[2753] <= 8'h28;
            reg_file[2754] <= 8'h21;
            reg_file[2755] <= 8'h01;
            reg_file[2756] <= 8'h23;
            reg_file[2757] <= 8'h26;
            reg_file[2758] <= 8'h31;
            reg_file[2759] <= 8'h01;
            reg_file[2760] <= 8'h23;
            reg_file[2761] <= 8'h24;
            reg_file[2762] <= 8'h41;
            reg_file[2763] <= 8'h01;
            reg_file[2764] <= 8'hF3;
            reg_file[2765] <= 8'h29;
            reg_file[2766] <= 8'h20;
            reg_file[2767] <= 8'h00;
            reg_file[2768] <= 8'hB7;
            reg_file[2769] <= 8'h08;
            reg_file[2770] <= 8'h10;
            reg_file[2771] <= 8'h00;
            reg_file[2772] <= 8'h93;
            reg_file[2773] <= 8'h88;
            reg_file[2774] <= 8'hF8;
            reg_file[2775] <= 8'hFF;
            reg_file[2776] <= 8'hB3;
            reg_file[2777] <= 8'hF7;
            reg_file[2778] <= 8'hB8;
            reg_file[2779] <= 8'h00;
            reg_file[2780] <= 8'h13;
            reg_file[2781] <= 8'hD4;
            reg_file[2782] <= 8'h45;
            reg_file[2783] <= 8'h01;
            reg_file[2784] <= 8'h93;
            reg_file[2785] <= 8'hD4;
            reg_file[2786] <= 8'hF5;
            reg_file[2787] <= 8'h01;
            reg_file[2788] <= 8'hB3;
            reg_file[2789] <= 8'hF5;
            reg_file[2790] <= 8'hD8;
            reg_file[2791] <= 8'h00;
            reg_file[2792] <= 8'h93;
            reg_file[2793] <= 8'hD8;
            reg_file[2794] <= 8'h46;
            reg_file[2795] <= 8'h01;
            reg_file[2796] <= 8'h13;
            reg_file[2797] <= 8'h57;
            reg_file[2798] <= 8'hD5;
            reg_file[2799] <= 8'h01;
            reg_file[2800] <= 8'h13;
            reg_file[2801] <= 8'h74;
            reg_file[2802] <= 8'hF4;
            reg_file[2803] <= 8'h7F;
            reg_file[2804] <= 8'h93;
            reg_file[2805] <= 8'h97;
            reg_file[2806] <= 8'h37;
            reg_file[2807] <= 8'h00;
            reg_file[2808] <= 8'h93;
            reg_file[2809] <= 8'hF8;
            reg_file[2810] <= 8'hF8;
            reg_file[2811] <= 8'h7F;
            reg_file[2812] <= 8'hB3;
            reg_file[2813] <= 8'h67;
            reg_file[2814] <= 8'hF7;
            reg_file[2815] <= 8'h00;
            reg_file[2816] <= 8'h13;
            reg_file[2817] <= 8'hDE;
            reg_file[2818] <= 8'hF6;
            reg_file[2819] <= 8'h01;
            reg_file[2820] <= 8'h13;
            reg_file[2821] <= 8'h57;
            reg_file[2822] <= 8'hD6;
            reg_file[2823] <= 8'h01;
            reg_file[2824] <= 8'h93;
            reg_file[2825] <= 8'h95;
            reg_file[2826] <= 8'h35;
            reg_file[2827] <= 8'h00;
            reg_file[2828] <= 8'hB3;
            reg_file[2829] <= 8'h06;
            reg_file[2830] <= 8'h14;
            reg_file[2831] <= 8'h41;
            reg_file[2832] <= 8'h13;
            reg_file[2833] <= 8'h15;
            reg_file[2834] <= 8'h35;
            reg_file[2835] <= 8'h00;
            reg_file[2836] <= 8'h33;
            reg_file[2837] <= 8'h67;
            reg_file[2838] <= 8'hB7;
            reg_file[2839] <= 8'h00;
            reg_file[2840] <= 8'h13;
            reg_file[2841] <= 8'h16;
            reg_file[2842] <= 8'h36;
            reg_file[2843] <= 8'h00;
            reg_file[2844] <= 8'h13;
            reg_file[2845] <= 8'h88;
            reg_file[2846] <= 8'h06;
            reg_file[2847] <= 8'h00;
            reg_file[2848] <= 8'h63;
            reg_file[2849] <= 8'h94;
            reg_file[2850] <= 8'hC4;
            reg_file[2851] <= 8'h43;
            reg_file[2852] <= 8'h63;
            reg_file[2853] <= 8'h56;
            reg_file[2854] <= 8'hD0;
            reg_file[2855] <= 8'h14;
            reg_file[2856] <= 8'h63;
            reg_file[2857] <= 8'h9E;
            reg_file[2858] <= 8'h08;
            reg_file[2859] <= 8'h04;
            reg_file[2860] <= 8'hB3;
            reg_file[2861] <= 8'h66;
            reg_file[2862] <= 8'hC7;
            reg_file[2863] <= 8'h00;
            reg_file[2864] <= 8'h63;
            reg_file[2865] <= 8'h98;
            reg_file[2866] <= 8'h06;
            reg_file[2867] <= 8'h00;
            reg_file[2868] <= 8'h13;
            reg_file[2869] <= 8'h07;
            reg_file[2870] <= 8'hF0;
            reg_file[2871] <= 8'h7F;
            reg_file[2872] <= 8'h63;
            reg_file[2873] <= 8'h14;
            reg_file[2874] <= 8'hE8;
            reg_file[2875] <= 8'h36;
            reg_file[2876] <= 8'h6F;
            reg_file[2877] <= 8'h00;
            reg_file[2878] <= 8'hC0;
            reg_file[2879] <= 8'h02;
            reg_file[2880] <= 8'h93;
            reg_file[2881] <= 8'h06;
            reg_file[2882] <= 8'hF8;
            reg_file[2883] <= 8'hFF;
            reg_file[2884] <= 8'h63;
            reg_file[2885] <= 8'h9E;
            reg_file[2886] <= 8'h06;
            reg_file[2887] <= 8'h00;
            reg_file[2888] <= 8'h33;
            reg_file[2889] <= 8'h06;
            reg_file[2890] <= 8'hA6;
            reg_file[2891] <= 8'h00;
            reg_file[2892] <= 8'hB3;
            reg_file[2893] <= 8'h87;
            reg_file[2894] <= 8'hE7;
            reg_file[2895] <= 8'h00;
            reg_file[2896] <= 8'hB3;
            reg_file[2897] <= 8'h36;
            reg_file[2898] <= 8'hA6;
            reg_file[2899] <= 8'h00;
            reg_file[2900] <= 8'h33;
            reg_file[2901] <= 8'h87;
            reg_file[2902] <= 8'hD7;
            reg_file[2903] <= 8'h00;
            reg_file[2904] <= 8'h13;
            reg_file[2905] <= 8'h08;
            reg_file[2906] <= 8'h10;
            reg_file[2907] <= 8'h00;
            reg_file[2908] <= 8'h6F;
            reg_file[2909] <= 8'h00;
            reg_file[2910] <= 8'h00;
            reg_file[2911] <= 8'h0A;
            reg_file[2912] <= 8'h93;
            reg_file[2913] <= 8'h05;
            reg_file[2914] <= 8'hF0;
            reg_file[2915] <= 8'h7F;
            reg_file[2916] <= 8'h63;
            reg_file[2917] <= 8'h18;
            reg_file[2918] <= 8'hB8;
            reg_file[2919] <= 8'h04;
            reg_file[2920] <= 8'h33;
            reg_file[2921] <= 8'hE7;
            reg_file[2922] <= 8'hA7;
            reg_file[2923] <= 8'h00;
            reg_file[2924] <= 8'hE3;
            reg_file[2925] <= 8'h02;
            reg_file[2926] <= 8'h07;
            reg_file[2927] <= 8'h0E;
            reg_file[2928] <= 8'h13;
            reg_file[2929] <= 8'h97;
            reg_file[2930] <= 8'h97;
            reg_file[2931] <= 8'h00;
            reg_file[2932] <= 8'h13;
            reg_file[2933] <= 8'h04;
            reg_file[2934] <= 8'h00;
            reg_file[2935] <= 8'h00;
            reg_file[2936] <= 8'h63;
            reg_file[2937] <= 8'h40;
            reg_file[2938] <= 8'h07;
            reg_file[2939] <= 8'h28;
            reg_file[2940] <= 8'h93;
            reg_file[2941] <= 8'h08;
            reg_file[2942] <= 8'h00;
            reg_file[2943] <= 8'h01;
            reg_file[2944] <= 8'h6F;
            reg_file[2945] <= 8'h00;
            reg_file[2946] <= 8'h80;
            reg_file[2947] <= 8'h27;
            reg_file[2948] <= 8'h93;
            reg_file[2949] <= 8'h05;
            reg_file[2950] <= 8'hF0;
            reg_file[2951] <= 8'h7F;
            reg_file[2952] <= 8'h63;
            reg_file[2953] <= 8'h12;
            reg_file[2954] <= 8'hB4;
            reg_file[2955] <= 8'h02;
            reg_file[2956] <= 8'h33;
            reg_file[2957] <= 8'hE7;
            reg_file[2958] <= 8'hA7;
            reg_file[2959] <= 8'h00;
            reg_file[2960] <= 8'hE3;
            reg_file[2961] <= 8'h06;
            reg_file[2962] <= 8'h07;
            reg_file[2963] <= 8'h0C;
            reg_file[2964] <= 8'h13;
            reg_file[2965] <= 8'h97;
            reg_file[2966] <= 8'h97;
            reg_file[2967] <= 8'h00;
            reg_file[2968] <= 8'h13;
            reg_file[2969] <= 8'h08;
            reg_file[2970] <= 8'hF0;
            reg_file[2971] <= 8'h7F;
            reg_file[2972] <= 8'h13;
            reg_file[2973] <= 8'h04;
            reg_file[2974] <= 8'h00;
            reg_file[2975] <= 8'h00;
            reg_file[2976] <= 8'hE3;
            reg_file[2977] <= 8'h5E;
            reg_file[2978] <= 8'h07;
            reg_file[2979] <= 8'hFC;
            reg_file[2980] <= 8'h93;
            reg_file[2981] <= 8'h08;
            reg_file[2982] <= 8'h00;
            reg_file[2983] <= 8'h00;
            reg_file[2984] <= 8'h6F;
            reg_file[2985] <= 8'h00;
            reg_file[2986] <= 8'h00;
            reg_file[2987] <= 8'h25;
            reg_file[2988] <= 8'hB7;
            reg_file[2989] <= 8'h05;
            reg_file[2990] <= 8'h80;
            reg_file[2991] <= 8'h00;
            reg_file[2992] <= 8'h33;
            reg_file[2993] <= 8'h67;
            reg_file[2994] <= 8'hB7;
            reg_file[2995] <= 8'h00;
            reg_file[2996] <= 8'h93;
            reg_file[2997] <= 8'h05;
            reg_file[2998] <= 8'h80;
            reg_file[2999] <= 8'h03;
            reg_file[3000] <= 8'h63;
            reg_file[3001] <= 8'hC6;
            reg_file[3002] <= 8'hD5;
            reg_file[3003] <= 8'h0A;
            reg_file[3004] <= 8'h93;
            reg_file[3005] <= 8'h05;
            reg_file[3006] <= 8'hF0;
            reg_file[3007] <= 8'h01;
            reg_file[3008] <= 8'h63;
            reg_file[3009] <= 8'hC8;
            reg_file[3010] <= 8'hD5;
            reg_file[3011] <= 8'h06;
            reg_file[3012] <= 8'h13;
            reg_file[3013] <= 8'h08;
            reg_file[3014] <= 8'h00;
            reg_file[3015] <= 8'h02;
            reg_file[3016] <= 8'h33;
            reg_file[3017] <= 8'h08;
            reg_file[3018] <= 8'hD8;
            reg_file[3019] <= 8'h40;
            reg_file[3020] <= 8'hB3;
            reg_file[3021] <= 8'h58;
            reg_file[3022] <= 8'hD6;
            reg_file[3023] <= 8'h00;
            reg_file[3024] <= 8'hB3;
            reg_file[3025] <= 8'h15;
            reg_file[3026] <= 8'h07;
            reg_file[3027] <= 8'h01;
            reg_file[3028] <= 8'h33;
            reg_file[3029] <= 8'h16;
            reg_file[3030] <= 8'h06;
            reg_file[3031] <= 8'h01;
            reg_file[3032] <= 8'hB3;
            reg_file[3033] <= 8'hE5;
            reg_file[3034] <= 8'h15;
            reg_file[3035] <= 8'h01;
            reg_file[3036] <= 8'h33;
            reg_file[3037] <= 8'h36;
            reg_file[3038] <= 8'hC0;
            reg_file[3039] <= 8'h00;
            reg_file[3040] <= 8'h33;
            reg_file[3041] <= 8'hE6;
            reg_file[3042] <= 8'hC5;
            reg_file[3043] <= 8'h00;
            reg_file[3044] <= 8'hB3;
            reg_file[3045] <= 8'h56;
            reg_file[3046] <= 8'hD7;
            reg_file[3047] <= 8'h00;
            reg_file[3048] <= 8'h33;
            reg_file[3049] <= 8'h06;
            reg_file[3050] <= 8'hA6;
            reg_file[3051] <= 8'h00;
            reg_file[3052] <= 8'hB3;
            reg_file[3053] <= 8'h86;
            reg_file[3054] <= 8'hF6;
            reg_file[3055] <= 8'h00;
            reg_file[3056] <= 8'hB3;
            reg_file[3057] <= 8'h37;
            reg_file[3058] <= 8'hA6;
            reg_file[3059] <= 8'h00;
            reg_file[3060] <= 8'h33;
            reg_file[3061] <= 8'h87;
            reg_file[3062] <= 8'hF6;
            reg_file[3063] <= 8'h00;
            reg_file[3064] <= 8'h13;
            reg_file[3065] <= 8'h08;
            reg_file[3066] <= 8'h04;
            reg_file[3067] <= 8'h00;
            reg_file[3068] <= 8'h93;
            reg_file[3069] <= 8'h17;
            reg_file[3070] <= 8'h87;
            reg_file[3071] <= 8'h00;
            reg_file[3072] <= 8'h63;
            reg_file[3073] <= 8'hD6;
            reg_file[3074] <= 8'h07;
            reg_file[3075] <= 8'h08;
            reg_file[3076] <= 8'h13;
            reg_file[3077] <= 8'h08;
            reg_file[3078] <= 8'h18;
            reg_file[3079] <= 8'h00;
            reg_file[3080] <= 8'h93;
            reg_file[3081] <= 8'h07;
            reg_file[3082] <= 8'hF0;
            reg_file[3083] <= 8'h7F;
            reg_file[3084] <= 8'h63;
            reg_file[3085] <= 8'h06;
            reg_file[3086] <= 8'hF8;
            reg_file[3087] <= 8'h30;
            reg_file[3088] <= 8'hB7;
            reg_file[3089] <= 8'h07;
            reg_file[3090] <= 8'h80;
            reg_file[3091] <= 8'hFF;
            reg_file[3092] <= 8'h93;
            reg_file[3093] <= 8'h87;
            reg_file[3094] <= 8'hF7;
            reg_file[3095] <= 8'hFF;
            reg_file[3096] <= 8'h13;
            reg_file[3097] <= 8'h55;
            reg_file[3098] <= 8'h16;
            reg_file[3099] <= 8'h00;
            reg_file[3100] <= 8'hB3;
            reg_file[3101] <= 8'h77;
            reg_file[3102] <= 8'hF7;
            reg_file[3103] <= 8'h00;
            reg_file[3104] <= 8'h13;
            reg_file[3105] <= 8'h76;
            reg_file[3106] <= 8'h16;
            reg_file[3107] <= 8'h00;
            reg_file[3108] <= 8'h33;
            reg_file[3109] <= 8'h66;
            reg_file[3110] <= 8'hC5;
            reg_file[3111] <= 8'h00;
            reg_file[3112] <= 8'h13;
            reg_file[3113] <= 8'h95;
            reg_file[3114] <= 8'hF7;
            reg_file[3115] <= 8'h01;
            reg_file[3116] <= 8'h6F;
            reg_file[3117] <= 8'h00;
            reg_file[3118] <= 8'hC0;
            reg_file[3119] <= 8'h26;
            reg_file[3120] <= 8'h93;
            reg_file[3121] <= 8'h85;
            reg_file[3122] <= 8'h06;
            reg_file[3123] <= 8'hFE;
            reg_file[3124] <= 8'h93;
            reg_file[3125] <= 8'h08;
            reg_file[3126] <= 8'h00;
            reg_file[3127] <= 8'h02;
            reg_file[3128] <= 8'hB3;
            reg_file[3129] <= 8'h55;
            reg_file[3130] <= 8'hB7;
            reg_file[3131] <= 8'h00;
            reg_file[3132] <= 8'h13;
            reg_file[3133] <= 8'h08;
            reg_file[3134] <= 8'h00;
            reg_file[3135] <= 8'h00;
            reg_file[3136] <= 8'h63;
            reg_file[3137] <= 8'h88;
            reg_file[3138] <= 8'h16;
            reg_file[3139] <= 8'h01;
            reg_file[3140] <= 8'h13;
            reg_file[3141] <= 8'h08;
            reg_file[3142] <= 8'h00;
            reg_file[3143] <= 8'h04;
            reg_file[3144] <= 8'hB3;
            reg_file[3145] <= 8'h06;
            reg_file[3146] <= 8'hD8;
            reg_file[3147] <= 8'h40;
            reg_file[3148] <= 8'h33;
            reg_file[3149] <= 8'h18;
            reg_file[3150] <= 8'hD7;
            reg_file[3151] <= 8'h00;
            reg_file[3152] <= 8'h33;
            reg_file[3153] <= 8'h66;
            reg_file[3154] <= 8'hC8;
            reg_file[3155] <= 8'h00;
            reg_file[3156] <= 8'h33;
            reg_file[3157] <= 8'h36;
            reg_file[3158] <= 8'hC0;
            reg_file[3159] <= 8'h00;
            reg_file[3160] <= 8'h33;
            reg_file[3161] <= 8'hE6;
            reg_file[3162] <= 8'hC5;
            reg_file[3163] <= 8'h00;
            reg_file[3164] <= 8'h93;
            reg_file[3165] <= 8'h06;
            reg_file[3166] <= 8'h00;
            reg_file[3167] <= 8'h00;
            reg_file[3168] <= 8'h6F;
            reg_file[3169] <= 8'hF0;
            reg_file[3170] <= 8'h9F;
            reg_file[3171] <= 8'hF8;
            reg_file[3172] <= 8'h33;
            reg_file[3173] <= 8'h66;
            reg_file[3174] <= 8'hC7;
            reg_file[3175] <= 8'h00;
            reg_file[3176] <= 8'h33;
            reg_file[3177] <= 8'h36;
            reg_file[3178] <= 8'hC0;
            reg_file[3179] <= 8'h00;
            reg_file[3180] <= 8'h6F;
            reg_file[3181] <= 8'hF0;
            reg_file[3182] <= 8'h1F;
            reg_file[3183] <= 8'hFF;
            reg_file[3184] <= 8'h63;
            reg_file[3185] <= 8'h8C;
            reg_file[3186] <= 8'h06;
            reg_file[3187] <= 8'h12;
            reg_file[3188] <= 8'h33;
            reg_file[3189] <= 8'h88;
            reg_file[3190] <= 8'h88;
            reg_file[3191] <= 8'h40;
            reg_file[3192] <= 8'h63;
            reg_file[3193] <= 8'h14;
            reg_file[3194] <= 8'h04;
            reg_file[3195] <= 8'h06;
            reg_file[3196] <= 8'hB3;
            reg_file[3197] <= 8'hE6;
            reg_file[3198] <= 8'hA7;
            reg_file[3199] <= 8'h00;
            reg_file[3200] <= 8'h63;
            reg_file[3201] <= 8'h9E;
            reg_file[3202] <= 8'h06;
            reg_file[3203] <= 8'h00;
            reg_file[3204] <= 8'h93;
            reg_file[3205] <= 8'h07;
            reg_file[3206] <= 8'hF0;
            reg_file[3207] <= 8'h7F;
            reg_file[3208] <= 8'h63;
            reg_file[3209] <= 8'h0E;
            reg_file[3210] <= 8'hF8;
            reg_file[3211] <= 8'h02;
            reg_file[3212] <= 8'h93;
            reg_file[3213] <= 8'h07;
            reg_file[3214] <= 8'h07;
            reg_file[3215] <= 8'h00;
            reg_file[3216] <= 8'h13;
            reg_file[3217] <= 8'h05;
            reg_file[3218] <= 8'h06;
            reg_file[3219] <= 8'h00;
            reg_file[3220] <= 8'h63;
            reg_file[3221] <= 8'h08;
            reg_file[3222] <= 8'h08;
            reg_file[3223] <= 8'h50;
            reg_file[3224] <= 8'h6F;
            reg_file[3225] <= 8'h00;
            reg_file[3226] <= 8'h80;
            reg_file[3227] <= 8'h20;
            reg_file[3228] <= 8'h93;
            reg_file[3229] <= 8'h05;
            reg_file[3230] <= 8'hF8;
            reg_file[3231] <= 8'hFF;
            reg_file[3232] <= 8'h63;
            reg_file[3233] <= 8'h9E;
            reg_file[3234] <= 8'h05;
            reg_file[3235] <= 8'h00;
            reg_file[3236] <= 8'hB3;
            reg_file[3237] <= 8'h05;
            reg_file[3238] <= 8'hC5;
            reg_file[3239] <= 8'h00;
            reg_file[3240] <= 8'h33;
            reg_file[3241] <= 8'hB6;
            reg_file[3242] <= 8'hC5;
            reg_file[3243] <= 8'h00;
            reg_file[3244] <= 8'hB3;
            reg_file[3245] <= 8'h87;
            reg_file[3246] <= 8'hE7;
            reg_file[3247] <= 8'h00;
            reg_file[3248] <= 8'h33;
            reg_file[3249] <= 8'h87;
            reg_file[3250] <= 8'hC7;
            reg_file[3251] <= 8'h00;
            reg_file[3252] <= 8'h13;
            reg_file[3253] <= 8'h86;
            reg_file[3254] <= 8'h05;
            reg_file[3255] <= 8'h00;
            reg_file[3256] <= 8'h6F;
            reg_file[3257] <= 8'hF0;
            reg_file[3258] <= 8'h1F;
            reg_file[3259] <= 8'hEA;
            reg_file[3260] <= 8'h93;
            reg_file[3261] <= 8'h06;
            reg_file[3262] <= 8'hF0;
            reg_file[3263] <= 8'h7F;
            reg_file[3264] <= 8'h63;
            reg_file[3265] <= 8'h1C;
            reg_file[3266] <= 8'hD8;
            reg_file[3267] <= 8'h04;
            reg_file[3268] <= 8'h33;
            reg_file[3269] <= 8'h65;
            reg_file[3270] <= 8'hC7;
            reg_file[3271] <= 8'h00;
            reg_file[3272] <= 8'h63;
            reg_file[3273] <= 8'h00;
            reg_file[3274] <= 8'h05;
            reg_file[3275] <= 8'h7A;
            reg_file[3276] <= 8'h93;
            reg_file[3277] <= 8'h17;
            reg_file[3278] <= 8'h97;
            reg_file[3279] <= 8'h00;
            reg_file[3280] <= 8'h63;
            reg_file[3281] <= 8'hC0;
            reg_file[3282] <= 8'h07;
            reg_file[3283] <= 8'h7A;
            reg_file[3284] <= 8'h93;
            reg_file[3285] <= 8'h07;
            reg_file[3286] <= 8'h07;
            reg_file[3287] <= 8'h00;
            reg_file[3288] <= 8'h13;
            reg_file[3289] <= 8'h05;
            reg_file[3290] <= 8'h06;
            reg_file[3291] <= 8'h00;
            reg_file[3292] <= 8'h6F;
            reg_file[3293] <= 8'hF0;
            reg_file[3294] <= 8'h1F;
            reg_file[3295] <= 8'hEA;
            reg_file[3296] <= 8'h93;
            reg_file[3297] <= 8'h06;
            reg_file[3298] <= 8'hF0;
            reg_file[3299] <= 8'h7F;
            reg_file[3300] <= 8'h63;
            reg_file[3301] <= 8'h94;
            reg_file[3302] <= 8'hD8;
            reg_file[3303] <= 8'h02;
            reg_file[3304] <= 8'h33;
            reg_file[3305] <= 8'h65;
            reg_file[3306] <= 8'hC7;
            reg_file[3307] <= 8'h00;
            reg_file[3308] <= 8'h63;
            reg_file[3309] <= 8'h08;
            reg_file[3310] <= 8'h05;
            reg_file[3311] <= 8'h72;
            reg_file[3312] <= 8'h93;
            reg_file[3313] <= 8'h17;
            reg_file[3314] <= 8'h97;
            reg_file[3315] <= 8'h00;
            reg_file[3316] <= 8'h63;
            reg_file[3317] <= 8'hCC;
            reg_file[3318] <= 8'h07;
            reg_file[3319] <= 8'h72;
            reg_file[3320] <= 8'h93;
            reg_file[3321] <= 8'h07;
            reg_file[3322] <= 8'h07;
            reg_file[3323] <= 8'h00;
            reg_file[3324] <= 8'h13;
            reg_file[3325] <= 8'h05;
            reg_file[3326] <= 8'h06;
            reg_file[3327] <= 8'h00;
            reg_file[3328] <= 8'h13;
            reg_file[3329] <= 8'h08;
            reg_file[3330] <= 8'hF0;
            reg_file[3331] <= 8'h7F;
            reg_file[3332] <= 8'h13;
            reg_file[3333] <= 8'h04;
            reg_file[3334] <= 8'h00;
            reg_file[3335] <= 8'h00;
            reg_file[3336] <= 8'h6F;
            reg_file[3337] <= 8'hF0;
            reg_file[3338] <= 8'h5F;
            reg_file[3339] <= 8'hE7;
            reg_file[3340] <= 8'hB7;
            reg_file[3341] <= 8'h06;
            reg_file[3342] <= 8'h80;
            reg_file[3343] <= 8'h00;
            reg_file[3344] <= 8'hB3;
            reg_file[3345] <= 8'hE7;
            reg_file[3346] <= 8'hD7;
            reg_file[3347] <= 8'h00;
            reg_file[3348] <= 8'h93;
            reg_file[3349] <= 8'h05;
            reg_file[3350] <= 8'h08;
            reg_file[3351] <= 8'h00;
            reg_file[3352] <= 8'h93;
            reg_file[3353] <= 8'h06;
            reg_file[3354] <= 8'h80;
            reg_file[3355] <= 8'h03;
            reg_file[3356] <= 8'h63;
            reg_file[3357] <= 8'hC0;
            reg_file[3358] <= 8'hB6;
            reg_file[3359] <= 8'h08;
            reg_file[3360] <= 8'h93;
            reg_file[3361] <= 8'h06;
            reg_file[3362] <= 8'hF0;
            reg_file[3363] <= 8'h01;
            reg_file[3364] <= 8'h63;
            reg_file[3365] <= 8'hC2;
            reg_file[3366] <= 8'hB6;
            reg_file[3367] <= 8'h04;
            reg_file[3368] <= 8'h13;
            reg_file[3369] <= 8'h08;
            reg_file[3370] <= 8'h00;
            reg_file[3371] <= 8'h02;
            reg_file[3372] <= 8'h33;
            reg_file[3373] <= 8'h08;
            reg_file[3374] <= 8'hB8;
            reg_file[3375] <= 8'h40;
            reg_file[3376] <= 8'hB3;
            reg_file[3377] <= 8'h96;
            reg_file[3378] <= 8'h07;
            reg_file[3379] <= 8'h01;
            reg_file[3380] <= 8'h33;
            reg_file[3381] <= 8'h53;
            reg_file[3382] <= 8'hB5;
            reg_file[3383] <= 8'h00;
            reg_file[3384] <= 8'h33;
            reg_file[3385] <= 8'h15;
            reg_file[3386] <= 8'h05;
            reg_file[3387] <= 8'h01;
            reg_file[3388] <= 8'hB3;
            reg_file[3389] <= 8'hE6;
            reg_file[3390] <= 8'h66;
            reg_file[3391] <= 8'h00;
            reg_file[3392] <= 8'h33;
            reg_file[3393] <= 8'h35;
            reg_file[3394] <= 8'hA0;
            reg_file[3395] <= 8'h00;
            reg_file[3396] <= 8'h33;
            reg_file[3397] <= 8'hE5;
            reg_file[3398] <= 8'hA6;
            reg_file[3399] <= 8'h00;
            reg_file[3400] <= 8'hB3;
            reg_file[3401] <= 8'hD7;
            reg_file[3402] <= 8'hB7;
            reg_file[3403] <= 8'h00;
            reg_file[3404] <= 8'hB3;
            reg_file[3405] <= 8'h06;
            reg_file[3406] <= 8'hC5;
            reg_file[3407] <= 8'h00;
            reg_file[3408] <= 8'hB3;
            reg_file[3409] <= 8'h87;
            reg_file[3410] <= 8'hE7;
            reg_file[3411] <= 8'h00;
            reg_file[3412] <= 8'h33;
            reg_file[3413] <= 8'hB7;
            reg_file[3414] <= 8'hC6;
            reg_file[3415] <= 8'h00;
            reg_file[3416] <= 8'h33;
            reg_file[3417] <= 8'h87;
            reg_file[3418] <= 8'hE7;
            reg_file[3419] <= 8'h00;
            reg_file[3420] <= 8'h13;
            reg_file[3421] <= 8'h86;
            reg_file[3422] <= 8'h06;
            reg_file[3423] <= 8'h00;
            reg_file[3424] <= 8'h13;
            reg_file[3425] <= 8'h88;
            reg_file[3426] <= 8'h08;
            reg_file[3427] <= 8'h00;
            reg_file[3428] <= 8'h6F;
            reg_file[3429] <= 8'hF0;
            reg_file[3430] <= 8'h9F;
            reg_file[3431] <= 8'hE9;
            reg_file[3432] <= 8'h93;
            reg_file[3433] <= 8'h86;
            reg_file[3434] <= 8'h05;
            reg_file[3435] <= 8'hFE;
            reg_file[3436] <= 8'h13;
            reg_file[3437] <= 8'h03;
            reg_file[3438] <= 8'h00;
            reg_file[3439] <= 8'h02;
            reg_file[3440] <= 8'hB3;
            reg_file[3441] <= 8'hD6;
            reg_file[3442] <= 8'hD7;
            reg_file[3443] <= 8'h00;
            reg_file[3444] <= 8'h13;
            reg_file[3445] <= 8'h08;
            reg_file[3446] <= 8'h00;
            reg_file[3447] <= 8'h00;
            reg_file[3448] <= 8'h63;
            reg_file[3449] <= 8'h88;
            reg_file[3450] <= 8'h65;
            reg_file[3451] <= 8'h00;
            reg_file[3452] <= 8'h13;
            reg_file[3453] <= 8'h08;
            reg_file[3454] <= 8'h00;
            reg_file[3455] <= 8'h04;
            reg_file[3456] <= 8'hB3;
            reg_file[3457] <= 8'h05;
            reg_file[3458] <= 8'hB8;
            reg_file[3459] <= 8'h40;
            reg_file[3460] <= 8'h33;
            reg_file[3461] <= 8'h98;
            reg_file[3462] <= 8'hB7;
            reg_file[3463] <= 8'h00;
            reg_file[3464] <= 8'h33;
            reg_file[3465] <= 8'h65;
            reg_file[3466] <= 8'hA8;
            reg_file[3467] <= 8'h00;
            reg_file[3468] <= 8'h33;
            reg_file[3469] <= 8'h35;
            reg_file[3470] <= 8'hA0;
            reg_file[3471] <= 8'h00;
            reg_file[3472] <= 8'h33;
            reg_file[3473] <= 8'hE5;
            reg_file[3474] <= 8'hA6;
            reg_file[3475] <= 8'h00;
            reg_file[3476] <= 8'h93;
            reg_file[3477] <= 8'h07;
            reg_file[3478] <= 8'h00;
            reg_file[3479] <= 8'h00;
            reg_file[3480] <= 8'h6F;
            reg_file[3481] <= 8'hF0;
            reg_file[3482] <= 8'h5F;
            reg_file[3483] <= 8'hFB;
            reg_file[3484] <= 8'h33;
            reg_file[3485] <= 8'hE5;
            reg_file[3486] <= 8'hA7;
            reg_file[3487] <= 8'h00;
            reg_file[3488] <= 8'h33;
            reg_file[3489] <= 8'h35;
            reg_file[3490] <= 8'hA0;
            reg_file[3491] <= 8'h00;
            reg_file[3492] <= 8'h6F;
            reg_file[3493] <= 8'hF0;
            reg_file[3494] <= 8'h1F;
            reg_file[3495] <= 8'hFF;
            reg_file[3496] <= 8'h13;
            reg_file[3497] <= 8'h08;
            reg_file[3498] <= 8'h14;
            reg_file[3499] <= 8'h00;
            reg_file[3500] <= 8'h93;
            reg_file[3501] <= 8'h76;
            reg_file[3502] <= 8'hE8;
            reg_file[3503] <= 8'h7F;
            reg_file[3504] <= 8'h63;
            reg_file[3505] <= 8'h94;
            reg_file[3506] <= 8'h06;
            reg_file[3507] <= 8'h0C;
            reg_file[3508] <= 8'hB3;
            reg_file[3509] <= 8'hE5;
            reg_file[3510] <= 8'hA7;
            reg_file[3511] <= 8'h00;
            reg_file[3512] <= 8'h63;
            reg_file[3513] <= 8'h1E;
            reg_file[3514] <= 8'h04;
            reg_file[3515] <= 8'h04;
            reg_file[3516] <= 8'h63;
            reg_file[3517] <= 8'h82;
            reg_file[3518] <= 8'h05;
            reg_file[3519] <= 8'h60;
            reg_file[3520] <= 8'hB3;
            reg_file[3521] <= 8'h66;
            reg_file[3522] <= 8'hC7;
            reg_file[3523] <= 8'h00;
            reg_file[3524] <= 8'h63;
            reg_file[3525] <= 8'h80;
            reg_file[3526] <= 8'h06;
            reg_file[3527] <= 8'h3E;
            reg_file[3528] <= 8'h33;
            reg_file[3529] <= 8'h06;
            reg_file[3530] <= 8'hC5;
            reg_file[3531] <= 8'h00;
            reg_file[3532] <= 8'hB3;
            reg_file[3533] <= 8'h87;
            reg_file[3534] <= 8'hE7;
            reg_file[3535] <= 8'h00;
            reg_file[3536] <= 8'h33;
            reg_file[3537] <= 8'h35;
            reg_file[3538] <= 8'hA6;
            reg_file[3539] <= 8'h00;
            reg_file[3540] <= 8'hB3;
            reg_file[3541] <= 8'h87;
            reg_file[3542] <= 8'hA7;
            reg_file[3543] <= 8'h00;
            reg_file[3544] <= 8'h13;
            reg_file[3545] <= 8'h97;
            reg_file[3546] <= 8'h87;
            reg_file[3547] <= 8'h00;
            reg_file[3548] <= 8'h63;
            reg_file[3549] <= 8'h54;
            reg_file[3550] <= 8'h07;
            reg_file[3551] <= 8'h5E;
            reg_file[3552] <= 8'h37;
            reg_file[3553] <= 8'h07;
            reg_file[3554] <= 8'h80;
            reg_file[3555] <= 8'hFF;
            reg_file[3556] <= 8'h13;
            reg_file[3557] <= 8'h07;
            reg_file[3558] <= 8'hF7;
            reg_file[3559] <= 8'hFF;
            reg_file[3560] <= 8'hB3;
            reg_file[3561] <= 8'hF7;
            reg_file[3562] <= 8'hE7;
            reg_file[3563] <= 8'h00;
            reg_file[3564] <= 8'h13;
            reg_file[3565] <= 8'h05;
            reg_file[3566] <= 8'h06;
            reg_file[3567] <= 8'h00;
            reg_file[3568] <= 8'h93;
            reg_file[3569] <= 8'h08;
            reg_file[3570] <= 8'h00;
            reg_file[3571] <= 8'h00;
            reg_file[3572] <= 8'h13;
            reg_file[3573] <= 8'h08;
            reg_file[3574] <= 8'h10;
            reg_file[3575] <= 8'h00;
            reg_file[3576] <= 8'h13;
            reg_file[3577] <= 8'h77;
            reg_file[3578] <= 8'h75;
            reg_file[3579] <= 8'h00;
            reg_file[3580] <= 8'h63;
            reg_file[3581] <= 8'h12;
            reg_file[3582] <= 8'h07;
            reg_file[3583] <= 8'h0E;
            reg_file[3584] <= 8'h63;
            reg_file[3585] <= 8'h06;
            reg_file[3586] <= 8'h04;
            reg_file[3587] <= 8'h74;
            reg_file[3588] <= 8'h13;
            reg_file[3589] <= 8'hF7;
            reg_file[3590] <= 8'h18;
            reg_file[3591] <= 8'h00;
            reg_file[3592] <= 8'h63;
            reg_file[3593] <= 8'h02;
            reg_file[3594] <= 8'h07;
            reg_file[3595] <= 8'h74;
            reg_file[3596] <= 8'h93;
            reg_file[3597] <= 8'hE8;
            reg_file[3598] <= 8'h28;
            reg_file[3599] <= 8'h00;
            reg_file[3600] <= 8'h6F;
            reg_file[3601] <= 8'h00;
            reg_file[3602] <= 8'hC0;
            reg_file[3603] <= 8'h73;
            reg_file[3604] <= 8'h93;
            reg_file[3605] <= 8'h06;
            reg_file[3606] <= 8'hF0;
            reg_file[3607] <= 8'h7F;
            reg_file[3608] <= 8'h63;
            reg_file[3609] <= 8'h16;
            reg_file[3610] <= 8'hD4;
            reg_file[3611] <= 8'h04;
            reg_file[3612] <= 8'h63;
            reg_file[3613] <= 8'h82;
            reg_file[3614] <= 8'h05;
            reg_file[3615] <= 8'h7E;
            reg_file[3616] <= 8'hB7;
            reg_file[3617] <= 8'h06;
            reg_file[3618] <= 8'h40;
            reg_file[3619] <= 8'h00;
            reg_file[3620] <= 8'hB3;
            reg_file[3621] <= 8'hF6;
            reg_file[3622] <= 8'hD7;
            reg_file[3623] <= 8'h00;
            reg_file[3624] <= 8'h93;
            reg_file[3625] <= 8'hB6;
            reg_file[3626] <= 8'h16;
            reg_file[3627] <= 8'h00;
            reg_file[3628] <= 8'h93;
            reg_file[3629] <= 8'h96;
            reg_file[3630] <= 8'h46;
            reg_file[3631] <= 8'h00;
            reg_file[3632] <= 8'h63;
            reg_file[3633] <= 8'h90;
            reg_file[3634] <= 8'h88;
            reg_file[3635] <= 8'h70;
            reg_file[3636] <= 8'h93;
            reg_file[3637] <= 8'h88;
            reg_file[3638] <= 8'h06;
            reg_file[3639] <= 8'h00;
            reg_file[3640] <= 8'hB3;
            reg_file[3641] <= 8'h66;
            reg_file[3642] <= 8'hC7;
            reg_file[3643] <= 8'h00;
            reg_file[3644] <= 8'h63;
            reg_file[3645] <= 8'h88;
            reg_file[3646] <= 8'h06;
            reg_file[3647] <= 8'h00;
            reg_file[3648] <= 8'h93;
            reg_file[3649] <= 8'h16;
            reg_file[3650] <= 8'h97;
            reg_file[3651] <= 8'h00;
            reg_file[3652] <= 8'h63;
            reg_file[3653] <= 8'hC4;
            reg_file[3654] <= 8'h06;
            reg_file[3655] <= 8'h00;
            reg_file[3656] <= 8'h93;
            reg_file[3657] <= 8'h08;
            reg_file[3658] <= 8'h00;
            reg_file[3659] <= 8'h01;
            reg_file[3660] <= 8'h63;
            reg_file[3661] <= 8'h94;
            reg_file[3662] <= 8'h05;
            reg_file[3663] <= 8'h6E;
            reg_file[3664] <= 8'h93;
            reg_file[3665] <= 8'h07;
            reg_file[3666] <= 8'h07;
            reg_file[3667] <= 8'h00;
            reg_file[3668] <= 8'h13;
            reg_file[3669] <= 8'h05;
            reg_file[3670] <= 8'h06;
            reg_file[3671] <= 8'h00;
            reg_file[3672] <= 8'h13;
            reg_file[3673] <= 8'h04;
            reg_file[3674] <= 8'h00;
            reg_file[3675] <= 8'h00;
            reg_file[3676] <= 8'h13;
            reg_file[3677] <= 8'h08;
            reg_file[3678] <= 8'hF0;
            reg_file[3679] <= 8'h7F;
            reg_file[3680] <= 8'h6F;
            reg_file[3681] <= 8'hF0;
            reg_file[3682] <= 8'h9F;
            reg_file[3683] <= 8'hF9;
            reg_file[3684] <= 8'h63;
            reg_file[3685] <= 8'h96;
            reg_file[3686] <= 8'hD8;
            reg_file[3687] <= 8'h00;
            reg_file[3688] <= 8'h93;
            reg_file[3689] <= 8'h08;
            reg_file[3690] <= 8'h00;
            reg_file[3691] <= 8'h00;
            reg_file[3692] <= 8'h6F;
            reg_file[3693] <= 8'hF0;
            reg_file[3694] <= 8'hDF;
            reg_file[3695] <= 8'hFC;
            reg_file[3696] <= 8'h93;
            reg_file[3697] <= 8'h08;
            reg_file[3698] <= 8'h00;
            reg_file[3699] <= 8'h00;
            reg_file[3700] <= 8'h6F;
            reg_file[3701] <= 8'hF0;
            reg_file[3702] <= 8'h9F;
            reg_file[3703] <= 8'hFD;
            reg_file[3704] <= 8'h93;
            reg_file[3705] <= 8'h06;
            reg_file[3706] <= 8'hF0;
            reg_file[3707] <= 8'h7F;
            reg_file[3708] <= 8'h63;
            reg_file[3709] <= 8'h06;
            reg_file[3710] <= 8'hD8;
            reg_file[3711] <= 8'h02;
            reg_file[3712] <= 8'h33;
            reg_file[3713] <= 8'h06;
            reg_file[3714] <= 8'hC5;
            reg_file[3715] <= 8'h00;
            reg_file[3716] <= 8'h33;
            reg_file[3717] <= 8'h35;
            reg_file[3718] <= 8'hA6;
            reg_file[3719] <= 8'h00;
            reg_file[3720] <= 8'hB3;
            reg_file[3721] <= 8'h87;
            reg_file[3722] <= 8'hE7;
            reg_file[3723] <= 8'h00;
            reg_file[3724] <= 8'hB3;
            reg_file[3725] <= 8'h87;
            reg_file[3726] <= 8'hA7;
            reg_file[3727] <= 8'h00;
            reg_file[3728] <= 8'h13;
            reg_file[3729] <= 8'h95;
            reg_file[3730] <= 8'hF7;
            reg_file[3731] <= 8'h01;
            reg_file[3732] <= 8'h13;
            reg_file[3733] <= 8'h56;
            reg_file[3734] <= 8'h16;
            reg_file[3735] <= 8'h00;
            reg_file[3736] <= 8'h33;
            reg_file[3737] <= 8'h65;
            reg_file[3738] <= 8'hC5;
            reg_file[3739] <= 8'h00;
            reg_file[3740] <= 8'h93;
            reg_file[3741] <= 8'hD7;
            reg_file[3742] <= 8'h17;
            reg_file[3743] <= 8'h00;
            reg_file[3744] <= 8'h13;
            reg_file[3745] <= 8'h04;
            reg_file[3746] <= 8'h00;
            reg_file[3747] <= 8'h00;
            reg_file[3748] <= 8'h6F;
            reg_file[3749] <= 8'hF0;
            reg_file[3750] <= 8'h1F;
            reg_file[3751] <= 8'hD0;
            reg_file[3752] <= 8'h63;
            reg_file[3753] <= 8'h88;
            reg_file[3754] <= 8'h09;
            reg_file[3755] <= 8'h00;
            reg_file[3756] <= 8'h93;
            reg_file[3757] <= 8'h07;
            reg_file[3758] <= 8'h30;
            reg_file[3759] <= 8'h00;
            reg_file[3760] <= 8'h63;
            reg_file[3761] <= 8'h98;
            reg_file[3762] <= 8'hF9;
            reg_file[3763] <= 8'h00;
            reg_file[3764] <= 8'h63;
            reg_file[3765] <= 8'h9C;
            reg_file[3766] <= 8'h04;
            reg_file[3767] <= 8'h00;
            reg_file[3768] <= 8'h13;
            reg_file[3769] <= 8'h08;
            reg_file[3770] <= 8'hF0;
            reg_file[3771] <= 8'h7F;
            reg_file[3772] <= 8'h6F;
            reg_file[3773] <= 8'h00;
            reg_file[3774] <= 8'hC0;
            reg_file[3775] <= 8'h06;
            reg_file[3776] <= 8'h93;
            reg_file[3777] <= 8'h07;
            reg_file[3778] <= 8'h20;
            reg_file[3779] <= 8'h00;
            reg_file[3780] <= 8'h63;
            reg_file[3781] <= 8'h94;
            reg_file[3782] <= 8'hF9;
            reg_file[3783] <= 8'h00;
            reg_file[3784] <= 8'hE3;
            reg_file[3785] <= 8'h98;
            reg_file[3786] <= 8'h04;
            reg_file[3787] <= 8'hFE;
            reg_file[3788] <= 8'h13;
            reg_file[3789] <= 8'h04;
            reg_file[3790] <= 8'h00;
            reg_file[3791] <= 8'h00;
            reg_file[3792] <= 8'h93;
            reg_file[3793] <= 8'h07;
            reg_file[3794] <= 8'hF0;
            reg_file[3795] <= 8'hFF;
            reg_file[3796] <= 8'h13;
            reg_file[3797] <= 8'h05;
            reg_file[3798] <= 8'hF0;
            reg_file[3799] <= 8'hFF;
            reg_file[3800] <= 8'h13;
            reg_file[3801] <= 8'h08;
            reg_file[3802] <= 8'hE0;
            reg_file[3803] <= 8'h7F;
            reg_file[3804] <= 8'h93;
            reg_file[3805] <= 8'h08;
            reg_file[3806] <= 8'h50;
            reg_file[3807] <= 8'h00;
            reg_file[3808] <= 8'h13;
            reg_file[3809] <= 8'h07;
            reg_file[3810] <= 8'h20;
            reg_file[3811] <= 8'h00;
            reg_file[3812] <= 8'h93;
            reg_file[3813] <= 8'hE8;
            reg_file[3814] <= 8'h18;
            reg_file[3815] <= 8'h00;
            reg_file[3816] <= 8'h63;
            reg_file[3817] <= 8'h82;
            reg_file[3818] <= 8'hE9;
            reg_file[3819] <= 8'h60;
            reg_file[3820] <= 8'h13;
            reg_file[3821] <= 8'h07;
            reg_file[3822] <= 8'h30;
            reg_file[3823] <= 8'h00;
            reg_file[3824] <= 8'h63;
            reg_file[3825] <= 8'h88;
            reg_file[3826] <= 8'hE9;
            reg_file[3827] <= 8'h5E;
            reg_file[3828] <= 8'h63;
            reg_file[3829] <= 8'h9E;
            reg_file[3830] <= 8'h09;
            reg_file[3831] <= 8'h5E;
            reg_file[3832] <= 8'h13;
            reg_file[3833] <= 8'h77;
            reg_file[3834] <= 8'hF5;
            reg_file[3835] <= 8'h00;
            reg_file[3836] <= 8'h93;
            reg_file[3837] <= 8'h06;
            reg_file[3838] <= 8'h40;
            reg_file[3839] <= 8'h00;
            reg_file[3840] <= 8'h63;
            reg_file[3841] <= 8'h08;
            reg_file[3842] <= 8'hD7;
            reg_file[3843] <= 8'h5E;
            reg_file[3844] <= 8'h13;
            reg_file[3845] <= 8'h07;
            reg_file[3846] <= 8'h45;
            reg_file[3847] <= 8'h00;
            reg_file[3848] <= 8'h33;
            reg_file[3849] <= 8'h35;
            reg_file[3850] <= 8'hA7;
            reg_file[3851] <= 8'h00;
            reg_file[3852] <= 8'hB3;
            reg_file[3853] <= 8'h87;
            reg_file[3854] <= 8'hA7;
            reg_file[3855] <= 8'h00;
            reg_file[3856] <= 8'h13;
            reg_file[3857] <= 8'h05;
            reg_file[3858] <= 8'h07;
            reg_file[3859] <= 8'h00;
            reg_file[3860] <= 8'h6F;
            reg_file[3861] <= 8'h00;
            reg_file[3862] <= 8'hC0;
            reg_file[3863] <= 8'h5D;
            reg_file[3864] <= 8'h63;
            reg_file[3865] <= 8'h88;
            reg_file[3866] <= 8'h09;
            reg_file[3867] <= 8'h00;
            reg_file[3868] <= 8'h93;
            reg_file[3869] <= 8'h07;
            reg_file[3870] <= 8'h30;
            reg_file[3871] <= 8'h00;
            reg_file[3872] <= 8'h63;
            reg_file[3873] <= 8'h9C;
            reg_file[3874] <= 8'hF9;
            reg_file[3875] <= 8'h00;
            reg_file[3876] <= 8'h63;
            reg_file[3877] <= 8'h9C;
            reg_file[3878] <= 8'h04;
            reg_file[3879] <= 8'h50;
            reg_file[3880] <= 8'h93;
            reg_file[3881] <= 8'h07;
            reg_file[3882] <= 8'h00;
            reg_file[3883] <= 8'h00;
            reg_file[3884] <= 8'h13;
            reg_file[3885] <= 8'h05;
            reg_file[3886] <= 8'h00;
            reg_file[3887] <= 8'h00;
            reg_file[3888] <= 8'h93;
            reg_file[3889] <= 8'h08;
            reg_file[3890] <= 8'h50;
            reg_file[3891] <= 8'h00;
            reg_file[3892] <= 8'h6F;
            reg_file[3893] <= 8'h00;
            reg_file[3894] <= 8'h80;
            reg_file[3895] <= 8'h61;
            reg_file[3896] <= 8'h93;
            reg_file[3897] <= 8'h07;
            reg_file[3898] <= 8'h20;
            reg_file[3899] <= 8'h00;
            reg_file[3900] <= 8'h63;
            reg_file[3901] <= 8'h90;
            reg_file[3902] <= 8'hF9;
            reg_file[3903] <= 8'h50;
            reg_file[3904] <= 8'hE3;
            reg_file[3905] <= 8'h94;
            reg_file[3906] <= 8'h04;
            reg_file[3907] <= 8'hFE;
            reg_file[3908] <= 8'h6F;
            reg_file[3909] <= 8'hF0;
            reg_file[3910] <= 8'h9F;
            reg_file[3911] <= 8'hF8;
            reg_file[3912] <= 8'h63;
            reg_file[3913] <= 8'h5A;
            reg_file[3914] <= 8'hD0;
            reg_file[3915] <= 8'h0E;
            reg_file[3916] <= 8'h63;
            reg_file[3917] <= 8'h9E;
            reg_file[3918] <= 8'h08;
            reg_file[3919] <= 8'h08;
            reg_file[3920] <= 8'hB3;
            reg_file[3921] <= 8'h66;
            reg_file[3922] <= 8'hC7;
            reg_file[3923] <= 8'h00;
            reg_file[3924] <= 8'hE3;
            reg_file[3925] <= 8'h80;
            reg_file[3926] <= 8'h06;
            reg_file[3927] <= 8'hBE;
            reg_file[3928] <= 8'h93;
            reg_file[3929] <= 8'h06;
            reg_file[3930] <= 8'hF8;
            reg_file[3931] <= 8'hFF;
            reg_file[3932] <= 8'h63;
            reg_file[3933] <= 8'h9E;
            reg_file[3934] <= 8'h06;
            reg_file[3935] <= 8'h00;
            reg_file[3936] <= 8'h33;
            reg_file[3937] <= 8'h06;
            reg_file[3938] <= 8'hC5;
            reg_file[3939] <= 8'h40;
            reg_file[3940] <= 8'hB3;
            reg_file[3941] <= 8'h87;
            reg_file[3942] <= 8'hE7;
            reg_file[3943] <= 8'h40;
            reg_file[3944] <= 8'hB3;
            reg_file[3945] <= 8'h36;
            reg_file[3946] <= 8'hC5;
            reg_file[3947] <= 8'h00;
            reg_file[3948] <= 8'h33;
            reg_file[3949] <= 8'h87;
            reg_file[3950] <= 8'hD7;
            reg_file[3951] <= 8'h40;
            reg_file[3952] <= 8'h13;
            reg_file[3953] <= 8'h08;
            reg_file[3954] <= 8'h10;
            reg_file[3955] <= 8'h00;
            reg_file[3956] <= 8'h6F;
            reg_file[3957] <= 8'h00;
            reg_file[3958] <= 8'h40;
            reg_file[3959] <= 8'h05;
            reg_file[3960] <= 8'h93;
            reg_file[3961] <= 8'h05;
            reg_file[3962] <= 8'hF0;
            reg_file[3963] <= 8'h7F;
            reg_file[3964] <= 8'hE3;
            reg_file[3965] <= 8'h06;
            reg_file[3966] <= 8'hB8;
            reg_file[3967] <= 8'hBE;
            reg_file[3968] <= 8'h93;
            reg_file[3969] <= 8'h05;
            reg_file[3970] <= 8'h80;
            reg_file[3971] <= 8'h03;
            reg_file[3972] <= 8'h63;
            reg_file[3973] <= 8'hC6;
            reg_file[3974] <= 8'hD5;
            reg_file[3975] <= 8'h0A;
            reg_file[3976] <= 8'h93;
            reg_file[3977] <= 8'h05;
            reg_file[3978] <= 8'hF0;
            reg_file[3979] <= 8'h01;
            reg_file[3980] <= 8'h63;
            reg_file[3981] <= 8'hC8;
            reg_file[3982] <= 8'hD5;
            reg_file[3983] <= 8'h06;
            reg_file[3984] <= 8'h13;
            reg_file[3985] <= 8'h08;
            reg_file[3986] <= 8'h00;
            reg_file[3987] <= 8'h02;
            reg_file[3988] <= 8'h33;
            reg_file[3989] <= 8'h08;
            reg_file[3990] <= 8'hD8;
            reg_file[3991] <= 8'h40;
            reg_file[3992] <= 8'hB3;
            reg_file[3993] <= 8'h58;
            reg_file[3994] <= 8'hD6;
            reg_file[3995] <= 8'h00;
            reg_file[3996] <= 8'hB3;
            reg_file[3997] <= 8'h15;
            reg_file[3998] <= 8'h07;
            reg_file[3999] <= 8'h01;
            reg_file[4000] <= 8'h33;
            reg_file[4001] <= 8'h16;
            reg_file[4002] <= 8'h06;
            reg_file[4003] <= 8'h01;
            reg_file[4004] <= 8'hB3;
            reg_file[4005] <= 8'hE5;
            reg_file[4006] <= 8'h15;
            reg_file[4007] <= 8'h01;
            reg_file[4008] <= 8'h33;
            reg_file[4009] <= 8'h36;
            reg_file[4010] <= 8'hC0;
            reg_file[4011] <= 8'h00;
            reg_file[4012] <= 8'h33;
            reg_file[4013] <= 8'hE6;
            reg_file[4014] <= 8'hC5;
            reg_file[4015] <= 8'h00;
            reg_file[4016] <= 8'hB3;
            reg_file[4017] <= 8'h56;
            reg_file[4018] <= 8'hD7;
            reg_file[4019] <= 8'h00;
            reg_file[4020] <= 8'h33;
            reg_file[4021] <= 8'h06;
            reg_file[4022] <= 8'hC5;
            reg_file[4023] <= 8'h40;
            reg_file[4024] <= 8'hB3;
            reg_file[4025] <= 8'h86;
            reg_file[4026] <= 8'hD7;
            reg_file[4027] <= 8'h40;
            reg_file[4028] <= 8'hB3;
            reg_file[4029] <= 8'h37;
            reg_file[4030] <= 8'hC5;
            reg_file[4031] <= 8'h00;
            reg_file[4032] <= 8'h33;
            reg_file[4033] <= 8'h87;
            reg_file[4034] <= 8'hF6;
            reg_file[4035] <= 8'h40;
            reg_file[4036] <= 8'h13;
            reg_file[4037] <= 8'h08;
            reg_file[4038] <= 8'h04;
            reg_file[4039] <= 8'h00;
            reg_file[4040] <= 8'h93;
            reg_file[4041] <= 8'h17;
            reg_file[4042] <= 8'h87;
            reg_file[4043] <= 8'h00;
            reg_file[4044] <= 8'hE3;
            reg_file[4045] <= 8'hD0;
            reg_file[4046] <= 8'h07;
            reg_file[4047] <= 8'hCC;
            reg_file[4048] <= 8'h37;
            reg_file[4049] <= 8'h09;
            reg_file[4050] <= 8'h80;
            reg_file[4051] <= 8'h00;
            reg_file[4052] <= 8'h13;
            reg_file[4053] <= 8'h09;
            reg_file[4054] <= 8'hF9;
            reg_file[4055] <= 8'hFF;
            reg_file[4056] <= 8'h33;
            reg_file[4057] <= 8'h79;
            reg_file[4058] <= 8'h27;
            reg_file[4059] <= 8'h01;
            reg_file[4060] <= 8'h13;
            reg_file[4061] <= 8'h0A;
            reg_file[4062] <= 8'h06;
            reg_file[4063] <= 8'h00;
            reg_file[4064] <= 8'h13;
            reg_file[4065] <= 8'h04;
            reg_file[4066] <= 8'h08;
            reg_file[4067] <= 8'h00;
            reg_file[4068] <= 8'h6F;
            reg_file[4069] <= 8'h00;
            reg_file[4070] <= 8'h00;
            reg_file[4071] <= 8'h30;
            reg_file[4072] <= 8'h93;
            reg_file[4073] <= 8'h05;
            reg_file[4074] <= 8'hF0;
            reg_file[4075] <= 8'h7F;
            reg_file[4076] <= 8'hE3;
            reg_file[4077] <= 8'h00;
            reg_file[4078] <= 8'hB4;
            reg_file[4079] <= 8'hBA;
            reg_file[4080] <= 8'hB7;
            reg_file[4081] <= 8'h05;
            reg_file[4082] <= 8'h80;
            reg_file[4083] <= 8'h00;
            reg_file[4084] <= 8'h33;
            reg_file[4085] <= 8'h67;
            reg_file[4086] <= 8'hB7;
            reg_file[4087] <= 8'h00;
            reg_file[4088] <= 8'h6F;
            reg_file[4089] <= 8'hF0;
            reg_file[4090] <= 8'h9F;
            reg_file[4091] <= 8'hF8;
            reg_file[4092] <= 8'h93;
            reg_file[4093] <= 8'h85;
            reg_file[4094] <= 8'h06;
            reg_file[4095] <= 8'hFE;
            reg_file[4096] <= 8'h93;
            reg_file[4097] <= 8'h08;
            reg_file[4098] <= 8'h00;
            reg_file[4099] <= 8'h02;
            reg_file[4100] <= 8'hB3;
            reg_file[4101] <= 8'h55;
            reg_file[4102] <= 8'hB7;
            reg_file[4103] <= 8'h00;
            reg_file[4104] <= 8'h13;
            reg_file[4105] <= 8'h08;
            reg_file[4106] <= 8'h00;
            reg_file[4107] <= 8'h00;
            reg_file[4108] <= 8'h63;
            reg_file[4109] <= 8'h88;
            reg_file[4110] <= 8'h16;
            reg_file[4111] <= 8'h01;
            reg_file[4112] <= 8'h13;
            reg_file[4113] <= 8'h08;
            reg_file[4114] <= 8'h00;
            reg_file[4115] <= 8'h04;
            reg_file[4116] <= 8'hB3;
            reg_file[4117] <= 8'h06;
            reg_file[4118] <= 8'hD8;
            reg_file[4119] <= 8'h40;
            reg_file[4120] <= 8'h33;
            reg_file[4121] <= 8'h18;
            reg_file[4122] <= 8'hD7;
            reg_file[4123] <= 8'h00;
            reg_file[4124] <= 8'h33;
            reg_file[4125] <= 8'h66;
            reg_file[4126] <= 8'hC8;
            reg_file[4127] <= 8'h00;
            reg_file[4128] <= 8'h33;
            reg_file[4129] <= 8'h36;
            reg_file[4130] <= 8'hC0;
            reg_file[4131] <= 8'h00;
            reg_file[4132] <= 8'h33;
            reg_file[4133] <= 8'hE6;
            reg_file[4134] <= 8'hC5;
            reg_file[4135] <= 8'h00;
            reg_file[4136] <= 8'h93;
            reg_file[4137] <= 8'h06;
            reg_file[4138] <= 8'h00;
            reg_file[4139] <= 8'h00;
            reg_file[4140] <= 8'h6F;
            reg_file[4141] <= 8'hF0;
            reg_file[4142] <= 8'h9F;
            reg_file[4143] <= 8'hF8;
            reg_file[4144] <= 8'h33;
            reg_file[4145] <= 8'h66;
            reg_file[4146] <= 8'hC7;
            reg_file[4147] <= 8'h00;
            reg_file[4148] <= 8'h33;
            reg_file[4149] <= 8'h36;
            reg_file[4150] <= 8'hC0;
            reg_file[4151] <= 8'h00;
            reg_file[4152] <= 8'h6F;
            reg_file[4153] <= 8'hF0;
            reg_file[4154] <= 8'h1F;
            reg_file[4155] <= 8'hFF;
            reg_file[4156] <= 8'h63;
            reg_file[4157] <= 8'h8C;
            reg_file[4158] <= 8'h06;
            reg_file[4159] <= 8'h12;
            reg_file[4160] <= 8'h33;
            reg_file[4161] <= 8'h88;
            reg_file[4162] <= 8'h88;
            reg_file[4163] <= 8'h40;
            reg_file[4164] <= 8'h63;
            reg_file[4165] <= 8'h12;
            reg_file[4166] <= 8'h04;
            reg_file[4167] <= 8'h06;
            reg_file[4168] <= 8'hB3;
            reg_file[4169] <= 8'hE6;
            reg_file[4170] <= 8'hA7;
            reg_file[4171] <= 8'h00;
            reg_file[4172] <= 8'h63;
            reg_file[4173] <= 8'h98;
            reg_file[4174] <= 8'h06;
            reg_file[4175] <= 8'h00;
            reg_file[4176] <= 8'h93;
            reg_file[4177] <= 8'h07;
            reg_file[4178] <= 8'hF0;
            reg_file[4179] <= 8'h7F;
            reg_file[4180] <= 8'h93;
            reg_file[4181] <= 8'h04;
            reg_file[4182] <= 8'h0E;
            reg_file[4183] <= 8'h00;
            reg_file[4184] <= 8'h6F;
            reg_file[4185] <= 8'hF0;
            reg_file[4186] <= 8'h1F;
            reg_file[4187] <= 8'hC3;
            reg_file[4188] <= 8'h13;
            reg_file[4189] <= 8'h03;
            reg_file[4190] <= 8'hF8;
            reg_file[4191] <= 8'hFF;
            reg_file[4192] <= 8'h63;
            reg_file[4193] <= 8'h10;
            reg_file[4194] <= 8'h03;
            reg_file[4195] <= 8'h02;
            reg_file[4196] <= 8'hB3;
            reg_file[4197] <= 8'h05;
            reg_file[4198] <= 8'hA6;
            reg_file[4199] <= 8'h40;
            reg_file[4200] <= 8'h33;
            reg_file[4201] <= 8'h36;
            reg_file[4202] <= 8'hB6;
            reg_file[4203] <= 8'h00;
            reg_file[4204] <= 8'hB3;
            reg_file[4205] <= 8'h07;
            reg_file[4206] <= 8'hF7;
            reg_file[4207] <= 8'h40;
            reg_file[4208] <= 8'h33;
            reg_file[4209] <= 8'h87;
            reg_file[4210] <= 8'hC7;
            reg_file[4211] <= 8'h40;
            reg_file[4212] <= 8'h93;
            reg_file[4213] <= 8'h04;
            reg_file[4214] <= 8'h0E;
            reg_file[4215] <= 8'h00;
            reg_file[4216] <= 8'h13;
            reg_file[4217] <= 8'h86;
            reg_file[4218] <= 8'h05;
            reg_file[4219] <= 8'h00;
            reg_file[4220] <= 8'h6F;
            reg_file[4221] <= 8'hF0;
            reg_file[4222] <= 8'h5F;
            reg_file[4223] <= 8'hEF;
            reg_file[4224] <= 8'h93;
            reg_file[4225] <= 8'h06;
            reg_file[4226] <= 8'hF0;
            reg_file[4227] <= 8'h7F;
            reg_file[4228] <= 8'h63;
            reg_file[4229] <= 8'h1E;
            reg_file[4230] <= 8'hD8;
            reg_file[4231] <= 8'h04;
            reg_file[4232] <= 8'h33;
            reg_file[4233] <= 8'h65;
            reg_file[4234] <= 8'hC7;
            reg_file[4235] <= 8'h00;
            reg_file[4236] <= 8'h63;
            reg_file[4237] <= 8'h08;
            reg_file[4238] <= 8'h05;
            reg_file[4239] <= 8'h3E;
            reg_file[4240] <= 8'h93;
            reg_file[4241] <= 8'h17;
            reg_file[4242] <= 8'h97;
            reg_file[4243] <= 8'h00;
            reg_file[4244] <= 8'h63;
            reg_file[4245] <= 8'hCA;
            reg_file[4246] <= 8'h07;
            reg_file[4247] <= 8'h3E;
            reg_file[4248] <= 8'h93;
            reg_file[4249] <= 8'h07;
            reg_file[4250] <= 8'h07;
            reg_file[4251] <= 8'h00;
            reg_file[4252] <= 8'h13;
            reg_file[4253] <= 8'h05;
            reg_file[4254] <= 8'h06;
            reg_file[4255] <= 8'h00;
            reg_file[4256] <= 8'h93;
            reg_file[4257] <= 8'h04;
            reg_file[4258] <= 8'h0E;
            reg_file[4259] <= 8'h00;
            reg_file[4260] <= 8'h6F;
            reg_file[4261] <= 8'hF0;
            reg_file[4262] <= 8'h9F;
            reg_file[4263] <= 8'hAD;
            reg_file[4264] <= 8'h93;
            reg_file[4265] <= 8'h06;
            reg_file[4266] <= 8'hF0;
            reg_file[4267] <= 8'h7F;
            reg_file[4268] <= 8'h63;
            reg_file[4269] <= 8'h94;
            reg_file[4270] <= 8'hD8;
            reg_file[4271] <= 8'h02;
            reg_file[4272] <= 8'h33;
            reg_file[4273] <= 8'h65;
            reg_file[4274] <= 8'hC7;
            reg_file[4275] <= 8'h00;
            reg_file[4276] <= 8'h63;
            reg_file[4277] <= 8'h02;
            reg_file[4278] <= 8'h05;
            reg_file[4279] <= 8'h3E;
            reg_file[4280] <= 8'h93;
            reg_file[4281] <= 8'h17;
            reg_file[4282] <= 8'h97;
            reg_file[4283] <= 8'h00;
            reg_file[4284] <= 8'h63;
            reg_file[4285] <= 8'hC4;
            reg_file[4286] <= 8'h07;
            reg_file[4287] <= 8'h3E;
            reg_file[4288] <= 8'h93;
            reg_file[4289] <= 8'h07;
            reg_file[4290] <= 8'h07;
            reg_file[4291] <= 8'h00;
            reg_file[4292] <= 8'h13;
            reg_file[4293] <= 8'h05;
            reg_file[4294] <= 8'h06;
            reg_file[4295] <= 8'h00;
            reg_file[4296] <= 8'h13;
            reg_file[4297] <= 8'h08;
            reg_file[4298] <= 8'hF0;
            reg_file[4299] <= 8'h7F;
            reg_file[4300] <= 8'h93;
            reg_file[4301] <= 8'h04;
            reg_file[4302] <= 8'h0E;
            reg_file[4303] <= 8'h00;
            reg_file[4304] <= 8'h6F;
            reg_file[4305] <= 8'hF0;
            reg_file[4306] <= 8'h5F;
            reg_file[4307] <= 8'hC3;
            reg_file[4308] <= 8'hB7;
            reg_file[4309] <= 8'h06;
            reg_file[4310] <= 8'h80;
            reg_file[4311] <= 8'h00;
            reg_file[4312] <= 8'hB3;
            reg_file[4313] <= 8'hE7;
            reg_file[4314] <= 8'hD7;
            reg_file[4315] <= 8'h00;
            reg_file[4316] <= 8'h13;
            reg_file[4317] <= 8'h03;
            reg_file[4318] <= 8'h08;
            reg_file[4319] <= 8'h00;
            reg_file[4320] <= 8'h93;
            reg_file[4321] <= 8'h06;
            reg_file[4322] <= 8'h80;
            reg_file[4323] <= 8'h03;
            reg_file[4324] <= 8'h63;
            reg_file[4325] <= 8'hC2;
            reg_file[4326] <= 8'h66;
            reg_file[4327] <= 8'h08;
            reg_file[4328] <= 8'h93;
            reg_file[4329] <= 8'h06;
            reg_file[4330] <= 8'hF0;
            reg_file[4331] <= 8'h01;
            reg_file[4332] <= 8'h63;
            reg_file[4333] <= 8'hC4;
            reg_file[4334] <= 8'h66;
            reg_file[4335] <= 8'h04;
            reg_file[4336] <= 8'h93;
            reg_file[4337] <= 8'h06;
            reg_file[4338] <= 8'h00;
            reg_file[4339] <= 8'h02;
            reg_file[4340] <= 8'hB3;
            reg_file[4341] <= 8'h86;
            reg_file[4342] <= 8'h66;
            reg_file[4343] <= 8'h40;
            reg_file[4344] <= 8'hB3;
            reg_file[4345] <= 8'h95;
            reg_file[4346] <= 8'hD7;
            reg_file[4347] <= 8'h00;
            reg_file[4348] <= 8'h33;
            reg_file[4349] <= 8'h58;
            reg_file[4350] <= 8'h65;
            reg_file[4351] <= 8'h00;
            reg_file[4352] <= 8'h33;
            reg_file[4353] <= 8'h15;
            reg_file[4354] <= 8'hD5;
            reg_file[4355] <= 8'h00;
            reg_file[4356] <= 8'hB3;
            reg_file[4357] <= 8'hE5;
            reg_file[4358] <= 8'h05;
            reg_file[4359] <= 8'h01;
            reg_file[4360] <= 8'h33;
            reg_file[4361] <= 8'h35;
            reg_file[4362] <= 8'hA0;
            reg_file[4363] <= 8'h00;
            reg_file[4364] <= 8'h33;
            reg_file[4365] <= 8'hE5;
            reg_file[4366] <= 8'hA5;
            reg_file[4367] <= 8'h00;
            reg_file[4368] <= 8'hB3;
            reg_file[4369] <= 8'hD7;
            reg_file[4370] <= 8'h67;
            reg_file[4371] <= 8'h00;
            reg_file[4372] <= 8'hB3;
            reg_file[4373] <= 8'h05;
            reg_file[4374] <= 8'hA6;
            reg_file[4375] <= 8'h40;
            reg_file[4376] <= 8'hB3;
            reg_file[4377] <= 8'h07;
            reg_file[4378] <= 8'hF7;
            reg_file[4379] <= 8'h40;
            reg_file[4380] <= 8'h33;
            reg_file[4381] <= 8'h37;
            reg_file[4382] <= 8'hB6;
            reg_file[4383] <= 8'h00;
            reg_file[4384] <= 8'h33;
            reg_file[4385] <= 8'h87;
            reg_file[4386] <= 8'hE7;
            reg_file[4387] <= 8'h40;
            reg_file[4388] <= 8'h13;
            reg_file[4389] <= 8'h86;
            reg_file[4390] <= 8'h05;
            reg_file[4391] <= 8'h00;
            reg_file[4392] <= 8'h13;
            reg_file[4393] <= 8'h88;
            reg_file[4394] <= 8'h08;
            reg_file[4395] <= 8'h00;
            reg_file[4396] <= 8'h93;
            reg_file[4397] <= 8'h04;
            reg_file[4398] <= 8'h0E;
            reg_file[4399] <= 8'h00;
            reg_file[4400] <= 8'h6F;
            reg_file[4401] <= 8'hF0;
            reg_file[4402] <= 8'h9F;
            reg_file[4403] <= 8'hE9;
            reg_file[4404] <= 8'h93;
            reg_file[4405] <= 8'h05;
            reg_file[4406] <= 8'h03;
            reg_file[4407] <= 8'hFE;
            reg_file[4408] <= 8'h13;
            reg_file[4409] <= 8'h08;
            reg_file[4410] <= 8'h00;
            reg_file[4411] <= 8'h02;
            reg_file[4412] <= 8'hB3;
            reg_file[4413] <= 8'hD5;
            reg_file[4414] <= 8'hB7;
            reg_file[4415] <= 8'h00;
            reg_file[4416] <= 8'h93;
            reg_file[4417] <= 8'h06;
            reg_file[4418] <= 8'h00;
            reg_file[4419] <= 8'h00;
            reg_file[4420] <= 8'h63;
            reg_file[4421] <= 8'h08;
            reg_file[4422] <= 8'h03;
            reg_file[4423] <= 8'h01;
            reg_file[4424] <= 8'h93;
            reg_file[4425] <= 8'h06;
            reg_file[4426] <= 8'h00;
            reg_file[4427] <= 8'h04;
            reg_file[4428] <= 8'h33;
            reg_file[4429] <= 8'h83;
            reg_file[4430] <= 8'h66;
            reg_file[4431] <= 8'h40;
            reg_file[4432] <= 8'hB3;
            reg_file[4433] <= 8'h96;
            reg_file[4434] <= 8'h67;
            reg_file[4435] <= 8'h00;
            reg_file[4436] <= 8'h33;
            reg_file[4437] <= 8'hE5;
            reg_file[4438] <= 8'hA6;
            reg_file[4439] <= 8'h00;
            reg_file[4440] <= 8'h33;
            reg_file[4441] <= 8'h35;
            reg_file[4442] <= 8'hA0;
            reg_file[4443] <= 8'h00;
            reg_file[4444] <= 8'h33;
            reg_file[4445] <= 8'hE5;
            reg_file[4446] <= 8'hA5;
            reg_file[4447] <= 8'h00;
            reg_file[4448] <= 8'h93;
            reg_file[4449] <= 8'h07;
            reg_file[4450] <= 8'h00;
            reg_file[4451] <= 8'h00;
            reg_file[4452] <= 8'h6F;
            reg_file[4453] <= 8'hF0;
            reg_file[4454] <= 8'h1F;
            reg_file[4455] <= 8'hFB;
            reg_file[4456] <= 8'h33;
            reg_file[4457] <= 8'hE5;
            reg_file[4458] <= 8'hA7;
            reg_file[4459] <= 8'h00;
            reg_file[4460] <= 8'h33;
            reg_file[4461] <= 8'h35;
            reg_file[4462] <= 8'hA0;
            reg_file[4463] <= 8'h00;
            reg_file[4464] <= 8'h6F;
            reg_file[4465] <= 8'hF0;
            reg_file[4466] <= 8'h1F;
            reg_file[4467] <= 8'hFF;
            reg_file[4468] <= 8'h93;
            reg_file[4469] <= 8'h06;
            reg_file[4470] <= 8'h14;
            reg_file[4471] <= 8'h00;
            reg_file[4472] <= 8'h93;
            reg_file[4473] <= 8'hF6;
            reg_file[4474] <= 8'hE6;
            reg_file[4475] <= 8'h7F;
            reg_file[4476] <= 8'h63;
            reg_file[4477] <= 8'h9E;
            reg_file[4478] <= 8'h06;
            reg_file[4479] <= 8'h12;
            reg_file[4480] <= 8'h33;
            reg_file[4481] <= 8'hE8;
            reg_file[4482] <= 8'hA7;
            reg_file[4483] <= 8'h00;
            reg_file[4484] <= 8'hB3;
            reg_file[4485] <= 8'h65;
            reg_file[4486] <= 8'hC7;
            reg_file[4487] <= 8'h00;
            reg_file[4488] <= 8'h63;
            reg_file[4489] <= 8'h18;
            reg_file[4490] <= 8'h04;
            reg_file[4491] <= 8'h0C;
            reg_file[4492] <= 8'h63;
            reg_file[4493] <= 8'h10;
            reg_file[4494] <= 8'h08;
            reg_file[4495] <= 8'h08;
            reg_file[4496] <= 8'h63;
            reg_file[4497] <= 8'h9E;
            reg_file[4498] <= 8'h05;
            reg_file[4499] <= 8'h22;
            reg_file[4500] <= 8'h93;
            reg_file[4501] <= 8'h84;
            reg_file[4502] <= 8'hE9;
            reg_file[4503] <= 8'hFF;
            reg_file[4504] <= 8'h93;
            reg_file[4505] <= 8'hB4;
            reg_file[4506] <= 8'h14;
            reg_file[4507] <= 8'h00;
            reg_file[4508] <= 8'h93;
            reg_file[4509] <= 8'h07;
            reg_file[4510] <= 8'h00;
            reg_file[4511] <= 8'h00;
            reg_file[4512] <= 8'h13;
            reg_file[4513] <= 8'h05;
            reg_file[4514] <= 8'h00;
            reg_file[4515] <= 8'h00;
            reg_file[4516] <= 8'h33;
            reg_file[4517] <= 8'h67;
            reg_file[4518] <= 8'hF5;
            reg_file[4519] <= 8'h00;
            reg_file[4520] <= 8'h63;
            reg_file[4521] <= 8'h04;
            reg_file[4522] <= 8'h07;
            reg_file[4523] <= 8'h32;
            reg_file[4524] <= 8'h13;
            reg_file[4525] <= 8'h57;
            reg_file[4526] <= 8'hF5;
            reg_file[4527] <= 8'h01;
            reg_file[4528] <= 8'h13;
            reg_file[4529] <= 8'h94;
            reg_file[4530] <= 8'h17;
            reg_file[4531] <= 8'h00;
            reg_file[4532] <= 8'h33;
            reg_file[4533] <= 8'h04;
            reg_file[4534] <= 8'hE4;
            reg_file[4535] <= 8'h00;
            reg_file[4536] <= 8'h13;
            reg_file[4537] <= 8'h17;
            reg_file[4538] <= 8'h15;
            reg_file[4539] <= 8'h00;
            reg_file[4540] <= 8'h93;
            reg_file[4541] <= 8'h76;
            reg_file[4542] <= 8'h77;
            reg_file[4543] <= 8'h00;
            reg_file[4544] <= 8'h93;
            reg_file[4545] <= 8'h08;
            reg_file[4546] <= 8'h00;
            reg_file[4547] <= 8'h00;
            reg_file[4548] <= 8'h63;
            reg_file[4549] <= 8'h8A;
            reg_file[4550] <= 8'h06;
            reg_file[4551] <= 8'h02;
            reg_file[4552] <= 8'h93;
            reg_file[4553] <= 8'h06;
            reg_file[4554] <= 8'h20;
            reg_file[4555] <= 8'h00;
            reg_file[4556] <= 8'h63;
            reg_file[4557] <= 8'h8A;
            reg_file[4558] <= 8'hD9;
            reg_file[4559] <= 8'h22;
            reg_file[4560] <= 8'h93;
            reg_file[4561] <= 8'h06;
            reg_file[4562] <= 8'h30;
            reg_file[4563] <= 8'h00;
            reg_file[4564] <= 8'h63;
            reg_file[4565] <= 8'h88;
            reg_file[4566] <= 8'hD9;
            reg_file[4567] <= 8'h20;
            reg_file[4568] <= 8'h93;
            reg_file[4569] <= 8'h08;
            reg_file[4570] <= 8'h10;
            reg_file[4571] <= 8'h00;
            reg_file[4572] <= 8'h63;
            reg_file[4573] <= 8'h9E;
            reg_file[4574] <= 8'h09;
            reg_file[4575] <= 8'h00;
            reg_file[4576] <= 8'h93;
            reg_file[4577] <= 8'h76;
            reg_file[4578] <= 8'hF7;
            reg_file[4579] <= 8'h00;
            reg_file[4580] <= 8'h13;
            reg_file[4581] <= 8'h06;
            reg_file[4582] <= 8'h40;
            reg_file[4583] <= 8'h00;
            reg_file[4584] <= 8'h63;
            reg_file[4585] <= 8'h88;
            reg_file[4586] <= 8'hC6;
            reg_file[4587] <= 8'h00;
            reg_file[4588] <= 8'h13;
            reg_file[4589] <= 8'h37;
            reg_file[4590] <= 8'hC7;
            reg_file[4591] <= 8'hFF;
            reg_file[4592] <= 8'h13;
            reg_file[4593] <= 8'h47;
            reg_file[4594] <= 8'h17;
            reg_file[4595] <= 8'h00;
            reg_file[4596] <= 8'h33;
            reg_file[4597] <= 8'h04;
            reg_file[4598] <= 8'hE4;
            reg_file[4599] <= 8'h00;
            reg_file[4600] <= 8'h13;
            reg_file[4601] <= 8'h54;
            reg_file[4602] <= 8'h84;
            reg_file[4603] <= 8'h01;
            reg_file[4604] <= 8'h13;
            reg_file[4605] <= 8'h44;
            reg_file[4606] <= 8'h14;
            reg_file[4607] <= 8'h00;
            reg_file[4608] <= 8'h13;
            reg_file[4609] <= 8'h74;
            reg_file[4610] <= 8'h14;
            reg_file[4611] <= 8'h00;
            reg_file[4612] <= 8'h13;
            reg_file[4613] <= 8'h08;
            reg_file[4614] <= 8'h00;
            reg_file[4615] <= 8'h00;
            reg_file[4616] <= 8'h6F;
            reg_file[4617] <= 8'hF0;
            reg_file[4618] <= 8'h1F;
            reg_file[4619] <= 8'hBF;
            reg_file[4620] <= 8'hE3;
            reg_file[4621] <= 8'h8C;
            reg_file[4622] <= 8'h05;
            reg_file[4623] <= 8'hF8;
            reg_file[4624] <= 8'hB3;
            reg_file[4625] <= 8'h05;
            reg_file[4626] <= 8'hC5;
            reg_file[4627] <= 8'h40;
            reg_file[4628] <= 8'h33;
            reg_file[4629] <= 8'h38;
            reg_file[4630] <= 8'hB5;
            reg_file[4631] <= 8'h00;
            reg_file[4632] <= 8'hB3;
            reg_file[4633] <= 8'h86;
            reg_file[4634] <= 8'hE7;
            reg_file[4635] <= 8'h40;
            reg_file[4636] <= 8'hB3;
            reg_file[4637] <= 8'h86;
            reg_file[4638] <= 8'h06;
            reg_file[4639] <= 8'h41;
            reg_file[4640] <= 8'h13;
            reg_file[4641] <= 8'h98;
            reg_file[4642] <= 8'h86;
            reg_file[4643] <= 8'h00;
            reg_file[4644] <= 8'h63;
            reg_file[4645] <= 8'h5E;
            reg_file[4646] <= 8'h08;
            reg_file[4647] <= 8'h00;
            reg_file[4648] <= 8'h33;
            reg_file[4649] <= 8'h05;
            reg_file[4650] <= 8'hA6;
            reg_file[4651] <= 8'h40;
            reg_file[4652] <= 8'hB3;
            reg_file[4653] <= 8'h07;
            reg_file[4654] <= 8'hF7;
            reg_file[4655] <= 8'h40;
            reg_file[4656] <= 8'h33;
            reg_file[4657] <= 8'h36;
            reg_file[4658] <= 8'hA6;
            reg_file[4659] <= 8'h00;
            reg_file[4660] <= 8'hB3;
            reg_file[4661] <= 8'h87;
            reg_file[4662] <= 8'hC7;
            reg_file[4663] <= 8'h40;
            reg_file[4664] <= 8'h93;
            reg_file[4665] <= 8'h04;
            reg_file[4666] <= 8'h0E;
            reg_file[4667] <= 8'h00;
            reg_file[4668] <= 8'h6F;
            reg_file[4669] <= 8'hF0;
            reg_file[4670] <= 8'h9F;
            reg_file[4671] <= 8'hF6;
            reg_file[4672] <= 8'h33;
            reg_file[4673] <= 8'hE5;
            reg_file[4674] <= 8'hD5;
            reg_file[4675] <= 8'h00;
            reg_file[4676] <= 8'h63;
            reg_file[4677] <= 8'h1A;
            reg_file[4678] <= 8'h05;
            reg_file[4679] <= 8'h18;
            reg_file[4680] <= 8'h93;
            reg_file[4681] <= 8'h84;
            reg_file[4682] <= 8'hE9;
            reg_file[4683] <= 8'hFF;
            reg_file[4684] <= 8'h93;
            reg_file[4685] <= 8'hB4;
            reg_file[4686] <= 8'h14;
            reg_file[4687] <= 8'h00;
            reg_file[4688] <= 8'h93;
            reg_file[4689] <= 8'h07;
            reg_file[4690] <= 8'h00;
            reg_file[4691] <= 8'h00;
            reg_file[4692] <= 8'h6F;
            reg_file[4693] <= 8'hF0;
            reg_file[4694] <= 8'h1F;
            reg_file[4695] <= 8'hF5;
            reg_file[4696] <= 8'h93;
            reg_file[4697] <= 8'h06;
            reg_file[4698] <= 8'hF0;
            reg_file[4699] <= 8'h7F;
            reg_file[4700] <= 8'h63;
            reg_file[4701] <= 8'h12;
            reg_file[4702] <= 8'hD4;
            reg_file[4703] <= 8'h02;
            reg_file[4704] <= 8'h63;
            reg_file[4705] <= 8'h04;
            reg_file[4706] <= 8'h08;
            reg_file[4707] <= 8'h38;
            reg_file[4708] <= 8'hB7;
            reg_file[4709] <= 8'h06;
            reg_file[4710] <= 8'h40;
            reg_file[4711] <= 8'h00;
            reg_file[4712] <= 8'hB3;
            reg_file[4713] <= 8'hF6;
            reg_file[4714] <= 8'hD7;
            reg_file[4715] <= 8'h00;
            reg_file[4716] <= 8'h93;
            reg_file[4717] <= 8'hB6;
            reg_file[4718] <= 8'h16;
            reg_file[4719] <= 8'h00;
            reg_file[4720] <= 8'h93;
            reg_file[4721] <= 8'h96;
            reg_file[4722] <= 8'h46;
            reg_file[4723] <= 8'h00;
            reg_file[4724] <= 8'h63;
            reg_file[4725] <= 8'h90;
            reg_file[4726] <= 8'h88;
            reg_file[4727] <= 8'h38;
            reg_file[4728] <= 8'h93;
            reg_file[4729] <= 8'h88;
            reg_file[4730] <= 8'h06;
            reg_file[4731] <= 8'h00;
            reg_file[4732] <= 8'h6F;
            reg_file[4733] <= 8'h00;
            reg_file[4734] <= 8'hC0;
            reg_file[4735] <= 8'h00;
            reg_file[4736] <= 8'h63;
            reg_file[4737] <= 8'h98;
            reg_file[4738] <= 8'hD8;
            reg_file[4739] <= 8'h02;
            reg_file[4740] <= 8'h93;
            reg_file[4741] <= 8'h08;
            reg_file[4742] <= 8'h00;
            reg_file[4743] <= 8'h00;
            reg_file[4744] <= 8'h63;
            reg_file[4745] <= 8'h88;
            reg_file[4746] <= 8'h05;
            reg_file[4747] <= 8'h00;
            reg_file[4748] <= 8'h93;
            reg_file[4749] <= 8'h16;
            reg_file[4750] <= 8'h97;
            reg_file[4751] <= 8'h00;
            reg_file[4752] <= 8'h63;
            reg_file[4753] <= 8'hC4;
            reg_file[4754] <= 8'h06;
            reg_file[4755] <= 8'h00;
            reg_file[4756] <= 8'h93;
            reg_file[4757] <= 8'h08;
            reg_file[4758] <= 8'h00;
            reg_file[4759] <= 8'h01;
            reg_file[4760] <= 8'h63;
            reg_file[4761] <= 8'h10;
            reg_file[4762] <= 8'h08;
            reg_file[4763] <= 8'h36;
            reg_file[4764] <= 8'h63;
            reg_file[4765] <= 8'h8E;
            reg_file[4766] <= 8'h05;
            reg_file[4767] <= 8'h20;
            reg_file[4768] <= 8'h93;
            reg_file[4769] <= 8'h07;
            reg_file[4770] <= 8'h07;
            reg_file[4771] <= 8'h00;
            reg_file[4772] <= 8'h13;
            reg_file[4773] <= 8'h05;
            reg_file[4774] <= 8'h06;
            reg_file[4775] <= 8'h00;
            reg_file[4776] <= 8'h93;
            reg_file[4777] <= 8'h04;
            reg_file[4778] <= 8'h0E;
            reg_file[4779] <= 8'h00;
            reg_file[4780] <= 8'h6F;
            reg_file[4781] <= 8'hF0;
            reg_file[4782] <= 8'hDF;
            reg_file[4783] <= 8'hBA;
            reg_file[4784] <= 8'h93;
            reg_file[4785] <= 8'h08;
            reg_file[4786] <= 8'h00;
            reg_file[4787] <= 8'h00;
            reg_file[4788] <= 8'h6F;
            reg_file[4789] <= 8'hF0;
            reg_file[4790] <= 8'h5F;
            reg_file[4791] <= 8'hFE;
            reg_file[4792] <= 8'h33;
            reg_file[4793] <= 8'h0A;
            reg_file[4794] <= 8'hC5;
            reg_file[4795] <= 8'h40;
            reg_file[4796] <= 8'hB3;
            reg_file[4797] <= 8'h36;
            reg_file[4798] <= 8'h45;
            reg_file[4799] <= 8'h01;
            reg_file[4800] <= 8'h33;
            reg_file[4801] <= 8'h89;
            reg_file[4802] <= 8'hE7;
            reg_file[4803] <= 8'h40;
            reg_file[4804] <= 8'h33;
            reg_file[4805] <= 8'h09;
            reg_file[4806] <= 8'hD9;
            reg_file[4807] <= 8'h40;
            reg_file[4808] <= 8'h93;
            reg_file[4809] <= 8'h16;
            reg_file[4810] <= 8'h89;
            reg_file[4811] <= 8'h00;
            reg_file[4812] <= 8'h63;
            reg_file[4813] <= 8'hD2;
            reg_file[4814] <= 8'h06;
            reg_file[4815] <= 8'h08;
            reg_file[4816] <= 8'h33;
            reg_file[4817] <= 8'h0A;
            reg_file[4818] <= 8'hA6;
            reg_file[4819] <= 8'h40;
            reg_file[4820] <= 8'hB3;
            reg_file[4821] <= 8'h07;
            reg_file[4822] <= 8'hF7;
            reg_file[4823] <= 8'h40;
            reg_file[4824] <= 8'h33;
            reg_file[4825] <= 8'h37;
            reg_file[4826] <= 8'h46;
            reg_file[4827] <= 8'h01;
            reg_file[4828] <= 8'h33;
            reg_file[4829] <= 8'h89;
            reg_file[4830] <= 8'hE7;
            reg_file[4831] <= 8'h40;
            reg_file[4832] <= 8'h93;
            reg_file[4833] <= 8'h04;
            reg_file[4834] <= 8'h0E;
            reg_file[4835] <= 8'h00;
            reg_file[4836] <= 8'h63;
            reg_file[4837] <= 8'h0C;
            reg_file[4838] <= 8'h09;
            reg_file[4839] <= 8'h06;
            reg_file[4840] <= 8'h13;
            reg_file[4841] <= 8'h05;
            reg_file[4842] <= 8'h09;
            reg_file[4843] <= 8'h00;
            reg_file[4844] <= 8'hEF;
            reg_file[4845] <= 8'h10;
            reg_file[4846] <= 8'h50;
            reg_file[4847] <= 8'h70;
            reg_file[4848] <= 8'h13;
            reg_file[4849] <= 8'h08;
            reg_file[4850] <= 8'h85;
            reg_file[4851] <= 8'hFF;
            reg_file[4852] <= 8'h93;
            reg_file[4853] <= 8'h07;
            reg_file[4854] <= 8'hF0;
            reg_file[4855] <= 8'h01;
            reg_file[4856] <= 8'h63;
            reg_file[4857] <= 8'hCA;
            reg_file[4858] <= 8'h07;
            reg_file[4859] <= 8'h07;
            reg_file[4860] <= 8'h93;
            reg_file[4861] <= 8'h07;
            reg_file[4862] <= 8'h00;
            reg_file[4863] <= 8'h02;
            reg_file[4864] <= 8'hB3;
            reg_file[4865] <= 8'h87;
            reg_file[4866] <= 8'h07;
            reg_file[4867] <= 8'h41;
            reg_file[4868] <= 8'h33;
            reg_file[4869] <= 8'h17;
            reg_file[4870] <= 8'h09;
            reg_file[4871] <= 8'h01;
            reg_file[4872] <= 8'hB3;
            reg_file[4873] <= 8'h57;
            reg_file[4874] <= 8'hFA;
            reg_file[4875] <= 8'h00;
            reg_file[4876] <= 8'hB3;
            reg_file[4877] <= 8'hE7;
            reg_file[4878] <= 8'hE7;
            reg_file[4879] <= 8'h00;
            reg_file[4880] <= 8'h33;
            reg_file[4881] <= 8'h16;
            reg_file[4882] <= 8'h0A;
            reg_file[4883] <= 8'h01;
            reg_file[4884] <= 8'h63;
            reg_file[4885] <= 8'h4C;
            reg_file[4886] <= 8'h88;
            reg_file[4887] <= 8'h08;
            reg_file[4888] <= 8'h33;
            reg_file[4889] <= 8'h08;
            reg_file[4890] <= 8'h88;
            reg_file[4891] <= 8'h40;
            reg_file[4892] <= 8'h93;
            reg_file[4893] <= 8'h05;
            reg_file[4894] <= 8'h18;
            reg_file[4895] <= 8'h00;
            reg_file[4896] <= 8'h13;
            reg_file[4897] <= 8'h07;
            reg_file[4898] <= 8'hF0;
            reg_file[4899] <= 8'h01;
            reg_file[4900] <= 8'h63;
            reg_file[4901] <= 8'h4C;
            reg_file[4902] <= 8'hB7;
            reg_file[4903] <= 8'h04;
            reg_file[4904] <= 8'h93;
            reg_file[4905] <= 8'h06;
            reg_file[4906] <= 8'h00;
            reg_file[4907] <= 8'h02;
            reg_file[4908] <= 8'hB3;
            reg_file[4909] <= 8'h86;
            reg_file[4910] <= 8'hB6;
            reg_file[4911] <= 8'h40;
            reg_file[4912] <= 8'h33;
            reg_file[4913] <= 8'h95;
            reg_file[4914] <= 8'hD7;
            reg_file[4915] <= 8'h00;
            reg_file[4916] <= 8'h33;
            reg_file[4917] <= 8'h57;
            reg_file[4918] <= 8'hB6;
            reg_file[4919] <= 8'h00;
            reg_file[4920] <= 8'h33;
            reg_file[4921] <= 8'h16;
            reg_file[4922] <= 8'hD6;
            reg_file[4923] <= 8'h00;
            reg_file[4924] <= 8'h33;
            reg_file[4925] <= 8'h65;
            reg_file[4926] <= 8'hE5;
            reg_file[4927] <= 8'h00;
            reg_file[4928] <= 8'h33;
            reg_file[4929] <= 8'h36;
            reg_file[4930] <= 8'hC0;
            reg_file[4931] <= 8'h00;
            reg_file[4932] <= 8'h33;
            reg_file[4933] <= 8'h65;
            reg_file[4934] <= 8'hC5;
            reg_file[4935] <= 8'h00;
            reg_file[4936] <= 8'hB3;
            reg_file[4937] <= 8'hD7;
            reg_file[4938] <= 8'hB7;
            reg_file[4939] <= 8'h00;
            reg_file[4940] <= 8'h6F;
            reg_file[4941] <= 8'hF0;
            reg_file[4942] <= 8'h9F;
            reg_file[4943] <= 8'hE5;
            reg_file[4944] <= 8'h33;
            reg_file[4945] <= 8'h65;
            reg_file[4946] <= 8'h2A;
            reg_file[4947] <= 8'h01;
            reg_file[4948] <= 8'hE3;
            reg_file[4949] <= 8'h18;
            reg_file[4950] <= 8'h05;
            reg_file[4951] <= 8'hF8;
            reg_file[4952] <= 8'h6F;
            reg_file[4953] <= 8'hF0;
            reg_file[4954] <= 8'h1F;
            reg_file[4955] <= 8'hEF;
            reg_file[4956] <= 8'h13;
            reg_file[4957] <= 8'h05;
            reg_file[4958] <= 8'h0A;
            reg_file[4959] <= 8'h00;
            reg_file[4960] <= 8'hEF;
            reg_file[4961] <= 8'h10;
            reg_file[4962] <= 8'h10;
            reg_file[4963] <= 8'h69;
            reg_file[4964] <= 8'h13;
            reg_file[4965] <= 8'h05;
            reg_file[4966] <= 8'h05;
            reg_file[4967] <= 8'h02;
            reg_file[4968] <= 8'h6F;
            reg_file[4969] <= 8'hF0;
            reg_file[4970] <= 8'h9F;
            reg_file[4971] <= 8'hF8;
            reg_file[4972] <= 8'h93;
            reg_file[4973] <= 8'h07;
            reg_file[4974] <= 8'h85;
            reg_file[4975] <= 8'hFD;
            reg_file[4976] <= 8'hB3;
            reg_file[4977] <= 8'h17;
            reg_file[4978] <= 8'hFA;
            reg_file[4979] <= 8'h00;
            reg_file[4980] <= 8'h13;
            reg_file[4981] <= 8'h06;
            reg_file[4982] <= 8'h00;
            reg_file[4983] <= 8'h00;
            reg_file[4984] <= 8'h6F;
            reg_file[4985] <= 8'hF0;
            reg_file[4986] <= 8'hDF;
            reg_file[4987] <= 8'hF9;
            reg_file[4988] <= 8'h13;
            reg_file[4989] <= 8'h08;
            reg_file[4990] <= 8'h18;
            reg_file[4991] <= 8'hFE;
            reg_file[4992] <= 8'h93;
            reg_file[4993] <= 8'h06;
            reg_file[4994] <= 8'h00;
            reg_file[4995] <= 8'h02;
            reg_file[4996] <= 8'h33;
            reg_file[4997] <= 8'hD8;
            reg_file[4998] <= 8'h07;
            reg_file[4999] <= 8'h01;
            reg_file[5000] <= 8'h13;
            reg_file[5001] <= 8'h07;
            reg_file[5002] <= 8'h00;
            reg_file[5003] <= 8'h00;
            reg_file[5004] <= 8'h63;
            reg_file[5005] <= 8'h88;
            reg_file[5006] <= 8'hD5;
            reg_file[5007] <= 8'h00;
            reg_file[5008] <= 8'h13;
            reg_file[5009] <= 8'h07;
            reg_file[5010] <= 8'h00;
            reg_file[5011] <= 8'h04;
            reg_file[5012] <= 8'h33;
            reg_file[5013] <= 8'h07;
            reg_file[5014] <= 8'hB7;
            reg_file[5015] <= 8'h40;
            reg_file[5016] <= 8'h33;
            reg_file[5017] <= 8'h97;
            reg_file[5018] <= 8'hE7;
            reg_file[5019] <= 8'h00;
            reg_file[5020] <= 8'h33;
            reg_file[5021] <= 8'h67;
            reg_file[5022] <= 8'hE6;
            reg_file[5023] <= 8'h00;
            reg_file[5024] <= 8'h33;
            reg_file[5025] <= 8'h35;
            reg_file[5026] <= 8'hE0;
            reg_file[5027] <= 8'h00;
            reg_file[5028] <= 8'h33;
            reg_file[5029] <= 8'h65;
            reg_file[5030] <= 8'hA8;
            reg_file[5031] <= 8'h00;
            reg_file[5032] <= 8'h6F;
            reg_file[5033] <= 8'hF0;
            reg_file[5034] <= 8'h9F;
            reg_file[5035] <= 8'hEA;
            reg_file[5036] <= 8'h37;
            reg_file[5037] <= 8'h07;
            reg_file[5038] <= 8'h80;
            reg_file[5039] <= 8'hFF;
            reg_file[5040] <= 8'h13;
            reg_file[5041] <= 8'h05;
            reg_file[5042] <= 8'hF7;
            reg_file[5043] <= 8'hFF;
            reg_file[5044] <= 8'h33;
            reg_file[5045] <= 8'h08;
            reg_file[5046] <= 8'h04;
            reg_file[5047] <= 8'h41;
            reg_file[5048] <= 8'h33;
            reg_file[5049] <= 8'hF7;
            reg_file[5050] <= 8'hA7;
            reg_file[5051] <= 8'h00;
            reg_file[5052] <= 8'h6F;
            reg_file[5053] <= 8'hF0;
            reg_file[5054] <= 8'h1F;
            reg_file[5055] <= 8'h8D;
            reg_file[5056] <= 8'h93;
            reg_file[5057] <= 8'h07;
            reg_file[5058] <= 8'h07;
            reg_file[5059] <= 8'h00;
            reg_file[5060] <= 8'h13;
            reg_file[5061] <= 8'h05;
            reg_file[5062] <= 8'h06;
            reg_file[5063] <= 8'h00;
            reg_file[5064] <= 8'h6F;
            reg_file[5065] <= 8'hF0;
            reg_file[5066] <= 8'hDF;
            reg_file[5067] <= 8'hDD;
            reg_file[5068] <= 8'h93;
            reg_file[5069] <= 8'h07;
            reg_file[5070] <= 8'h07;
            reg_file[5071] <= 8'h00;
            reg_file[5072] <= 8'h13;
            reg_file[5073] <= 8'h05;
            reg_file[5074] <= 8'h06;
            reg_file[5075] <= 8'h00;
            reg_file[5076] <= 8'h6F;
            reg_file[5077] <= 8'hF0;
            reg_file[5078] <= 8'h5F;
            reg_file[5079] <= 8'hE6;
            reg_file[5080] <= 8'h93;
            reg_file[5081] <= 8'h87;
            reg_file[5082] <= 8'h06;
            reg_file[5083] <= 8'h00;
            reg_file[5084] <= 8'h13;
            reg_file[5085] <= 8'h85;
            reg_file[5086] <= 8'h05;
            reg_file[5087] <= 8'h00;
            reg_file[5088] <= 8'h6F;
            reg_file[5089] <= 8'hF0;
            reg_file[5090] <= 8'h5F;
            reg_file[5091] <= 8'hDC;
            reg_file[5092] <= 8'h93;
            reg_file[5093] <= 8'h88;
            reg_file[5094] <= 8'h04;
            reg_file[5095] <= 8'h00;
            reg_file[5096] <= 8'hE3;
            reg_file[5097] <= 8'h98;
            reg_file[5098] <= 8'h04;
            reg_file[5099] <= 8'hE0;
            reg_file[5100] <= 8'h13;
            reg_file[5101] <= 8'h37;
            reg_file[5102] <= 8'h87;
            reg_file[5103] <= 8'hFF;
            reg_file[5104] <= 8'h13;
            reg_file[5105] <= 8'h47;
            reg_file[5106] <= 8'h17;
            reg_file[5107] <= 8'h00;
            reg_file[5108] <= 8'h33;
            reg_file[5109] <= 8'h04;
            reg_file[5110] <= 8'hE4;
            reg_file[5111] <= 8'h00;
            reg_file[5112] <= 8'h93;
            reg_file[5113] <= 8'h08;
            reg_file[5114] <= 8'h10;
            reg_file[5115] <= 8'h00;
            reg_file[5116] <= 8'h6F;
            reg_file[5117] <= 8'hF0;
            reg_file[5118] <= 8'hDF;
            reg_file[5119] <= 8'hDF;
            reg_file[5120] <= 8'h93;
            reg_file[5121] <= 8'h08;
            reg_file[5122] <= 8'h10;
            reg_file[5123] <= 8'h00;
            reg_file[5124] <= 8'hE3;
            reg_file[5125] <= 8'h8A;
            reg_file[5126] <= 8'h04;
            reg_file[5127] <= 8'hDE;
            reg_file[5128] <= 8'h13;
            reg_file[5129] <= 8'h37;
            reg_file[5130] <= 8'h87;
            reg_file[5131] <= 8'hFF;
            reg_file[5132] <= 8'h13;
            reg_file[5133] <= 8'h47;
            reg_file[5134] <= 8'h17;
            reg_file[5135] <= 8'h00;
            reg_file[5136] <= 8'h33;
            reg_file[5137] <= 8'h04;
            reg_file[5138] <= 8'hE4;
            reg_file[5139] <= 8'h00;
            reg_file[5140] <= 8'h93;
            reg_file[5141] <= 8'h88;
            reg_file[5142] <= 8'h04;
            reg_file[5143] <= 8'h00;
            reg_file[5144] <= 8'h6F;
            reg_file[5145] <= 8'hF0;
            reg_file[5146] <= 8'h1F;
            reg_file[5147] <= 8'hDE;
            reg_file[5148] <= 8'h93;
            reg_file[5149] <= 8'h07;
            reg_file[5150] <= 8'h00;
            reg_file[5151] <= 8'h00;
            reg_file[5152] <= 8'h13;
            reg_file[5153] <= 8'h08;
            reg_file[5154] <= 8'hF0;
            reg_file[5155] <= 8'h7F;
            reg_file[5156] <= 8'h93;
            reg_file[5157] <= 8'h08;
            reg_file[5158] <= 8'h00;
            reg_file[5159] <= 8'h00;
            reg_file[5160] <= 8'h6F;
            reg_file[5161] <= 8'h00;
            reg_file[5162] <= 8'h40;
            reg_file[5163] <= 8'h12;
            reg_file[5164] <= 8'h93;
            reg_file[5165] <= 8'h07;
            reg_file[5166] <= 8'h07;
            reg_file[5167] <= 8'h00;
            reg_file[5168] <= 8'h13;
            reg_file[5169] <= 8'h05;
            reg_file[5170] <= 8'h06;
            reg_file[5171] <= 8'h00;
            reg_file[5172] <= 8'h13;
            reg_file[5173] <= 8'h08;
            reg_file[5174] <= 8'hF0;
            reg_file[5175] <= 8'h7F;
            reg_file[5176] <= 8'h6F;
            reg_file[5177] <= 8'hF0;
            reg_file[5178] <= 8'h9F;
            reg_file[5179] <= 8'hA6;
            reg_file[5180] <= 8'h93;
            reg_file[5181] <= 8'h07;
            reg_file[5182] <= 8'hF0;
            reg_file[5183] <= 8'hFF;
            reg_file[5184] <= 8'h13;
            reg_file[5185] <= 8'h05;
            reg_file[5186] <= 8'hF0;
            reg_file[5187] <= 8'hFF;
            reg_file[5188] <= 8'h13;
            reg_file[5189] <= 8'h08;
            reg_file[5190] <= 8'hE0;
            reg_file[5191] <= 8'h7F;
            reg_file[5192] <= 8'h13;
            reg_file[5193] <= 8'h04;
            reg_file[5194] <= 8'h00;
            reg_file[5195] <= 8'h00;
            reg_file[5196] <= 8'h6F;
            reg_file[5197] <= 8'hF0;
            reg_file[5198] <= 8'h1F;
            reg_file[5199] <= 8'hA9;
            reg_file[5200] <= 8'h93;
            reg_file[5201] <= 8'h07;
            reg_file[5202] <= 8'h00;
            reg_file[5203] <= 8'h00;
            reg_file[5204] <= 8'h13;
            reg_file[5205] <= 8'h05;
            reg_file[5206] <= 8'h00;
            reg_file[5207] <= 8'h00;
            reg_file[5208] <= 8'h6F;
            reg_file[5209] <= 8'h00;
            reg_file[5210] <= 8'h40;
            reg_file[5211] <= 8'h0F;
            reg_file[5212] <= 8'h93;
            reg_file[5213] <= 8'h07;
            reg_file[5214] <= 8'h00;
            reg_file[5215] <= 8'h00;
            reg_file[5216] <= 8'h13;
            reg_file[5217] <= 8'h05;
            reg_file[5218] <= 8'h00;
            reg_file[5219] <= 8'h00;
            reg_file[5220] <= 8'h6F;
            reg_file[5221] <= 8'hF0;
            reg_file[5222] <= 8'hDF;
            reg_file[5223] <= 8'hFB;
            reg_file[5224] <= 8'h93;
            reg_file[5225] <= 8'h07;
            reg_file[5226] <= 8'h00;
            reg_file[5227] <= 8'h00;
            reg_file[5228] <= 8'h6F;
            reg_file[5229] <= 8'hF0;
            reg_file[5230] <= 8'h9F;
            reg_file[5231] <= 8'hFB;
            reg_file[5232] <= 8'h93;
            reg_file[5233] <= 8'h07;
            reg_file[5234] <= 8'h07;
            reg_file[5235] <= 8'h00;
            reg_file[5236] <= 8'h13;
            reg_file[5237] <= 8'h05;
            reg_file[5238] <= 8'h06;
            reg_file[5239] <= 8'h00;
            reg_file[5240] <= 8'h6F;
            reg_file[5241] <= 8'hF0;
            reg_file[5242] <= 8'hCF;
            reg_file[5243] <= 8'hF2;
            reg_file[5244] <= 8'h93;
            reg_file[5245] <= 8'h07;
            reg_file[5246] <= 8'h00;
            reg_file[5247] <= 8'h00;
            reg_file[5248] <= 8'h93;
            reg_file[5249] <= 8'h04;
            reg_file[5250] <= 8'h0E;
            reg_file[5251] <= 8'h00;
            reg_file[5252] <= 8'h6F;
            reg_file[5253] <= 8'hF0;
            reg_file[5254] <= 8'h1F;
            reg_file[5255] <= 8'hFA;
            reg_file[5256] <= 8'h93;
            reg_file[5257] <= 8'h07;
            reg_file[5258] <= 8'h07;
            reg_file[5259] <= 8'h00;
            reg_file[5260] <= 8'h13;
            reg_file[5261] <= 8'h05;
            reg_file[5262] <= 8'h06;
            reg_file[5263] <= 8'h00;
            reg_file[5264] <= 8'h93;
            reg_file[5265] <= 8'h04;
            reg_file[5266] <= 8'h0E;
            reg_file[5267] <= 8'h00;
            reg_file[5268] <= 8'h6F;
            reg_file[5269] <= 8'hF0;
            reg_file[5270] <= 8'h0F;
            reg_file[5271] <= 8'hF1;
            reg_file[5272] <= 8'h93;
            reg_file[5273] <= 8'h07;
            reg_file[5274] <= 8'h00;
            reg_file[5275] <= 8'h00;
            reg_file[5276] <= 8'h13;
            reg_file[5277] <= 8'h08;
            reg_file[5278] <= 8'hF0;
            reg_file[5279] <= 8'h7F;
            reg_file[5280] <= 8'h6F;
            reg_file[5281] <= 8'hF0;
            reg_file[5282] <= 8'h1F;
            reg_file[5283] <= 8'hFE;
            reg_file[5284] <= 8'h93;
            reg_file[5285] <= 8'h07;
            reg_file[5286] <= 8'h07;
            reg_file[5287] <= 8'h00;
            reg_file[5288] <= 8'h13;
            reg_file[5289] <= 8'h05;
            reg_file[5290] <= 8'h06;
            reg_file[5291] <= 8'h00;
            reg_file[5292] <= 8'h13;
            reg_file[5293] <= 8'h08;
            reg_file[5294] <= 8'hF0;
            reg_file[5295] <= 8'h7F;
            reg_file[5296] <= 8'h93;
            reg_file[5297] <= 8'h04;
            reg_file[5298] <= 8'h0E;
            reg_file[5299] <= 8'h00;
            reg_file[5300] <= 8'h6F;
            reg_file[5301] <= 8'hF0;
            reg_file[5302] <= 8'hDF;
            reg_file[5303] <= 8'h9E;
            reg_file[5304] <= 8'h13;
            reg_file[5305] <= 8'h05;
            reg_file[5306] <= 8'h00;
            reg_file[5307] <= 8'h00;
            reg_file[5308] <= 8'h93;
            reg_file[5309] <= 8'h04;
            reg_file[5310] <= 8'h00;
            reg_file[5311] <= 8'h00;
            reg_file[5312] <= 8'hB7;
            reg_file[5313] <= 8'h07;
            reg_file[5314] <= 8'h40;
            reg_file[5315] <= 8'h00;
            reg_file[5316] <= 8'h13;
            reg_file[5317] <= 8'h08;
            reg_file[5318] <= 8'hF0;
            reg_file[5319] <= 8'h7F;
            reg_file[5320] <= 8'h93;
            reg_file[5321] <= 8'h08;
            reg_file[5322] <= 8'h00;
            reg_file[5323] <= 8'h01;
            reg_file[5324] <= 8'h6F;
            reg_file[5325] <= 8'h00;
            reg_file[5326] <= 8'h00;
            reg_file[5327] <= 8'h08;
            reg_file[5328] <= 8'h93;
            reg_file[5329] <= 8'h07;
            reg_file[5330] <= 8'h00;
            reg_file[5331] <= 8'h00;
            reg_file[5332] <= 8'h13;
            reg_file[5333] <= 8'h05;
            reg_file[5334] <= 8'h00;
            reg_file[5335] <= 8'h00;
            reg_file[5336] <= 8'h13;
            reg_file[5337] <= 8'h08;
            reg_file[5338] <= 8'h00;
            reg_file[5339] <= 8'h00;
            reg_file[5340] <= 8'h6F;
            reg_file[5341] <= 8'hF0;
            reg_file[5342] <= 8'h9F;
            reg_file[5343] <= 8'hF4;
            reg_file[5344] <= 8'h63;
            reg_file[5345] <= 8'h98;
            reg_file[5346] <= 8'h04;
            reg_file[5347] <= 8'h00;
            reg_file[5348] <= 8'h13;
            reg_file[5349] <= 8'h07;
            reg_file[5350] <= 8'h85;
            reg_file[5351] <= 8'h00;
            reg_file[5352] <= 8'h6F;
            reg_file[5353] <= 8'hF0;
            reg_file[5354] <= 8'h1F;
            reg_file[5355] <= 8'hA2;
            reg_file[5356] <= 8'hE3;
            reg_file[5357] <= 8'h9C;
            reg_file[5358] <= 8'h04;
            reg_file[5359] <= 8'hFE;
            reg_file[5360] <= 8'hE3;
            reg_file[5361] <= 8'h1E;
            reg_file[5362] <= 8'h04;
            reg_file[5363] <= 8'h90;
            reg_file[5364] <= 8'h6F;
            reg_file[5365] <= 8'h00;
            reg_file[5366] <= 8'h80;
            reg_file[5367] <= 8'h05;
            reg_file[5368] <= 8'h13;
            reg_file[5369] <= 8'h05;
            reg_file[5370] <= 8'h00;
            reg_file[5371] <= 8'h00;
            reg_file[5372] <= 8'h63;
            reg_file[5373] <= 8'h84;
            reg_file[5374] <= 8'h09;
            reg_file[5375] <= 8'h02;
            reg_file[5376] <= 8'h93;
            reg_file[5377] <= 8'h07;
            reg_file[5378] <= 8'h30;
            reg_file[5379] <= 8'h00;
            reg_file[5380] <= 8'h63;
            reg_file[5381] <= 8'h9A;
            reg_file[5382] <= 8'hF9;
            reg_file[5383] <= 8'h00;
            reg_file[5384] <= 8'h63;
            reg_file[5385] <= 8'h8E;
            reg_file[5386] <= 8'h04;
            reg_file[5387] <= 8'h00;
            reg_file[5388] <= 8'h13;
            reg_file[5389] <= 8'h05;
            reg_file[5390] <= 8'hF0;
            reg_file[5391] <= 8'hFF;
            reg_file[5392] <= 8'h13;
            reg_file[5393] <= 8'h08;
            reg_file[5394] <= 8'hE0;
            reg_file[5395] <= 8'h7F;
            reg_file[5396] <= 8'h6F;
            reg_file[5397] <= 8'h00;
            reg_file[5398] <= 8'h00;
            reg_file[5399] <= 8'h01;
            reg_file[5400] <= 8'h93;
            reg_file[5401] <= 8'h07;
            reg_file[5402] <= 8'h20;
            reg_file[5403] <= 8'h00;
            reg_file[5404] <= 8'hE3;
            reg_file[5405] <= 8'h98;
            reg_file[5406] <= 8'hF9;
            reg_file[5407] <= 8'hFE;
            reg_file[5408] <= 8'hE3;
            reg_file[5409] <= 8'h86;
            reg_file[5410] <= 8'h04;
            reg_file[5411] <= 8'hFE;
            reg_file[5412] <= 8'h93;
            reg_file[5413] <= 8'hE8;
            reg_file[5414] <= 8'h58;
            reg_file[5415] <= 8'h00;
            reg_file[5416] <= 8'h93;
            reg_file[5417] <= 8'h07;
            reg_file[5418] <= 8'h05;
            reg_file[5419] <= 8'h00;
            reg_file[5420] <= 8'h6F;
            reg_file[5421] <= 8'h00;
            reg_file[5422] <= 8'h00;
            reg_file[5423] <= 8'h04;
            reg_file[5424] <= 8'h93;
            reg_file[5425] <= 8'h88;
            reg_file[5426] <= 8'h06;
            reg_file[5427] <= 8'h00;
            reg_file[5428] <= 8'h33;
            reg_file[5429] <= 8'h67;
            reg_file[5430] <= 8'hC7;
            reg_file[5431] <= 8'h00;
            reg_file[5432] <= 8'hE3;
            reg_file[5433] <= 8'h00;
            reg_file[5434] <= 8'h07;
            reg_file[5435] <= 8'h92;
            reg_file[5436] <= 8'h93;
            reg_file[5437] <= 8'h04;
            reg_file[5438] <= 8'h00;
            reg_file[5439] <= 8'h00;
            reg_file[5440] <= 8'hB7;
            reg_file[5441] <= 8'h07;
            reg_file[5442] <= 8'h40;
            reg_file[5443] <= 8'h00;
            reg_file[5444] <= 8'h13;
            reg_file[5445] <= 8'h05;
            reg_file[5446] <= 8'h00;
            reg_file[5447] <= 8'h00;
            reg_file[5448] <= 8'h13;
            reg_file[5449] <= 8'h08;
            reg_file[5450] <= 8'hF0;
            reg_file[5451] <= 8'h7F;
            reg_file[5452] <= 8'h13;
            reg_file[5453] <= 8'h97;
            reg_file[5454] <= 8'h87;
            reg_file[5455] <= 8'h00;
            reg_file[5456] <= 8'h63;
            reg_file[5457] <= 8'h5E;
            reg_file[5458] <= 8'h07;
            reg_file[5459] <= 8'h00;
            reg_file[5460] <= 8'h13;
            reg_file[5461] <= 8'h08;
            reg_file[5462] <= 8'h18;
            reg_file[5463] <= 8'h00;
            reg_file[5464] <= 8'h13;
            reg_file[5465] <= 8'h07;
            reg_file[5466] <= 8'hF0;
            reg_file[5467] <= 8'h7F;
            reg_file[5468] <= 8'hE3;
            reg_file[5469] <= 8'h0E;
            reg_file[5470] <= 8'hE8;
            reg_file[5471] <= 8'hF8;
            reg_file[5472] <= 8'h37;
            reg_file[5473] <= 8'h07;
            reg_file[5474] <= 8'h80;
            reg_file[5475] <= 8'hFF;
            reg_file[5476] <= 8'h13;
            reg_file[5477] <= 8'h07;
            reg_file[5478] <= 8'hF7;
            reg_file[5479] <= 8'hFF;
            reg_file[5480] <= 8'hB3;
            reg_file[5481] <= 8'hF7;
            reg_file[5482] <= 8'hE7;
            reg_file[5483] <= 8'h00;
            reg_file[5484] <= 8'h13;
            reg_file[5485] <= 8'h97;
            reg_file[5486] <= 8'hD7;
            reg_file[5487] <= 8'h01;
            reg_file[5488] <= 8'h13;
            reg_file[5489] <= 8'h55;
            reg_file[5490] <= 8'h35;
            reg_file[5491] <= 8'h00;
            reg_file[5492] <= 8'h33;
            reg_file[5493] <= 8'h65;
            reg_file[5494] <= 8'hA7;
            reg_file[5495] <= 8'h00;
            reg_file[5496] <= 8'h13;
            reg_file[5497] <= 8'h07;
            reg_file[5498] <= 8'hF0;
            reg_file[5499] <= 8'h7F;
            reg_file[5500] <= 8'h93;
            reg_file[5501] <= 8'hD7;
            reg_file[5502] <= 8'h37;
            reg_file[5503] <= 8'h00;
            reg_file[5504] <= 8'h63;
            reg_file[5505] <= 8'h1E;
            reg_file[5506] <= 8'hE8;
            reg_file[5507] <= 8'h00;
            reg_file[5508] <= 8'h33;
            reg_file[5509] <= 8'h65;
            reg_file[5510] <= 8'hF5;
            reg_file[5511] <= 8'h00;
            reg_file[5512] <= 8'h93;
            reg_file[5513] <= 8'h07;
            reg_file[5514] <= 8'h00;
            reg_file[5515] <= 8'h00;
            reg_file[5516] <= 8'h63;
            reg_file[5517] <= 8'h08;
            reg_file[5518] <= 8'h05;
            reg_file[5519] <= 8'h00;
            reg_file[5520] <= 8'hB7;
            reg_file[5521] <= 8'h07;
            reg_file[5522] <= 8'h08;
            reg_file[5523] <= 8'h00;
            reg_file[5524] <= 8'h13;
            reg_file[5525] <= 8'h05;
            reg_file[5526] <= 8'h00;
            reg_file[5527] <= 8'h00;
            reg_file[5528] <= 8'h93;
            reg_file[5529] <= 8'h04;
            reg_file[5530] <= 8'h00;
            reg_file[5531] <= 8'h00;
            reg_file[5532] <= 8'h37;
            reg_file[5533] <= 8'h07;
            reg_file[5534] <= 8'hF0;
            reg_file[5535] <= 8'h7F;
            reg_file[5536] <= 8'h13;
            reg_file[5537] <= 8'h18;
            reg_file[5538] <= 8'h48;
            reg_file[5539] <= 8'h01;
            reg_file[5540] <= 8'h93;
            reg_file[5541] <= 8'h97;
            reg_file[5542] <= 8'hC7;
            reg_file[5543] <= 8'h00;
            reg_file[5544] <= 8'h33;
            reg_file[5545] <= 8'h78;
            reg_file[5546] <= 8'hE8;
            reg_file[5547] <= 8'h00;
            reg_file[5548] <= 8'h93;
            reg_file[5549] <= 8'hD7;
            reg_file[5550] <= 8'hC7;
            reg_file[5551] <= 8'h00;
            reg_file[5552] <= 8'hB3;
            reg_file[5553] <= 8'h67;
            reg_file[5554] <= 8'hF8;
            reg_file[5555] <= 8'h00;
            reg_file[5556] <= 8'h93;
            reg_file[5557] <= 8'h94;
            reg_file[5558] <= 8'hF4;
            reg_file[5559] <= 8'h01;
            reg_file[5560] <= 8'h33;
            reg_file[5561] <= 8'hE7;
            reg_file[5562] <= 8'h97;
            reg_file[5563] <= 8'h00;
            reg_file[5564] <= 8'h93;
            reg_file[5565] <= 8'h05;
            reg_file[5566] <= 8'h07;
            reg_file[5567] <= 8'h00;
            reg_file[5568] <= 8'h63;
            reg_file[5569] <= 8'h84;
            reg_file[5570] <= 8'h08;
            reg_file[5571] <= 8'h00;
            reg_file[5572] <= 8'h73;
            reg_file[5573] <= 8'hA0;
            reg_file[5574] <= 8'h18;
            reg_file[5575] <= 8'h00;
            reg_file[5576] <= 8'h83;
            reg_file[5577] <= 8'h20;
            reg_file[5578] <= 8'hC1;
            reg_file[5579] <= 8'h01;
            reg_file[5580] <= 8'h03;
            reg_file[5581] <= 8'h24;
            reg_file[5582] <= 8'h81;
            reg_file[5583] <= 8'h01;
            reg_file[5584] <= 8'h83;
            reg_file[5585] <= 8'h24;
            reg_file[5586] <= 8'h41;
            reg_file[5587] <= 8'h01;
            reg_file[5588] <= 8'h03;
            reg_file[5589] <= 8'h29;
            reg_file[5590] <= 8'h01;
            reg_file[5591] <= 8'h01;
            reg_file[5592] <= 8'h83;
            reg_file[5593] <= 8'h29;
            reg_file[5594] <= 8'hC1;
            reg_file[5595] <= 8'h00;
            reg_file[5596] <= 8'h03;
            reg_file[5597] <= 8'h2A;
            reg_file[5598] <= 8'h81;
            reg_file[5599] <= 8'h00;
            reg_file[5600] <= 8'h13;
            reg_file[5601] <= 8'h01;
            reg_file[5602] <= 8'h01;
            reg_file[5603] <= 8'h02;
            reg_file[5604] <= 8'h67;
            reg_file[5605] <= 8'h80;
            reg_file[5606] <= 8'h00;
            reg_file[5607] <= 8'h00;
            reg_file[5608] <= 8'hE3;
            reg_file[5609] <= 8'h8E;
            reg_file[5610] <= 8'h88;
            reg_file[5611] <= 8'hC8;
            reg_file[5612] <= 8'h93;
            reg_file[5613] <= 8'h08;
            reg_file[5614] <= 8'h00;
            reg_file[5615] <= 8'h00;
            reg_file[5616] <= 8'h6F;
            reg_file[5617] <= 8'hF0;
            reg_file[5618] <= 8'hDF;
            reg_file[5619] <= 8'hCA;
            reg_file[5620] <= 8'h93;
            reg_file[5621] <= 8'h88;
            reg_file[5622] <= 8'h06;
            reg_file[5623] <= 8'h00;
            reg_file[5624] <= 8'hE3;
            reg_file[5625] <= 8'h80;
            reg_file[5626] <= 8'h05;
            reg_file[5627] <= 8'h86;
            reg_file[5628] <= 8'h6F;
            reg_file[5629] <= 8'hF0;
            reg_file[5630] <= 8'h1F;
            reg_file[5631] <= 8'hF4;
            reg_file[5632] <= 8'hE3;
            reg_file[5633] <= 8'h84;
            reg_file[5634] <= 8'h88;
            reg_file[5635] <= 8'h86;
            reg_file[5636] <= 8'h93;
            reg_file[5637] <= 8'h08;
            reg_file[5638] <= 8'h00;
            reg_file[5639] <= 8'h00;
            reg_file[5640] <= 8'h6F;
            reg_file[5641] <= 8'hF0;
            reg_file[5642] <= 8'h9F;
            reg_file[5643] <= 8'h84;
            reg_file[5644] <= 8'h13;
            reg_file[5645] <= 8'h01;
            reg_file[5646] <= 8'h01;
            reg_file[5647] <= 8'hFD;
            reg_file[5648] <= 8'h23;
            reg_file[5649] <= 8'h24;
            reg_file[5650] <= 8'h81;
            reg_file[5651] <= 8'h02;
            reg_file[5652] <= 8'h23;
            reg_file[5653] <= 8'h2A;
            reg_file[5654] <= 8'h51;
            reg_file[5655] <= 8'h01;
            reg_file[5656] <= 8'h23;
            reg_file[5657] <= 8'h24;
            reg_file[5658] <= 8'h81;
            reg_file[5659] <= 8'h01;
            reg_file[5660] <= 8'h23;
            reg_file[5661] <= 8'h26;
            reg_file[5662] <= 8'h11;
            reg_file[5663] <= 8'h02;
            reg_file[5664] <= 8'h23;
            reg_file[5665] <= 8'h22;
            reg_file[5666] <= 8'h91;
            reg_file[5667] <= 8'h02;
            reg_file[5668] <= 8'h23;
            reg_file[5669] <= 8'h20;
            reg_file[5670] <= 8'h21;
            reg_file[5671] <= 8'h03;
            reg_file[5672] <= 8'h23;
            reg_file[5673] <= 8'h2E;
            reg_file[5674] <= 8'h31;
            reg_file[5675] <= 8'h01;
            reg_file[5676] <= 8'h23;
            reg_file[5677] <= 8'h2C;
            reg_file[5678] <= 8'h41;
            reg_file[5679] <= 8'h01;
            reg_file[5680] <= 8'h23;
            reg_file[5681] <= 8'h28;
            reg_file[5682] <= 8'h61;
            reg_file[5683] <= 8'h01;
            reg_file[5684] <= 8'h23;
            reg_file[5685] <= 8'h26;
            reg_file[5686] <= 8'h71;
            reg_file[5687] <= 8'h01;
            reg_file[5688] <= 8'h23;
            reg_file[5689] <= 8'h22;
            reg_file[5690] <= 8'h91;
            reg_file[5691] <= 8'h01;
            reg_file[5692] <= 8'h13;
            reg_file[5693] <= 8'h04;
            reg_file[5694] <= 8'h05;
            reg_file[5695] <= 8'h00;
            reg_file[5696] <= 8'h13;
            reg_file[5697] <= 8'h0C;
            reg_file[5698] <= 8'h06;
            reg_file[5699] <= 8'h00;
            reg_file[5700] <= 8'h93;
            reg_file[5701] <= 8'h8A;
            reg_file[5702] <= 8'h06;
            reg_file[5703] <= 8'h00;
            reg_file[5704] <= 8'h73;
            reg_file[5705] <= 8'h29;
            reg_file[5706] <= 8'h20;
            reg_file[5707] <= 8'h00;
            reg_file[5708] <= 8'h93;
            reg_file[5709] <= 8'hD7;
            reg_file[5710] <= 8'h45;
            reg_file[5711] <= 8'h01;
            reg_file[5712] <= 8'h93;
            reg_file[5713] <= 8'h9B;
            reg_file[5714] <= 8'hC5;
            reg_file[5715] <= 8'h00;
            reg_file[5716] <= 8'h13;
            reg_file[5717] <= 8'h97;
            reg_file[5718] <= 8'h57;
            reg_file[5719] <= 8'h01;
            reg_file[5720] <= 8'h93;
            reg_file[5721] <= 8'hDB;
            reg_file[5722] <= 8'hCB;
            reg_file[5723] <= 8'h00;
            reg_file[5724] <= 8'h13;
            reg_file[5725] <= 8'hDA;
            reg_file[5726] <= 8'hF5;
            reg_file[5727] <= 8'h01;
            reg_file[5728] <= 8'h63;
            reg_file[5729] <= 8'h0C;
            reg_file[5730] <= 8'h07;
            reg_file[5731] <= 8'h02;
            reg_file[5732] <= 8'h13;
            reg_file[5733] <= 8'hFB;
            reg_file[5734] <= 8'hF7;
            reg_file[5735] <= 8'h7F;
            reg_file[5736] <= 8'h93;
            reg_file[5737] <= 8'h07;
            reg_file[5738] <= 8'hF0;
            reg_file[5739] <= 8'h7F;
            reg_file[5740] <= 8'h63;
            reg_file[5741] <= 8'h08;
            reg_file[5742] <= 8'hFB;
            reg_file[5743] <= 8'h08;
            reg_file[5744] <= 8'h13;
            reg_file[5745] <= 8'h57;
            reg_file[5746] <= 8'hD5;
            reg_file[5747] <= 8'h01;
            reg_file[5748] <= 8'h93;
            reg_file[5749] <= 8'h9B;
            reg_file[5750] <= 8'h3B;
            reg_file[5751] <= 8'h00;
            reg_file[5752] <= 8'hB3;
            reg_file[5753] <= 8'h6B;
            reg_file[5754] <= 8'h77;
            reg_file[5755] <= 8'h01;
            reg_file[5756] <= 8'hB7;
            reg_file[5757] <= 8'h07;
            reg_file[5758] <= 8'h80;
            reg_file[5759] <= 8'h00;
            reg_file[5760] <= 8'hB3;
            reg_file[5761] <= 8'hEB;
            reg_file[5762] <= 8'hFB;
            reg_file[5763] <= 8'h00;
            reg_file[5764] <= 8'h93;
            reg_file[5765] <= 8'h19;
            reg_file[5766] <= 8'h35;
            reg_file[5767] <= 8'h00;
            reg_file[5768] <= 8'h13;
            reg_file[5769] <= 8'h0B;
            reg_file[5770] <= 8'h1B;
            reg_file[5771] <= 8'hC0;
            reg_file[5772] <= 8'h93;
            reg_file[5773] <= 8'h0C;
            reg_file[5774] <= 8'h00;
            reg_file[5775] <= 8'h00;
            reg_file[5776] <= 8'h93;
            reg_file[5777] <= 8'h04;
            reg_file[5778] <= 8'h00;
            reg_file[5779] <= 8'h00;
            reg_file[5780] <= 8'h6F;
            reg_file[5781] <= 8'h00;
            reg_file[5782] <= 8'h80;
            reg_file[5783] <= 8'h08;
            reg_file[5784] <= 8'hB3;
            reg_file[5785] <= 8'hE7;
            reg_file[5786] <= 8'hAB;
            reg_file[5787] <= 8'h00;
            reg_file[5788] <= 8'h63;
            reg_file[5789] <= 8'h8E;
            reg_file[5790] <= 8'h07;
            reg_file[5791] <= 8'h0E;
            reg_file[5792] <= 8'h63;
            reg_file[5793] <= 8'h80;
            reg_file[5794] <= 8'h0B;
            reg_file[5795] <= 8'h04;
            reg_file[5796] <= 8'h13;
            reg_file[5797] <= 8'h85;
            reg_file[5798] <= 8'h0B;
            reg_file[5799] <= 8'h00;
            reg_file[5800] <= 8'hEF;
            reg_file[5801] <= 8'h10;
            reg_file[5802] <= 8'h90;
            reg_file[5803] <= 8'h34;
            reg_file[5804] <= 8'h13;
            reg_file[5805] <= 8'h07;
            reg_file[5806] <= 8'h55;
            reg_file[5807] <= 8'hFF;
            reg_file[5808] <= 8'h93;
            reg_file[5809] <= 8'h07;
            reg_file[5810] <= 8'hC0;
            reg_file[5811] <= 8'h01;
            reg_file[5812] <= 8'h63;
            reg_file[5813] <= 8'hCC;
            reg_file[5814] <= 8'hE7;
            reg_file[5815] <= 8'h02;
            reg_file[5816] <= 8'h93;
            reg_file[5817] <= 8'h06;
            reg_file[5818] <= 8'hD0;
            reg_file[5819] <= 8'h01;
            reg_file[5820] <= 8'h93;
            reg_file[5821] <= 8'h09;
            reg_file[5822] <= 8'h85;
            reg_file[5823] <= 8'hFF;
            reg_file[5824] <= 8'hB3;
            reg_file[5825] <= 8'h86;
            reg_file[5826] <= 8'hE6;
            reg_file[5827] <= 8'h40;
            reg_file[5828] <= 8'hB3;
            reg_file[5829] <= 8'h9B;
            reg_file[5830] <= 8'h3B;
            reg_file[5831] <= 8'h01;
            reg_file[5832] <= 8'hB3;
            reg_file[5833] <= 8'h56;
            reg_file[5834] <= 8'hD4;
            reg_file[5835] <= 8'h00;
            reg_file[5836] <= 8'hB3;
            reg_file[5837] <= 8'hEB;
            reg_file[5838] <= 8'h76;
            reg_file[5839] <= 8'h01;
            reg_file[5840] <= 8'hB3;
            reg_file[5841] <= 8'h19;
            reg_file[5842] <= 8'h34;
            reg_file[5843] <= 8'h01;
            reg_file[5844] <= 8'h93;
            reg_file[5845] <= 8'h05;
            reg_file[5846] <= 8'hD0;
            reg_file[5847] <= 8'hC0;
            reg_file[5848] <= 8'h33;
            reg_file[5849] <= 8'h8B;
            reg_file[5850] <= 8'hA5;
            reg_file[5851] <= 8'h40;
            reg_file[5852] <= 8'h6F;
            reg_file[5853] <= 8'hF0;
            reg_file[5854] <= 8'h1F;
            reg_file[5855] <= 8'hFB;
            reg_file[5856] <= 8'hEF;
            reg_file[5857] <= 8'h10;
            reg_file[5858] <= 8'h10;
            reg_file[5859] <= 8'h31;
            reg_file[5860] <= 8'h13;
            reg_file[5861] <= 8'h05;
            reg_file[5862] <= 8'h05;
            reg_file[5863] <= 8'h02;
            reg_file[5864] <= 8'h6F;
            reg_file[5865] <= 8'hF0;
            reg_file[5866] <= 8'h5F;
            reg_file[5867] <= 8'hFC;
            reg_file[5868] <= 8'h93;
            reg_file[5869] <= 8'h0B;
            reg_file[5870] <= 8'h85;
            reg_file[5871] <= 8'hFD;
            reg_file[5872] <= 8'hB3;
            reg_file[5873] <= 8'h1B;
            reg_file[5874] <= 8'h74;
            reg_file[5875] <= 8'h01;
            reg_file[5876] <= 8'h93;
            reg_file[5877] <= 8'h09;
            reg_file[5878] <= 8'h00;
            reg_file[5879] <= 8'h00;
            reg_file[5880] <= 8'h6F;
            reg_file[5881] <= 8'hF0;
            reg_file[5882] <= 8'hDF;
            reg_file[5883] <= 8'hFD;
            reg_file[5884] <= 8'h33;
            reg_file[5885] <= 8'hE4;
            reg_file[5886] <= 8'hAB;
            reg_file[5887] <= 8'h00;
            reg_file[5888] <= 8'h63;
            reg_file[5889] <= 8'h06;
            reg_file[5890] <= 8'h04;
            reg_file[5891] <= 8'h0A;
            reg_file[5892] <= 8'h93;
            reg_file[5893] <= 8'h97;
            reg_file[5894] <= 8'hCB;
            reg_file[5895] <= 8'h00;
            reg_file[5896] <= 8'h93;
            reg_file[5897] <= 8'h09;
            reg_file[5898] <= 8'h05;
            reg_file[5899] <= 8'h00;
            reg_file[5900] <= 8'h13;
            reg_file[5901] <= 8'h0B;
            reg_file[5902] <= 8'hF0;
            reg_file[5903] <= 8'h7F;
            reg_file[5904] <= 8'h93;
            reg_file[5905] <= 8'h0C;
            reg_file[5906] <= 8'h30;
            reg_file[5907] <= 8'h00;
            reg_file[5908] <= 8'h93;
            reg_file[5909] <= 8'h04;
            reg_file[5910] <= 8'h00;
            reg_file[5911] <= 8'h01;
            reg_file[5912] <= 8'hE3;
            reg_file[5913] <= 8'hCC;
            reg_file[5914] <= 8'h07;
            reg_file[5915] <= 8'hF6;
            reg_file[5916] <= 8'h13;
            reg_file[5917] <= 8'hD7;
            reg_file[5918] <= 8'h4A;
            reg_file[5919] <= 8'h01;
            reg_file[5920] <= 8'h13;
            reg_file[5921] <= 8'h95;
            reg_file[5922] <= 8'hCA;
            reg_file[5923] <= 8'h00;
            reg_file[5924] <= 8'h93;
            reg_file[5925] <= 8'h16;
            reg_file[5926] <= 8'h57;
            reg_file[5927] <= 8'h01;
            reg_file[5928] <= 8'h93;
            reg_file[5929] <= 8'h07;
            reg_file[5930] <= 8'h0C;
            reg_file[5931] <= 8'h00;
            reg_file[5932] <= 8'h13;
            reg_file[5933] <= 8'h54;
            reg_file[5934] <= 8'hC5;
            reg_file[5935] <= 8'h00;
            reg_file[5936] <= 8'h93;
            reg_file[5937] <= 8'h75;
            reg_file[5938] <= 8'hF7;
            reg_file[5939] <= 8'h7F;
            reg_file[5940] <= 8'h93;
            reg_file[5941] <= 8'hDA;
            reg_file[5942] <= 8'hFA;
            reg_file[5943] <= 8'h01;
            reg_file[5944] <= 8'h63;
            reg_file[5945] <= 8'h84;
            reg_file[5946] <= 8'h06;
            reg_file[5947] <= 8'h08;
            reg_file[5948] <= 8'h13;
            reg_file[5949] <= 8'h07;
            reg_file[5950] <= 8'hF0;
            reg_file[5951] <= 8'h7F;
            reg_file[5952] <= 8'h63;
            reg_file[5953] <= 8'h86;
            reg_file[5954] <= 8'hE5;
            reg_file[5955] <= 8'h0E;
            reg_file[5956] <= 8'h93;
            reg_file[5957] <= 8'h57;
            reg_file[5958] <= 8'hDC;
            reg_file[5959] <= 8'h01;
            reg_file[5960] <= 8'h13;
            reg_file[5961] <= 8'h15;
            reg_file[5962] <= 8'h34;
            reg_file[5963] <= 8'h00;
            reg_file[5964] <= 8'h33;
            reg_file[5965] <= 8'hE5;
            reg_file[5966] <= 8'hA7;
            reg_file[5967] <= 8'h00;
            reg_file[5968] <= 8'h37;
            reg_file[5969] <= 8'h04;
            reg_file[5970] <= 8'h80;
            reg_file[5971] <= 8'h00;
            reg_file[5972] <= 8'h33;
            reg_file[5973] <= 8'h64;
            reg_file[5974] <= 8'h85;
            reg_file[5975] <= 8'h00;
            reg_file[5976] <= 8'h93;
            reg_file[5977] <= 8'h17;
            reg_file[5978] <= 8'h3C;
            reg_file[5979] <= 8'h00;
            reg_file[5980] <= 8'h13;
            reg_file[5981] <= 8'h85;
            reg_file[5982] <= 8'h15;
            reg_file[5983] <= 8'hC0;
            reg_file[5984] <= 8'h13;
            reg_file[5985] <= 8'h07;
            reg_file[5986] <= 8'h00;
            reg_file[5987] <= 8'h00;
            reg_file[5988] <= 8'h93;
            reg_file[5989] <= 8'h96;
            reg_file[5990] <= 8'h2C;
            reg_file[5991] <= 8'h00;
            reg_file[5992] <= 8'hB3;
            reg_file[5993] <= 8'hE6;
            reg_file[5994] <= 8'hE6;
            reg_file[5995] <= 8'h00;
            reg_file[5996] <= 8'hB3;
            reg_file[5997] <= 8'h05;
            reg_file[5998] <= 8'hAB;
            reg_file[5999] <= 8'h40;
            reg_file[6000] <= 8'h93;
            reg_file[6001] <= 8'h86;
            reg_file[6002] <= 8'hF6;
            reg_file[6003] <= 8'hFF;
            reg_file[6004] <= 8'h13;
            reg_file[6005] <= 8'h05;
            reg_file[6006] <= 8'hE0;
            reg_file[6007] <= 8'h00;
            reg_file[6008] <= 8'h33;
            reg_file[6009] <= 8'h46;
            reg_file[6010] <= 8'h5A;
            reg_file[6011] <= 8'h01;
            reg_file[6012] <= 8'h63;
            reg_file[6013] <= 8'h60;
            reg_file[6014] <= 8'hD5;
            reg_file[6015] <= 8'h10;
            reg_file[6016] <= 8'h37;
            reg_file[6017] <= 8'h35;
            reg_file[6018] <= 8'h00;
            reg_file[6019] <= 8'h80;
            reg_file[6020] <= 8'h93;
            reg_file[6021] <= 8'h96;
            reg_file[6022] <= 8'h26;
            reg_file[6023] <= 8'h00;
            reg_file[6024] <= 8'h13;
            reg_file[6025] <= 8'h05;
            reg_file[6026] <= 8'hC5;
            reg_file[6027] <= 8'h63;
            reg_file[6028] <= 8'hB3;
            reg_file[6029] <= 8'h86;
            reg_file[6030] <= 8'hA6;
            reg_file[6031] <= 8'h00;
            reg_file[6032] <= 8'h83;
            reg_file[6033] <= 8'hA6;
            reg_file[6034] <= 8'h06;
            reg_file[6035] <= 8'h00;
            reg_file[6036] <= 8'h67;
            reg_file[6037] <= 8'h80;
            reg_file[6038] <= 8'h06;
            reg_file[6039] <= 8'h00;
            reg_file[6040] <= 8'h93;
            reg_file[6041] <= 8'h0B;
            reg_file[6042] <= 8'h00;
            reg_file[6043] <= 8'h00;
            reg_file[6044] <= 8'h93;
            reg_file[6045] <= 8'h09;
            reg_file[6046] <= 8'h00;
            reg_file[6047] <= 8'h00;
            reg_file[6048] <= 8'h13;
            reg_file[6049] <= 8'h0B;
            reg_file[6050] <= 8'h00;
            reg_file[6051] <= 8'h00;
            reg_file[6052] <= 8'h93;
            reg_file[6053] <= 8'h0C;
            reg_file[6054] <= 8'h10;
            reg_file[6055] <= 8'h00;
            reg_file[6056] <= 8'h6F;
            reg_file[6057] <= 8'hF0;
            reg_file[6058] <= 8'h9F;
            reg_file[6059] <= 8'hEE;
            reg_file[6060] <= 8'h93;
            reg_file[6061] <= 8'h0B;
            reg_file[6062] <= 8'h00;
            reg_file[6063] <= 8'h00;
            reg_file[6064] <= 8'h93;
            reg_file[6065] <= 8'h09;
            reg_file[6066] <= 8'h00;
            reg_file[6067] <= 8'h00;
            reg_file[6068] <= 8'h13;
            reg_file[6069] <= 8'h0B;
            reg_file[6070] <= 8'hF0;
            reg_file[6071] <= 8'h7F;
            reg_file[6072] <= 8'h93;
            reg_file[6073] <= 8'h0C;
            reg_file[6074] <= 8'h20;
            reg_file[6075] <= 8'h00;
            reg_file[6076] <= 8'h6F;
            reg_file[6077] <= 8'hF0;
            reg_file[6078] <= 8'h5F;
            reg_file[6079] <= 8'hED;
            reg_file[6080] <= 8'hB3;
            reg_file[6081] <= 8'h67;
            reg_file[6082] <= 8'h84;
            reg_file[6083] <= 8'h01;
            reg_file[6084] <= 8'h63;
            reg_file[6085] <= 8'h84;
            reg_file[6086] <= 8'h07;
            reg_file[6087] <= 8'h08;
            reg_file[6088] <= 8'h63;
            reg_file[6089] <= 8'h02;
            reg_file[6090] <= 8'h04;
            reg_file[6091] <= 8'h04;
            reg_file[6092] <= 8'h13;
            reg_file[6093] <= 8'h05;
            reg_file[6094] <= 8'h04;
            reg_file[6095] <= 8'h00;
            reg_file[6096] <= 8'hEF;
            reg_file[6097] <= 8'h10;
            reg_file[6098] <= 8'h10;
            reg_file[6099] <= 8'h22;
            reg_file[6100] <= 8'h93;
            reg_file[6101] <= 8'h05;
            reg_file[6102] <= 8'h05;
            reg_file[6103] <= 8'h00;
            reg_file[6104] <= 8'h93;
            reg_file[6105] <= 8'h86;
            reg_file[6106] <= 8'h55;
            reg_file[6107] <= 8'hFF;
            reg_file[6108] <= 8'h93;
            reg_file[6109] <= 8'h07;
            reg_file[6110] <= 8'hC0;
            reg_file[6111] <= 8'h01;
            reg_file[6112] <= 8'h63;
            reg_file[6113] <= 8'hCE;
            reg_file[6114] <= 8'hD7;
            reg_file[6115] <= 8'h02;
            reg_file[6116] <= 8'h13;
            reg_file[6117] <= 8'h07;
            reg_file[6118] <= 8'hD0;
            reg_file[6119] <= 8'h01;
            reg_file[6120] <= 8'h93;
            reg_file[6121] <= 8'h87;
            reg_file[6122] <= 8'h85;
            reg_file[6123] <= 8'hFF;
            reg_file[6124] <= 8'h33;
            reg_file[6125] <= 8'h07;
            reg_file[6126] <= 8'hD7;
            reg_file[6127] <= 8'h40;
            reg_file[6128] <= 8'h33;
            reg_file[6129] <= 8'h15;
            reg_file[6130] <= 8'hF4;
            reg_file[6131] <= 8'h00;
            reg_file[6132] <= 8'h33;
            reg_file[6133] <= 8'h57;
            reg_file[6134] <= 8'hEC;
            reg_file[6135] <= 8'h00;
            reg_file[6136] <= 8'h33;
            reg_file[6137] <= 8'h64;
            reg_file[6138] <= 8'hA7;
            reg_file[6139] <= 8'h00;
            reg_file[6140] <= 8'hB3;
            reg_file[6141] <= 8'h17;
            reg_file[6142] <= 8'hFC;
            reg_file[6143] <= 8'h00;
            reg_file[6144] <= 8'h13;
            reg_file[6145] <= 8'h07;
            reg_file[6146] <= 8'hD0;
            reg_file[6147] <= 8'hC0;
            reg_file[6148] <= 8'h33;
            reg_file[6149] <= 8'h05;
            reg_file[6150] <= 8'hB7;
            reg_file[6151] <= 8'h40;
            reg_file[6152] <= 8'h6F;
            reg_file[6153] <= 8'hF0;
            reg_file[6154] <= 8'h9F;
            reg_file[6155] <= 8'hF5;
            reg_file[6156] <= 8'h13;
            reg_file[6157] <= 8'h05;
            reg_file[6158] <= 8'h0C;
            reg_file[6159] <= 8'h00;
            reg_file[6160] <= 8'hEF;
            reg_file[6161] <= 8'h10;
            reg_file[6162] <= 8'h10;
            reg_file[6163] <= 8'h1E;
            reg_file[6164] <= 8'h93;
            reg_file[6165] <= 8'h05;
            reg_file[6166] <= 8'h05;
            reg_file[6167] <= 8'h02;
            reg_file[6168] <= 8'h6F;
            reg_file[6169] <= 8'hF0;
            reg_file[6170] <= 8'h1F;
            reg_file[6171] <= 8'hFC;
            reg_file[6172] <= 8'h13;
            reg_file[6173] <= 8'h85;
            reg_file[6174] <= 8'h85;
            reg_file[6175] <= 8'hFD;
            reg_file[6176] <= 8'h33;
            reg_file[6177] <= 8'h14;
            reg_file[6178] <= 8'hAC;
            reg_file[6179] <= 8'h00;
            reg_file[6180] <= 8'h93;
            reg_file[6181] <= 8'h07;
            reg_file[6182] <= 8'h00;
            reg_file[6183] <= 8'h00;
            reg_file[6184] <= 8'h6F;
            reg_file[6185] <= 8'hF0;
            reg_file[6186] <= 8'h9F;
            reg_file[6187] <= 8'hFD;
            reg_file[6188] <= 8'h33;
            reg_file[6189] <= 8'h66;
            reg_file[6190] <= 8'h84;
            reg_file[6191] <= 8'h01;
            reg_file[6192] <= 8'h63;
            reg_file[6193] <= 8'h08;
            reg_file[6194] <= 8'h06;
            reg_file[6195] <= 8'h02;
            reg_file[6196] <= 8'h13;
            reg_file[6197] <= 8'h17;
            reg_file[6198] <= 8'hC4;
            reg_file[6199] <= 8'h00;
            reg_file[6200] <= 8'h13;
            reg_file[6201] <= 8'h05;
            reg_file[6202] <= 8'hF0;
            reg_file[6203] <= 8'h7F;
            reg_file[6204] <= 8'h63;
            reg_file[6205] <= 8'h4C;
            reg_file[6206] <= 8'h07;
            reg_file[6207] <= 8'h02;
            reg_file[6208] <= 8'h13;
            reg_file[6209] <= 8'h07;
            reg_file[6210] <= 8'h30;
            reg_file[6211] <= 8'h00;
            reg_file[6212] <= 8'h93;
            reg_file[6213] <= 8'h04;
            reg_file[6214] <= 8'h00;
            reg_file[6215] <= 8'h01;
            reg_file[6216] <= 8'h6F;
            reg_file[6217] <= 8'hF0;
            reg_file[6218] <= 8'hDF;
            reg_file[6219] <= 8'hF1;
            reg_file[6220] <= 8'h13;
            reg_file[6221] <= 8'h04;
            reg_file[6222] <= 8'h00;
            reg_file[6223] <= 8'h00;
            reg_file[6224] <= 8'h93;
            reg_file[6225] <= 8'h07;
            reg_file[6226] <= 8'h00;
            reg_file[6227] <= 8'h00;
            reg_file[6228] <= 8'h13;
            reg_file[6229] <= 8'h05;
            reg_file[6230] <= 8'h00;
            reg_file[6231] <= 8'h00;
            reg_file[6232] <= 8'h13;
            reg_file[6233] <= 8'h07;
            reg_file[6234] <= 8'h10;
            reg_file[6235] <= 8'h00;
            reg_file[6236] <= 8'h6F;
            reg_file[6237] <= 8'hF0;
            reg_file[6238] <= 8'h9F;
            reg_file[6239] <= 8'hF0;
            reg_file[6240] <= 8'h13;
            reg_file[6241] <= 8'h04;
            reg_file[6242] <= 8'h00;
            reg_file[6243] <= 8'h00;
            reg_file[6244] <= 8'h93;
            reg_file[6245] <= 8'h07;
            reg_file[6246] <= 8'h00;
            reg_file[6247] <= 8'h00;
            reg_file[6248] <= 8'h13;
            reg_file[6249] <= 8'h05;
            reg_file[6250] <= 8'hF0;
            reg_file[6251] <= 8'h7F;
            reg_file[6252] <= 8'h13;
            reg_file[6253] <= 8'h07;
            reg_file[6254] <= 8'h20;
            reg_file[6255] <= 8'h00;
            reg_file[6256] <= 8'h6F;
            reg_file[6257] <= 8'hF0;
            reg_file[6258] <= 8'h5F;
            reg_file[6259] <= 8'hEF;
            reg_file[6260] <= 8'h13;
            reg_file[6261] <= 8'h07;
            reg_file[6262] <= 8'h30;
            reg_file[6263] <= 8'h00;
            reg_file[6264] <= 8'h6F;
            reg_file[6265] <= 8'hF0;
            reg_file[6266] <= 8'hDF;
            reg_file[6267] <= 8'hEE;
            reg_file[6268] <= 8'h63;
            reg_file[6269] <= 8'h66;
            reg_file[6270] <= 8'h74;
            reg_file[6271] <= 8'h01;
            reg_file[6272] <= 8'h63;
            reg_file[6273] <= 8'h96;
            reg_file[6274] <= 8'h8B;
            reg_file[6275] <= 8'h2E;
            reg_file[6276] <= 8'h63;
            reg_file[6277] <= 8'hE4;
            reg_file[6278] <= 8'hF9;
            reg_file[6279] <= 8'h2E;
            reg_file[6280] <= 8'h13;
            reg_file[6281] <= 8'h95;
            reg_file[6282] <= 8'hFB;
            reg_file[6283] <= 8'h01;
            reg_file[6284] <= 8'h13;
            reg_file[6285] <= 8'hD7;
            reg_file[6286] <= 8'h19;
            reg_file[6287] <= 8'h00;
            reg_file[6288] <= 8'h93;
            reg_file[6289] <= 8'h96;
            reg_file[6290] <= 8'hF9;
            reg_file[6291] <= 8'h01;
            reg_file[6292] <= 8'h93;
            reg_file[6293] <= 8'hDB;
            reg_file[6294] <= 8'h1B;
            reg_file[6295] <= 8'h00;
            reg_file[6296] <= 8'hB3;
            reg_file[6297] <= 8'h69;
            reg_file[6298] <= 8'hE5;
            reg_file[6299] <= 8'h00;
            reg_file[6300] <= 8'h13;
            reg_file[6301] <= 8'h15;
            reg_file[6302] <= 8'h84;
            reg_file[6303] <= 8'h00;
            reg_file[6304] <= 8'h13;
            reg_file[6305] <= 8'hD8;
            reg_file[6306] <= 8'h87;
            reg_file[6307] <= 8'h01;
            reg_file[6308] <= 8'h33;
            reg_file[6309] <= 8'h68;
            reg_file[6310] <= 8'hA8;
            reg_file[6311] <= 8'h00;
            reg_file[6312] <= 8'h13;
            reg_file[6313] <= 8'h55;
            reg_file[6314] <= 8'h05;
            reg_file[6315] <= 8'h01;
            reg_file[6316] <= 8'h33;
            reg_file[6317] <= 8'hD3;
            reg_file[6318] <= 8'hAB;
            reg_file[6319] <= 8'h02;
            reg_file[6320] <= 8'h13;
            reg_file[6321] <= 8'h1E;
            reg_file[6322] <= 8'h08;
            reg_file[6323] <= 8'h01;
            reg_file[6324] <= 8'h13;
            reg_file[6325] <= 8'h5E;
            reg_file[6326] <= 8'h0E;
            reg_file[6327] <= 8'h01;
            reg_file[6328] <= 8'h93;
            reg_file[6329] <= 8'h98;
            reg_file[6330] <= 8'h87;
            reg_file[6331] <= 8'h00;
            reg_file[6332] <= 8'h93;
            reg_file[6333] <= 8'hD7;
            reg_file[6334] <= 8'h09;
            reg_file[6335] <= 8'h01;
            reg_file[6336] <= 8'hB3;
            reg_file[6337] <= 8'hFB;
            reg_file[6338] <= 8'hAB;
            reg_file[6339] <= 8'h02;
            reg_file[6340] <= 8'h93;
            reg_file[6341] <= 8'h0F;
            reg_file[6342] <= 8'h03;
            reg_file[6343] <= 8'h00;
            reg_file[6344] <= 8'h33;
            reg_file[6345] <= 8'h07;
            reg_file[6346] <= 8'h6E;
            reg_file[6347] <= 8'h02;
            reg_file[6348] <= 8'h93;
            reg_file[6349] <= 8'h9B;
            reg_file[6350] <= 8'h0B;
            reg_file[6351] <= 8'h01;
            reg_file[6352] <= 8'hB3;
            reg_file[6353] <= 8'hE7;
            reg_file[6354] <= 8'h77;
            reg_file[6355] <= 8'h01;
            reg_file[6356] <= 8'h63;
            reg_file[6357] <= 8'hFE;
            reg_file[6358] <= 8'hE7;
            reg_file[6359] <= 8'h00;
            reg_file[6360] <= 8'hB3;
            reg_file[6361] <= 8'h87;
            reg_file[6362] <= 8'h07;
            reg_file[6363] <= 8'h01;
            reg_file[6364] <= 8'h93;
            reg_file[6365] <= 8'h0F;
            reg_file[6366] <= 8'hF3;
            reg_file[6367] <= 8'hFF;
            reg_file[6368] <= 8'h63;
            reg_file[6369] <= 8'hE8;
            reg_file[6370] <= 8'h07;
            reg_file[6371] <= 8'h01;
            reg_file[6372] <= 8'h63;
            reg_file[6373] <= 8'hF6;
            reg_file[6374] <= 8'hE7;
            reg_file[6375] <= 8'h00;
            reg_file[6376] <= 8'h93;
            reg_file[6377] <= 8'h0F;
            reg_file[6378] <= 8'hE3;
            reg_file[6379] <= 8'hFF;
            reg_file[6380] <= 8'hB3;
            reg_file[6381] <= 8'h87;
            reg_file[6382] <= 8'h07;
            reg_file[6383] <= 8'h01;
            reg_file[6384] <= 8'hB3;
            reg_file[6385] <= 8'h87;
            reg_file[6386] <= 8'hE7;
            reg_file[6387] <= 8'h40;
            reg_file[6388] <= 8'hB3;
            reg_file[6389] <= 8'hDE;
            reg_file[6390] <= 8'hA7;
            reg_file[6391] <= 8'h02;
            reg_file[6392] <= 8'h93;
            reg_file[6393] <= 8'h99;
            reg_file[6394] <= 8'h09;
            reg_file[6395] <= 8'h01;
            reg_file[6396] <= 8'h93;
            reg_file[6397] <= 8'hD9;
            reg_file[6398] <= 8'h09;
            reg_file[6399] <= 8'h01;
            reg_file[6400] <= 8'hB3;
            reg_file[6401] <= 8'hF7;
            reg_file[6402] <= 8'hA7;
            reg_file[6403] <= 8'h02;
            reg_file[6404] <= 8'h13;
            reg_file[6405] <= 8'h83;
            reg_file[6406] <= 8'h0E;
            reg_file[6407] <= 8'h00;
            reg_file[6408] <= 8'h33;
            reg_file[6409] <= 8'h07;
            reg_file[6410] <= 8'hDE;
            reg_file[6411] <= 8'h03;
            reg_file[6412] <= 8'h93;
            reg_file[6413] <= 8'h97;
            reg_file[6414] <= 8'h07;
            reg_file[6415] <= 8'h01;
            reg_file[6416] <= 8'hB3;
            reg_file[6417] <= 8'hE7;
            reg_file[6418] <= 8'hF9;
            reg_file[6419] <= 8'h00;
            reg_file[6420] <= 8'h63;
            reg_file[6421] <= 8'hFE;
            reg_file[6422] <= 8'hE7;
            reg_file[6423] <= 8'h00;
            reg_file[6424] <= 8'hB3;
            reg_file[6425] <= 8'h87;
            reg_file[6426] <= 8'h07;
            reg_file[6427] <= 8'h01;
            reg_file[6428] <= 8'h13;
            reg_file[6429] <= 8'h83;
            reg_file[6430] <= 8'hFE;
            reg_file[6431] <= 8'hFF;
            reg_file[6432] <= 8'h63;
            reg_file[6433] <= 8'hE8;
            reg_file[6434] <= 8'h07;
            reg_file[6435] <= 8'h01;
            reg_file[6436] <= 8'h63;
            reg_file[6437] <= 8'hF6;
            reg_file[6438] <= 8'hE7;
            reg_file[6439] <= 8'h00;
            reg_file[6440] <= 8'h13;
            reg_file[6441] <= 8'h83;
            reg_file[6442] <= 8'hEE;
            reg_file[6443] <= 8'hFF;
            reg_file[6444] <= 8'hB3;
            reg_file[6445] <= 8'h87;
            reg_file[6446] <= 8'h07;
            reg_file[6447] <= 8'h01;
            reg_file[6448] <= 8'h33;
            reg_file[6449] <= 8'h87;
            reg_file[6450] <= 8'hE7;
            reg_file[6451] <= 8'h40;
            reg_file[6452] <= 8'h93;
            reg_file[6453] <= 8'h9F;
            reg_file[6454] <= 8'h0F;
            reg_file[6455] <= 8'h01;
            reg_file[6456] <= 8'hB7;
            reg_file[6457] <= 8'h07;
            reg_file[6458] <= 8'h01;
            reg_file[6459] <= 8'h00;
            reg_file[6460] <= 8'hB3;
            reg_file[6461] <= 8'hEF;
            reg_file[6462] <= 8'h6F;
            reg_file[6463] <= 8'h00;
            reg_file[6464] <= 8'h13;
            reg_file[6465] <= 8'h83;
            reg_file[6466] <= 8'hF7;
            reg_file[6467] <= 8'hFF;
            reg_file[6468] <= 8'h33;
            reg_file[6469] <= 8'hFF;
            reg_file[6470] <= 8'h6F;
            reg_file[6471] <= 8'h00;
            reg_file[6472] <= 8'h93;
            reg_file[6473] <= 8'hD2;
            reg_file[6474] <= 8'h0F;
            reg_file[6475] <= 8'h01;
            reg_file[6476] <= 8'h93;
            reg_file[6477] <= 8'hDE;
            reg_file[6478] <= 8'h08;
            reg_file[6479] <= 8'h01;
            reg_file[6480] <= 8'h33;
            reg_file[6481] <= 8'hF3;
            reg_file[6482] <= 8'h68;
            reg_file[6483] <= 8'h00;
            reg_file[6484] <= 8'h33;
            reg_file[6485] <= 8'h04;
            reg_file[6486] <= 8'h6F;
            reg_file[6487] <= 8'h02;
            reg_file[6488] <= 8'hB3;
            reg_file[6489] <= 8'h89;
            reg_file[6490] <= 8'h62;
            reg_file[6491] <= 8'h02;
            reg_file[6492] <= 8'h33;
            reg_file[6493] <= 8'h8F;
            reg_file[6494] <= 8'hEE;
            reg_file[6495] <= 8'h03;
            reg_file[6496] <= 8'hB3;
            reg_file[6497] <= 8'h03;
            reg_file[6498] <= 8'h3F;
            reg_file[6499] <= 8'h01;
            reg_file[6500] <= 8'h13;
            reg_file[6501] <= 8'h5F;
            reg_file[6502] <= 8'h04;
            reg_file[6503] <= 8'h01;
            reg_file[6504] <= 8'h33;
            reg_file[6505] <= 8'h0F;
            reg_file[6506] <= 8'h7F;
            reg_file[6507] <= 8'h00;
            reg_file[6508] <= 8'hB3;
            reg_file[6509] <= 8'h82;
            reg_file[6510] <= 8'hD2;
            reg_file[6511] <= 8'h03;
            reg_file[6512] <= 8'h63;
            reg_file[6513] <= 8'h74;
            reg_file[6514] <= 8'h3F;
            reg_file[6515] <= 8'h01;
            reg_file[6516] <= 8'hB3;
            reg_file[6517] <= 8'h82;
            reg_file[6518] <= 8'hF2;
            reg_file[6519] <= 8'h00;
            reg_file[6520] <= 8'hB7;
            reg_file[6521] <= 8'h03;
            reg_file[6522] <= 8'h01;
            reg_file[6523] <= 8'h00;
            reg_file[6524] <= 8'h93;
            reg_file[6525] <= 8'h57;
            reg_file[6526] <= 8'h0F;
            reg_file[6527] <= 8'h01;
            reg_file[6528] <= 8'h93;
            reg_file[6529] <= 8'h83;
            reg_file[6530] <= 8'hF3;
            reg_file[6531] <= 8'hFF;
            reg_file[6532] <= 8'hB3;
            reg_file[6533] <= 8'h82;
            reg_file[6534] <= 8'h57;
            reg_file[6535] <= 8'h00;
            reg_file[6536] <= 8'hB3;
            reg_file[6537] <= 8'h77;
            reg_file[6538] <= 8'h7F;
            reg_file[6539] <= 8'h00;
            reg_file[6540] <= 8'h93;
            reg_file[6541] <= 8'h97;
            reg_file[6542] <= 8'h07;
            reg_file[6543] <= 8'h01;
            reg_file[6544] <= 8'h33;
            reg_file[6545] <= 8'h74;
            reg_file[6546] <= 8'h74;
            reg_file[6547] <= 8'h00;
            reg_file[6548] <= 8'hB3;
            reg_file[6549] <= 8'h87;
            reg_file[6550] <= 8'h87;
            reg_file[6551] <= 8'h00;
            reg_file[6552] <= 8'h63;
            reg_file[6553] <= 8'h68;
            reg_file[6554] <= 8'h57;
            reg_file[6555] <= 8'h00;
            reg_file[6556] <= 8'h13;
            reg_file[6557] <= 8'h84;
            reg_file[6558] <= 8'h0F;
            reg_file[6559] <= 8'h00;
            reg_file[6560] <= 8'h63;
            reg_file[6561] <= 8'h14;
            reg_file[6562] <= 8'h57;
            reg_file[6563] <= 8'h04;
            reg_file[6564] <= 8'h63;
            reg_file[6565] <= 8'hF2;
            reg_file[6566] <= 8'hF6;
            reg_file[6567] <= 8'h04;
            reg_file[6568] <= 8'hB3;
            reg_file[6569] <= 8'h86;
            reg_file[6570] <= 8'h16;
            reg_file[6571] <= 8'h01;
            reg_file[6572] <= 8'h33;
            reg_file[6573] <= 8'hBF;
            reg_file[6574] <= 8'h16;
            reg_file[6575] <= 8'h01;
            reg_file[6576] <= 8'h33;
            reg_file[6577] <= 8'h0F;
            reg_file[6578] <= 8'h0F;
            reg_file[6579] <= 8'h01;
            reg_file[6580] <= 8'h33;
            reg_file[6581] <= 8'h07;
            reg_file[6582] <= 8'hE7;
            reg_file[6583] <= 8'h01;
            reg_file[6584] <= 8'h13;
            reg_file[6585] <= 8'h84;
            reg_file[6586] <= 8'hFF;
            reg_file[6587] <= 8'hFF;
            reg_file[6588] <= 8'h63;
            reg_file[6589] <= 8'h66;
            reg_file[6590] <= 8'hE8;
            reg_file[6591] <= 8'h00;
            reg_file[6592] <= 8'h63;
            reg_file[6593] <= 8'h14;
            reg_file[6594] <= 8'hE8;
            reg_file[6595] <= 8'h02;
            reg_file[6596] <= 8'h63;
            reg_file[6597] <= 8'hE2;
            reg_file[6598] <= 8'h16;
            reg_file[6599] <= 8'h03;
            reg_file[6600] <= 8'h63;
            reg_file[6601] <= 8'h66;
            reg_file[6602] <= 8'h57;
            reg_file[6603] <= 8'h00;
            reg_file[6604] <= 8'h63;
            reg_file[6605] <= 8'h9E;
            reg_file[6606] <= 8'hE2;
            reg_file[6607] <= 8'h00;
            reg_file[6608] <= 8'h63;
            reg_file[6609] <= 8'hFC;
            reg_file[6610] <= 8'hF6;
            reg_file[6611] <= 8'h00;
            reg_file[6612] <= 8'hB3;
            reg_file[6613] <= 8'h86;
            reg_file[6614] <= 8'h16;
            reg_file[6615] <= 8'h01;
            reg_file[6616] <= 8'h33;
            reg_file[6617] <= 8'hBF;
            reg_file[6618] <= 8'h16;
            reg_file[6619] <= 8'h01;
            reg_file[6620] <= 8'h33;
            reg_file[6621] <= 8'h0F;
            reg_file[6622] <= 8'h0F;
            reg_file[6623] <= 8'h01;
            reg_file[6624] <= 8'h13;
            reg_file[6625] <= 8'h84;
            reg_file[6626] <= 8'hEF;
            reg_file[6627] <= 8'hFF;
            reg_file[6628] <= 8'h33;
            reg_file[6629] <= 8'h07;
            reg_file[6630] <= 8'hE7;
            reg_file[6631] <= 8'h01;
            reg_file[6632] <= 8'h33;
            reg_file[6633] <= 8'h8F;
            reg_file[6634] <= 8'hF6;
            reg_file[6635] <= 8'h40;
            reg_file[6636] <= 8'h33;
            reg_file[6637] <= 8'h07;
            reg_file[6638] <= 8'h57;
            reg_file[6639] <= 8'h40;
            reg_file[6640] <= 8'hB3;
            reg_file[6641] <= 8'hB6;
            reg_file[6642] <= 8'hE6;
            reg_file[6643] <= 8'h01;
            reg_file[6644] <= 8'h33;
            reg_file[6645] <= 8'h07;
            reg_file[6646] <= 8'hD7;
            reg_file[6647] <= 8'h40;
            reg_file[6648] <= 8'h93;
            reg_file[6649] <= 8'h07;
            reg_file[6650] <= 8'hF0;
            reg_file[6651] <= 8'hFF;
            reg_file[6652] <= 8'h63;
            reg_file[6653] <= 8'h04;
            reg_file[6654] <= 8'hE8;
            reg_file[6655] <= 8'h12;
            reg_file[6656] <= 8'hB3;
            reg_file[6657] <= 8'h52;
            reg_file[6658] <= 8'hA7;
            reg_file[6659] <= 8'h02;
            reg_file[6660] <= 8'h93;
            reg_file[6661] <= 8'h57;
            reg_file[6662] <= 8'h0F;
            reg_file[6663] <= 8'h01;
            reg_file[6664] <= 8'h33;
            reg_file[6665] <= 8'h77;
            reg_file[6666] <= 8'hA7;
            reg_file[6667] <= 8'h02;
            reg_file[6668] <= 8'h93;
            reg_file[6669] <= 8'h86;
            reg_file[6670] <= 8'h02;
            reg_file[6671] <= 8'h00;
            reg_file[6672] <= 8'hB3;
            reg_file[6673] <= 8'h0F;
            reg_file[6674] <= 8'h5E;
            reg_file[6675] <= 8'h02;
            reg_file[6676] <= 8'h13;
            reg_file[6677] <= 8'h17;
            reg_file[6678] <= 8'h07;
            reg_file[6679] <= 8'h01;
            reg_file[6680] <= 8'h33;
            reg_file[6681] <= 8'hE7;
            reg_file[6682] <= 8'hE7;
            reg_file[6683] <= 8'h00;
            reg_file[6684] <= 8'h63;
            reg_file[6685] <= 8'h7E;
            reg_file[6686] <= 8'hF7;
            reg_file[6687] <= 8'h01;
            reg_file[6688] <= 8'h33;
            reg_file[6689] <= 8'h07;
            reg_file[6690] <= 8'h07;
            reg_file[6691] <= 8'h01;
            reg_file[6692] <= 8'h93;
            reg_file[6693] <= 8'h86;
            reg_file[6694] <= 8'hF2;
            reg_file[6695] <= 8'hFF;
            reg_file[6696] <= 8'h63;
            reg_file[6697] <= 8'h68;
            reg_file[6698] <= 8'h07;
            reg_file[6699] <= 8'h01;
            reg_file[6700] <= 8'h63;
            reg_file[6701] <= 8'h76;
            reg_file[6702] <= 8'hF7;
            reg_file[6703] <= 8'h01;
            reg_file[6704] <= 8'h93;
            reg_file[6705] <= 8'h86;
            reg_file[6706] <= 8'hE2;
            reg_file[6707] <= 8'hFF;
            reg_file[6708] <= 8'h33;
            reg_file[6709] <= 8'h07;
            reg_file[6710] <= 8'h07;
            reg_file[6711] <= 8'h01;
            reg_file[6712] <= 8'h33;
            reg_file[6713] <= 8'h07;
            reg_file[6714] <= 8'hF7;
            reg_file[6715] <= 8'h41;
            reg_file[6716] <= 8'hB3;
            reg_file[6717] <= 8'h5F;
            reg_file[6718] <= 8'hA7;
            reg_file[6719] <= 8'h02;
            reg_file[6720] <= 8'h93;
            reg_file[6721] <= 8'h17;
            reg_file[6722] <= 8'h0F;
            reg_file[6723] <= 8'h01;
            reg_file[6724] <= 8'h93;
            reg_file[6725] <= 8'hD7;
            reg_file[6726] <= 8'h07;
            reg_file[6727] <= 8'h01;
            reg_file[6728] <= 8'h33;
            reg_file[6729] <= 8'h77;
            reg_file[6730] <= 8'hA7;
            reg_file[6731] <= 8'h02;
            reg_file[6732] <= 8'h33;
            reg_file[6733] <= 8'h0E;
            reg_file[6734] <= 8'hFE;
            reg_file[6735] <= 8'h03;
            reg_file[6736] <= 8'h13;
            reg_file[6737] <= 8'h17;
            reg_file[6738] <= 8'h07;
            reg_file[6739] <= 8'h01;
            reg_file[6740] <= 8'h33;
            reg_file[6741] <= 8'hE7;
            reg_file[6742] <= 8'hE7;
            reg_file[6743] <= 8'h00;
            reg_file[6744] <= 8'h93;
            reg_file[6745] <= 8'h87;
            reg_file[6746] <= 8'h0F;
            reg_file[6747] <= 8'h00;
            reg_file[6748] <= 8'h63;
            reg_file[6749] <= 8'h7E;
            reg_file[6750] <= 8'hC7;
            reg_file[6751] <= 8'h01;
            reg_file[6752] <= 8'h33;
            reg_file[6753] <= 8'h07;
            reg_file[6754] <= 8'h07;
            reg_file[6755] <= 8'h01;
            reg_file[6756] <= 8'h93;
            reg_file[6757] <= 8'h87;
            reg_file[6758] <= 8'hFF;
            reg_file[6759] <= 8'hFF;
            reg_file[6760] <= 8'h63;
            reg_file[6761] <= 8'h68;
            reg_file[6762] <= 8'h07;
            reg_file[6763] <= 8'h01;
            reg_file[6764] <= 8'h63;
            reg_file[6765] <= 8'h76;
            reg_file[6766] <= 8'hC7;
            reg_file[6767] <= 8'h01;
            reg_file[6768] <= 8'h93;
            reg_file[6769] <= 8'h87;
            reg_file[6770] <= 8'hEF;
            reg_file[6771] <= 8'hFF;
            reg_file[6772] <= 8'h33;
            reg_file[6773] <= 8'h07;
            reg_file[6774] <= 8'h07;
            reg_file[6775] <= 8'h01;
            reg_file[6776] <= 8'h93;
            reg_file[6777] <= 8'h96;
            reg_file[6778] <= 8'h06;
            reg_file[6779] <= 8'h01;
            reg_file[6780] <= 8'hB3;
            reg_file[6781] <= 8'hE6;
            reg_file[6782] <= 8'hF6;
            reg_file[6783] <= 8'h00;
            reg_file[6784] <= 8'h93;
            reg_file[6785] <= 8'h97;
            reg_file[6786] <= 8'h06;
            reg_file[6787] <= 8'h01;
            reg_file[6788] <= 8'h93;
            reg_file[6789] <= 8'hD7;
            reg_file[6790] <= 8'h07;
            reg_file[6791] <= 8'h01;
            reg_file[6792] <= 8'h33;
            reg_file[6793] <= 8'h07;
            reg_file[6794] <= 8'hC7;
            reg_file[6795] <= 8'h41;
            reg_file[6796] <= 8'h13;
            reg_file[6797] <= 8'hDE;
            reg_file[6798] <= 8'h06;
            reg_file[6799] <= 8'h01;
            reg_file[6800] <= 8'h33;
            reg_file[6801] <= 8'h0F;
            reg_file[6802] <= 8'hF3;
            reg_file[6803] <= 8'h02;
            reg_file[6804] <= 8'h33;
            reg_file[6805] <= 8'h03;
            reg_file[6806] <= 8'h6E;
            reg_file[6807] <= 8'h02;
            reg_file[6808] <= 8'h33;
            reg_file[6809] <= 8'h8E;
            reg_file[6810] <= 8'hCE;
            reg_file[6811] <= 8'h03;
            reg_file[6812] <= 8'hB3;
            reg_file[6813] <= 8'h8E;
            reg_file[6814] <= 8'hFE;
            reg_file[6815] <= 8'h02;
            reg_file[6816] <= 8'h93;
            reg_file[6817] <= 8'h57;
            reg_file[6818] <= 8'h0F;
            reg_file[6819] <= 8'h01;
            reg_file[6820] <= 8'hB3;
            reg_file[6821] <= 8'h8E;
            reg_file[6822] <= 8'h6E;
            reg_file[6823] <= 8'h00;
            reg_file[6824] <= 8'hB3;
            reg_file[6825] <= 8'h87;
            reg_file[6826] <= 8'hD7;
            reg_file[6827] <= 8'h01;
            reg_file[6828] <= 8'h63;
            reg_file[6829] <= 8'hF6;
            reg_file[6830] <= 8'h67;
            reg_file[6831] <= 8'h00;
            reg_file[6832] <= 8'h37;
            reg_file[6833] <= 8'h05;
            reg_file[6834] <= 8'h01;
            reg_file[6835] <= 8'h00;
            reg_file[6836] <= 8'h33;
            reg_file[6837] <= 8'h0E;
            reg_file[6838] <= 8'hAE;
            reg_file[6839] <= 8'h00;
            reg_file[6840] <= 8'h13;
            reg_file[6841] <= 8'hD3;
            reg_file[6842] <= 8'h07;
            reg_file[6843] <= 8'h01;
            reg_file[6844] <= 8'h33;
            reg_file[6845] <= 8'h03;
            reg_file[6846] <= 8'hC3;
            reg_file[6847] <= 8'h01;
            reg_file[6848] <= 8'h37;
            reg_file[6849] <= 8'h0E;
            reg_file[6850] <= 8'h01;
            reg_file[6851] <= 8'h00;
            reg_file[6852] <= 8'h13;
            reg_file[6853] <= 8'h0E;
            reg_file[6854] <= 8'hFE;
            reg_file[6855] <= 8'hFF;
            reg_file[6856] <= 8'h33;
            reg_file[6857] <= 8'hF5;
            reg_file[6858] <= 8'hC7;
            reg_file[6859] <= 8'h01;
            reg_file[6860] <= 8'h13;
            reg_file[6861] <= 8'h15;
            reg_file[6862] <= 8'h05;
            reg_file[6863] <= 8'h01;
            reg_file[6864] <= 8'h33;
            reg_file[6865] <= 8'h7F;
            reg_file[6866] <= 8'hCF;
            reg_file[6867] <= 8'h01;
            reg_file[6868] <= 8'h33;
            reg_file[6869] <= 8'h05;
            reg_file[6870] <= 8'hE5;
            reg_file[6871] <= 8'h01;
            reg_file[6872] <= 8'h63;
            reg_file[6873] <= 8'h68;
            reg_file[6874] <= 8'h67;
            reg_file[6875] <= 8'h00;
            reg_file[6876] <= 8'h63;
            reg_file[6877] <= 8'h14;
            reg_file[6878] <= 8'h67;
            reg_file[6879] <= 8'h3E;
            reg_file[6880] <= 8'h93;
            reg_file[6881] <= 8'h87;
            reg_file[6882] <= 8'h06;
            reg_file[6883] <= 8'h00;
            reg_file[6884] <= 8'h63;
            reg_file[6885] <= 8'h00;
            reg_file[6886] <= 8'h05;
            reg_file[6887] <= 8'h04;
            reg_file[6888] <= 8'h33;
            reg_file[6889] <= 8'h07;
            reg_file[6890] <= 8'hE8;
            reg_file[6891] <= 8'h00;
            reg_file[6892] <= 8'h93;
            reg_file[6893] <= 8'h87;
            reg_file[6894] <= 8'hF6;
            reg_file[6895] <= 8'hFF;
            reg_file[6896] <= 8'h63;
            reg_file[6897] <= 8'h64;
            reg_file[6898] <= 8'h07;
            reg_file[6899] <= 8'h03;
            reg_file[6900] <= 8'h63;
            reg_file[6901] <= 8'h66;
            reg_file[6902] <= 8'h67;
            reg_file[6903] <= 8'h00;
            reg_file[6904] <= 8'h63;
            reg_file[6905] <= 8'h14;
            reg_file[6906] <= 8'h67;
            reg_file[6907] <= 8'h3C;
            reg_file[6908] <= 8'h63;
            reg_file[6909] <= 8'hF0;
            reg_file[6910] <= 8'hA8;
            reg_file[6911] <= 8'h02;
            reg_file[6912] <= 8'h93;
            reg_file[6913] <= 8'h87;
            reg_file[6914] <= 8'hE6;
            reg_file[6915] <= 8'hFF;
            reg_file[6916] <= 8'h93;
            reg_file[6917] <= 8'h96;
            reg_file[6918] <= 8'h18;
            reg_file[6919] <= 8'h00;
            reg_file[6920] <= 8'hB3;
            reg_file[6921] <= 8'hB8;
            reg_file[6922] <= 8'h16;
            reg_file[6923] <= 8'h01;
            reg_file[6924] <= 8'h33;
            reg_file[6925] <= 8'h88;
            reg_file[6926] <= 8'h08;
            reg_file[6927] <= 8'h01;
            reg_file[6928] <= 8'h33;
            reg_file[6929] <= 8'h07;
            reg_file[6930] <= 8'h07;
            reg_file[6931] <= 8'h01;
            reg_file[6932] <= 8'h93;
            reg_file[6933] <= 8'h88;
            reg_file[6934] <= 8'h06;
            reg_file[6935] <= 8'h00;
            reg_file[6936] <= 8'h63;
            reg_file[6937] <= 8'h14;
            reg_file[6938] <= 8'h67;
            reg_file[6939] <= 8'h00;
            reg_file[6940] <= 8'h63;
            reg_file[6941] <= 8'h84;
            reg_file[6942] <= 8'hA8;
            reg_file[6943] <= 8'h00;
            reg_file[6944] <= 8'h93;
            reg_file[6945] <= 8'hE7;
            reg_file[6946] <= 8'h17;
            reg_file[6947] <= 8'h00;
            reg_file[6948] <= 8'h13;
            reg_file[6949] <= 8'h88;
            reg_file[6950] <= 8'hF5;
            reg_file[6951] <= 8'h3F;
            reg_file[6952] <= 8'h63;
            reg_file[6953] <= 8'h5A;
            reg_file[6954] <= 8'h00;
            reg_file[6955] <= 8'h19;
            reg_file[6956] <= 8'h13;
            reg_file[6957] <= 8'hF7;
            reg_file[6958] <= 8'h77;
            reg_file[6959] <= 8'h00;
            reg_file[6960] <= 8'h63;
            reg_file[6961] <= 8'h0A;
            reg_file[6962] <= 8'h07;
            reg_file[6963] <= 8'h0A;
            reg_file[6964] <= 8'h13;
            reg_file[6965] <= 8'h07;
            reg_file[6966] <= 8'h20;
            reg_file[6967] <= 8'h00;
            reg_file[6968] <= 8'h93;
            reg_file[6969] <= 8'hE4;
            reg_file[6970] <= 8'h14;
            reg_file[6971] <= 8'h00;
            reg_file[6972] <= 8'h63;
            reg_file[6973] <= 8'h02;
            reg_file[6974] <= 8'hE9;
            reg_file[6975] <= 8'h0A;
            reg_file[6976] <= 8'h13;
            reg_file[6977] <= 8'h07;
            reg_file[6978] <= 8'h30;
            reg_file[6979] <= 8'h00;
            reg_file[6980] <= 8'h63;
            reg_file[6981] <= 8'h08;
            reg_file[6982] <= 8'hE9;
            reg_file[6983] <= 8'h08;
            reg_file[6984] <= 8'h63;
            reg_file[6985] <= 8'h1E;
            reg_file[6986] <= 8'h09;
            reg_file[6987] <= 8'h08;
            reg_file[6988] <= 8'h13;
            reg_file[6989] <= 8'hF7;
            reg_file[6990] <= 8'hF7;
            reg_file[6991] <= 8'h00;
            reg_file[6992] <= 8'h93;
            reg_file[6993] <= 8'h06;
            reg_file[6994] <= 8'h40;
            reg_file[6995] <= 8'h00;
            reg_file[6996] <= 8'h63;
            reg_file[6997] <= 8'h08;
            reg_file[6998] <= 8'hD7;
            reg_file[6999] <= 8'h08;
            reg_file[7000] <= 8'h13;
            reg_file[7001] <= 8'h87;
            reg_file[7002] <= 8'h47;
            reg_file[7003] <= 8'h00;
            reg_file[7004] <= 8'hB3;
            reg_file[7005] <= 8'h37;
            reg_file[7006] <= 8'hF7;
            reg_file[7007] <= 8'h00;
            reg_file[7008] <= 8'h33;
            reg_file[7009] <= 8'h04;
            reg_file[7010] <= 8'hF4;
            reg_file[7011] <= 8'h00;
            reg_file[7012] <= 8'h93;
            reg_file[7013] <= 8'h07;
            reg_file[7014] <= 8'h07;
            reg_file[7015] <= 8'h00;
            reg_file[7016] <= 8'h6F;
            reg_file[7017] <= 8'h00;
            reg_file[7018] <= 8'hC0;
            reg_file[7019] <= 8'h07;
            reg_file[7020] <= 8'h93;
            reg_file[7021] <= 8'h85;
            reg_file[7022] <= 8'hF5;
            reg_file[7023] <= 8'hFF;
            reg_file[7024] <= 8'h93;
            reg_file[7025] <= 8'h06;
            reg_file[7026] <= 8'h00;
            reg_file[7027] <= 8'h00;
            reg_file[7028] <= 8'h6F;
            reg_file[7029] <= 8'hF0;
            reg_file[7030] <= 8'h9F;
            reg_file[7031] <= 8'hD2;
            reg_file[7032] <= 8'h13;
            reg_file[7033] <= 8'h06;
            reg_file[7034] <= 8'h0A;
            reg_file[7035] <= 8'h00;
            reg_file[7036] <= 8'h13;
            reg_file[7037] <= 8'h84;
            reg_file[7038] <= 8'h0B;
            reg_file[7039] <= 8'h00;
            reg_file[7040] <= 8'h93;
            reg_file[7041] <= 8'h87;
            reg_file[7042] <= 8'h09;
            reg_file[7043] <= 8'h00;
            reg_file[7044] <= 8'h13;
            reg_file[7045] <= 8'h87;
            reg_file[7046] <= 8'h0C;
            reg_file[7047] <= 8'h00;
            reg_file[7048] <= 8'h93;
            reg_file[7049] <= 8'h06;
            reg_file[7050] <= 8'h30;
            reg_file[7051] <= 8'h00;
            reg_file[7052] <= 8'h63;
            reg_file[7053] <= 8'h00;
            reg_file[7054] <= 8'hD7;
            reg_file[7055] <= 8'h32;
            reg_file[7056] <= 8'h93;
            reg_file[7057] <= 8'h06;
            reg_file[7058] <= 8'h10;
            reg_file[7059] <= 8'h00;
            reg_file[7060] <= 8'h63;
            reg_file[7061] <= 8'h06;
            reg_file[7062] <= 8'hD7;
            reg_file[7063] <= 8'h30;
            reg_file[7064] <= 8'h93;
            reg_file[7065] <= 8'h06;
            reg_file[7066] <= 8'h20;
            reg_file[7067] <= 8'h00;
            reg_file[7068] <= 8'hE3;
            reg_file[7069] <= 8'h14;
            reg_file[7070] <= 8'hD7;
            reg_file[7071] <= 8'hF8;
            reg_file[7072] <= 8'h6F;
            reg_file[7073] <= 8'h00;
            reg_file[7074] <= 8'h00;
            reg_file[7075] <= 8'h01;
            reg_file[7076] <= 8'h13;
            reg_file[7077] <= 8'h86;
            reg_file[7078] <= 8'h0A;
            reg_file[7079] <= 8'h00;
            reg_file[7080] <= 8'h6F;
            reg_file[7081] <= 8'hF0;
            reg_file[7082] <= 8'h1F;
            reg_file[7083] <= 8'hFE;
            reg_file[7084] <= 8'h93;
            reg_file[7085] <= 8'hE4;
            reg_file[7086] <= 8'h84;
            reg_file[7087] <= 8'h00;
            reg_file[7088] <= 8'h13;
            reg_file[7089] <= 8'h05;
            reg_file[7090] <= 8'h00;
            reg_file[7091] <= 8'h00;
            reg_file[7092] <= 8'h93;
            reg_file[7093] <= 8'h07;
            reg_file[7094] <= 8'h00;
            reg_file[7095] <= 8'h00;
            reg_file[7096] <= 8'h13;
            reg_file[7097] <= 8'h07;
            reg_file[7098] <= 8'hF0;
            reg_file[7099] <= 8'h7F;
            reg_file[7100] <= 8'h6F;
            reg_file[7101] <= 8'h00;
            reg_file[7102] <= 8'hC0;
            reg_file[7103] <= 8'h05;
            reg_file[7104] <= 8'h37;
            reg_file[7105] <= 8'h04;
            reg_file[7106] <= 8'h08;
            reg_file[7107] <= 8'h00;
            reg_file[7108] <= 8'h93;
            reg_file[7109] <= 8'h07;
            reg_file[7110] <= 8'h00;
            reg_file[7111] <= 8'h00;
            reg_file[7112] <= 8'h13;
            reg_file[7113] <= 8'h06;
            reg_file[7114] <= 8'h00;
            reg_file[7115] <= 8'h00;
            reg_file[7116] <= 8'h13;
            reg_file[7117] <= 8'h07;
            reg_file[7118] <= 8'h30;
            reg_file[7119] <= 8'h00;
            reg_file[7120] <= 8'h6F;
            reg_file[7121] <= 8'hF0;
            reg_file[7122] <= 8'h9F;
            reg_file[7123] <= 8'hFB;
            reg_file[7124] <= 8'h63;
            reg_file[7125] <= 8'h18;
            reg_file[7126] <= 8'h06;
            reg_file[7127] <= 8'h00;
            reg_file[7128] <= 8'h13;
            reg_file[7129] <= 8'h87;
            reg_file[7130] <= 8'h87;
            reg_file[7131] <= 8'h00;
            reg_file[7132] <= 8'h6F;
            reg_file[7133] <= 8'hF0;
            reg_file[7134] <= 8'h1F;
            reg_file[7135] <= 8'hF8;
            reg_file[7136] <= 8'hE3;
            reg_file[7137] <= 8'h1C;
            reg_file[7138] <= 8'h06;
            reg_file[7139] <= 8'hFE;
            reg_file[7140] <= 8'h13;
            reg_file[7141] <= 8'h17;
            reg_file[7142] <= 8'h74;
            reg_file[7143] <= 8'h00;
            reg_file[7144] <= 8'h63;
            reg_file[7145] <= 8'h5A;
            reg_file[7146] <= 8'h07;
            reg_file[7147] <= 8'h00;
            reg_file[7148] <= 8'h37;
            reg_file[7149] <= 8'h07;
            reg_file[7150] <= 8'h00;
            reg_file[7151] <= 8'hFF;
            reg_file[7152] <= 8'h13;
            reg_file[7153] <= 8'h07;
            reg_file[7154] <= 8'hF7;
            reg_file[7155] <= 8'hFF;
            reg_file[7156] <= 8'h33;
            reg_file[7157] <= 8'h74;
            reg_file[7158] <= 8'hE4;
            reg_file[7159] <= 8'h00;
            reg_file[7160] <= 8'h13;
            reg_file[7161] <= 8'h88;
            reg_file[7162] <= 8'h05;
            reg_file[7163] <= 8'h40;
            reg_file[7164] <= 8'h13;
            reg_file[7165] <= 8'h07;
            reg_file[7166] <= 8'hE0;
            reg_file[7167] <= 8'h7F;
            reg_file[7168] <= 8'h63;
            reg_file[7169] <= 8'h4E;
            reg_file[7170] <= 8'h07;
            reg_file[7171] <= 8'h07;
            reg_file[7172] <= 8'h13;
            reg_file[7173] <= 8'hD7;
            reg_file[7174] <= 8'h37;
            reg_file[7175] <= 8'h00;
            reg_file[7176] <= 8'h93;
            reg_file[7177] <= 8'h17;
            reg_file[7178] <= 8'hD4;
            reg_file[7179] <= 8'h01;
            reg_file[7180] <= 8'hB3;
            reg_file[7181] <= 8'hE7;
            reg_file[7182] <= 8'hE7;
            reg_file[7183] <= 8'h00;
            reg_file[7184] <= 8'h13;
            reg_file[7185] <= 8'h55;
            reg_file[7186] <= 8'h34;
            reg_file[7187] <= 8'h00;
            reg_file[7188] <= 8'h13;
            reg_file[7189] <= 8'h07;
            reg_file[7190] <= 8'h08;
            reg_file[7191] <= 8'h00;
            reg_file[7192] <= 8'h13;
            reg_file[7193] <= 8'h17;
            reg_file[7194] <= 8'h47;
            reg_file[7195] <= 8'h01;
            reg_file[7196] <= 8'hB7;
            reg_file[7197] <= 8'h06;
            reg_file[7198] <= 8'hF0;
            reg_file[7199] <= 8'h7F;
            reg_file[7200] <= 8'h13;
            reg_file[7201] <= 8'h15;
            reg_file[7202] <= 8'hC5;
            reg_file[7203] <= 8'h00;
            reg_file[7204] <= 8'h33;
            reg_file[7205] <= 8'h77;
            reg_file[7206] <= 8'hD7;
            reg_file[7207] <= 8'h00;
            reg_file[7208] <= 8'h13;
            reg_file[7209] <= 8'h55;
            reg_file[7210] <= 8'hC5;
            reg_file[7211] <= 8'h00;
            reg_file[7212] <= 8'h33;
            reg_file[7213] <= 8'h65;
            reg_file[7214] <= 8'hA7;
            reg_file[7215] <= 8'h00;
            reg_file[7216] <= 8'h13;
            reg_file[7217] <= 8'h16;
            reg_file[7218] <= 8'hF6;
            reg_file[7219] <= 8'h01;
            reg_file[7220] <= 8'h33;
            reg_file[7221] <= 8'h67;
            reg_file[7222] <= 8'hC5;
            reg_file[7223] <= 8'h00;
            reg_file[7224] <= 8'h93;
            reg_file[7225] <= 8'h05;
            reg_file[7226] <= 8'h07;
            reg_file[7227] <= 8'h00;
            reg_file[7228] <= 8'h13;
            reg_file[7229] <= 8'h85;
            reg_file[7230] <= 8'h07;
            reg_file[7231] <= 8'h00;
            reg_file[7232] <= 8'h63;
            reg_file[7233] <= 8'h84;
            reg_file[7234] <= 8'h04;
            reg_file[7235] <= 8'h00;
            reg_file[7236] <= 8'h73;
            reg_file[7237] <= 8'hA0;
            reg_file[7238] <= 8'h14;
            reg_file[7239] <= 8'h00;
            reg_file[7240] <= 8'h83;
            reg_file[7241] <= 8'h20;
            reg_file[7242] <= 8'hC1;
            reg_file[7243] <= 8'h02;
            reg_file[7244] <= 8'h03;
            reg_file[7245] <= 8'h24;
            reg_file[7246] <= 8'h81;
            reg_file[7247] <= 8'h02;
            reg_file[7248] <= 8'h83;
            reg_file[7249] <= 8'h24;
            reg_file[7250] <= 8'h41;
            reg_file[7251] <= 8'h02;
            reg_file[7252] <= 8'h03;
            reg_file[7253] <= 8'h29;
            reg_file[7254] <= 8'h01;
            reg_file[7255] <= 8'h02;
            reg_file[7256] <= 8'h83;
            reg_file[7257] <= 8'h29;
            reg_file[7258] <= 8'hC1;
            reg_file[7259] <= 8'h01;
            reg_file[7260] <= 8'h03;
            reg_file[7261] <= 8'h2A;
            reg_file[7262] <= 8'h81;
            reg_file[7263] <= 8'h01;
            reg_file[7264] <= 8'h83;
            reg_file[7265] <= 8'h2A;
            reg_file[7266] <= 8'h41;
            reg_file[7267] <= 8'h01;
            reg_file[7268] <= 8'h03;
            reg_file[7269] <= 8'h2B;
            reg_file[7270] <= 8'h01;
            reg_file[7271] <= 8'h01;
            reg_file[7272] <= 8'h83;
            reg_file[7273] <= 8'h2B;
            reg_file[7274] <= 8'hC1;
            reg_file[7275] <= 8'h00;
            reg_file[7276] <= 8'h03;
            reg_file[7277] <= 8'h2C;
            reg_file[7278] <= 8'h81;
            reg_file[7279] <= 8'h00;
            reg_file[7280] <= 8'h83;
            reg_file[7281] <= 8'h2C;
            reg_file[7282] <= 8'h41;
            reg_file[7283] <= 8'h00;
            reg_file[7284] <= 8'h13;
            reg_file[7285] <= 8'h01;
            reg_file[7286] <= 8'h01;
            reg_file[7287] <= 8'h03;
            reg_file[7288] <= 8'h67;
            reg_file[7289] <= 8'h80;
            reg_file[7290] <= 8'h00;
            reg_file[7291] <= 8'h00;
            reg_file[7292] <= 8'h93;
            reg_file[7293] <= 8'h07;
            reg_file[7294] <= 8'h20;
            reg_file[7295] <= 8'h00;
            reg_file[7296] <= 8'h63;
            reg_file[7297] <= 8'h0A;
            reg_file[7298] <= 8'hF9;
            reg_file[7299] <= 8'h02;
            reg_file[7300] <= 8'h93;
            reg_file[7301] <= 8'h07;
            reg_file[7302] <= 8'h30;
            reg_file[7303] <= 8'h00;
            reg_file[7304] <= 8'h63;
            reg_file[7305] <= 8'h0A;
            reg_file[7306] <= 8'hF9;
            reg_file[7307] <= 8'h00;
            reg_file[7308] <= 8'h63;
            reg_file[7309] <= 8'h1A;
            reg_file[7310] <= 8'h09;
            reg_file[7311] <= 8'h00;
            reg_file[7312] <= 8'h93;
            reg_file[7313] <= 8'h07;
            reg_file[7314] <= 8'h00;
            reg_file[7315] <= 8'h00;
            reg_file[7316] <= 8'h13;
            reg_file[7317] <= 8'h07;
            reg_file[7318] <= 8'hF0;
            reg_file[7319] <= 8'h7F;
            reg_file[7320] <= 8'h6F;
            reg_file[7321] <= 8'h00;
            reg_file[7322] <= 8'h00;
            reg_file[7323] <= 8'h01;
            reg_file[7324] <= 8'hE3;
            reg_file[7325] <= 8'h0A;
            reg_file[7326] <= 8'h06;
            reg_file[7327] <= 8'hFE;
            reg_file[7328] <= 8'h93;
            reg_file[7329] <= 8'h07;
            reg_file[7330] <= 8'hF0;
            reg_file[7331] <= 8'hFF;
            reg_file[7332] <= 8'h13;
            reg_file[7333] <= 8'h07;
            reg_file[7334] <= 8'hE0;
            reg_file[7335] <= 8'h7F;
            reg_file[7336] <= 8'h93;
            reg_file[7337] <= 8'hE4;
            reg_file[7338] <= 8'h54;
            reg_file[7339] <= 8'h00;
            reg_file[7340] <= 8'h13;
            reg_file[7341] <= 8'h85;
            reg_file[7342] <= 8'h07;
            reg_file[7343] <= 8'h00;
            reg_file[7344] <= 8'h6F;
            reg_file[7345] <= 8'hF0;
            reg_file[7346] <= 8'h9F;
            reg_file[7347] <= 8'hF6;
            reg_file[7348] <= 8'hE3;
            reg_file[7349] <= 8'h1E;
            reg_file[7350] <= 8'h06;
            reg_file[7351] <= 8'hFC;
            reg_file[7352] <= 8'h6F;
            reg_file[7353] <= 8'hF0;
            reg_file[7354] <= 8'h9F;
            reg_file[7355] <= 8'hFE;
            reg_file[7356] <= 8'h13;
            reg_file[7357] <= 8'h07;
            reg_file[7358] <= 8'h10;
            reg_file[7359] <= 8'h00;
            reg_file[7360] <= 8'h63;
            reg_file[7361] <= 8'h16;
            reg_file[7362] <= 8'h08;
            reg_file[7363] <= 8'h06;
            reg_file[7364] <= 8'h93;
            reg_file[7365] <= 8'hF6;
            reg_file[7366] <= 8'h77;
            reg_file[7367] <= 8'h00;
            reg_file[7368] <= 8'h13;
            reg_file[7369] <= 8'h07;
            reg_file[7370] <= 8'h04;
            reg_file[7371] <= 8'h00;
            reg_file[7372] <= 8'h63;
            reg_file[7373] <= 8'h8A;
            reg_file[7374] <= 8'h06;
            reg_file[7375] <= 8'h04;
            reg_file[7376] <= 8'h13;
            reg_file[7377] <= 8'h07;
            reg_file[7378] <= 8'h20;
            reg_file[7379] <= 8'h00;
            reg_file[7380] <= 8'h93;
            reg_file[7381] <= 8'hE4;
            reg_file[7382] <= 8'h14;
            reg_file[7383] <= 8'h00;
            reg_file[7384] <= 8'h63;
            reg_file[7385] <= 8'h00;
            reg_file[7386] <= 8'hE9;
            reg_file[7387] <= 8'h04;
            reg_file[7388] <= 8'h13;
            reg_file[7389] <= 8'h07;
            reg_file[7390] <= 8'h30;
            reg_file[7391] <= 8'h00;
            reg_file[7392] <= 8'h63;
            reg_file[7393] <= 8'h04;
            reg_file[7394] <= 8'hE9;
            reg_file[7395] <= 8'h02;
            reg_file[7396] <= 8'h13;
            reg_file[7397] <= 8'h07;
            reg_file[7398] <= 8'h04;
            reg_file[7399] <= 8'h00;
            reg_file[7400] <= 8'h63;
            reg_file[7401] <= 8'h1C;
            reg_file[7402] <= 8'h09;
            reg_file[7403] <= 8'h02;
            reg_file[7404] <= 8'h93;
            reg_file[7405] <= 8'hF6;
            reg_file[7406] <= 8'hF7;
            reg_file[7407] <= 8'h00;
            reg_file[7408] <= 8'h13;
            reg_file[7409] <= 8'h05;
            reg_file[7410] <= 8'h40;
            reg_file[7411] <= 8'h00;
            reg_file[7412] <= 8'h63;
            reg_file[7413] <= 8'h86;
            reg_file[7414] <= 8'hA6;
            reg_file[7415] <= 8'h02;
            reg_file[7416] <= 8'h13;
            reg_file[7417] <= 8'hB7;
            reg_file[7418] <= 8'hC7;
            reg_file[7419] <= 8'hFF;
            reg_file[7420] <= 8'h13;
            reg_file[7421] <= 8'h47;
            reg_file[7422] <= 8'h17;
            reg_file[7423] <= 8'h00;
            reg_file[7424] <= 8'h33;
            reg_file[7425] <= 8'h07;
            reg_file[7426] <= 8'h87;
            reg_file[7427] <= 8'h00;
            reg_file[7428] <= 8'h6F;
            reg_file[7429] <= 8'h00;
            reg_file[7430] <= 8'hC0;
            reg_file[7431] <= 8'h01;
            reg_file[7432] <= 8'h13;
            reg_file[7433] <= 8'h07;
            reg_file[7434] <= 8'h04;
            reg_file[7435] <= 8'h00;
            reg_file[7436] <= 8'h63;
            reg_file[7437] <= 8'h1A;
            reg_file[7438] <= 8'h06;
            reg_file[7439] <= 8'h00;
            reg_file[7440] <= 8'h13;
            reg_file[7441] <= 8'hB7;
            reg_file[7442] <= 8'h87;
            reg_file[7443] <= 8'hFF;
            reg_file[7444] <= 8'h6F;
            reg_file[7445] <= 8'hF0;
            reg_file[7446] <= 8'h9F;
            reg_file[7447] <= 8'hFE;
            reg_file[7448] <= 8'h13;
            reg_file[7449] <= 8'h07;
            reg_file[7450] <= 8'h04;
            reg_file[7451] <= 8'h00;
            reg_file[7452] <= 8'hE3;
            reg_file[7453] <= 8'h1A;
            reg_file[7454] <= 8'h06;
            reg_file[7455] <= 8'hFE;
            reg_file[7456] <= 8'h13;
            reg_file[7457] <= 8'h57;
            reg_file[7458] <= 8'h87;
            reg_file[7459] <= 8'h01;
            reg_file[7460] <= 8'h13;
            reg_file[7461] <= 8'h47;
            reg_file[7462] <= 8'h17;
            reg_file[7463] <= 8'h00;
            reg_file[7464] <= 8'h13;
            reg_file[7465] <= 8'h77;
            reg_file[7466] <= 8'h17;
            reg_file[7467] <= 8'h00;
            reg_file[7468] <= 8'h13;
            reg_file[7469] <= 8'h05;
            reg_file[7470] <= 8'h10;
            reg_file[7471] <= 8'h00;
            reg_file[7472] <= 8'h33;
            reg_file[7473] <= 8'h05;
            reg_file[7474] <= 8'h05;
            reg_file[7475] <= 8'h41;
            reg_file[7476] <= 8'h93;
            reg_file[7477] <= 8'h06;
            reg_file[7478] <= 8'h80;
            reg_file[7479] <= 8'h03;
            reg_file[7480] <= 8'h63;
            reg_file[7481] <= 8'hCC;
            reg_file[7482] <= 8'hA6;
            reg_file[7483] <= 8'h0E;
            reg_file[7484] <= 8'h93;
            reg_file[7485] <= 8'h06;
            reg_file[7486] <= 8'hF0;
            reg_file[7487] <= 8'h01;
            reg_file[7488] <= 8'h63;
            reg_file[7489] <= 8'hC2;
            reg_file[7490] <= 8'hA6;
            reg_file[7491] <= 8'h06;
            reg_file[7492] <= 8'h93;
            reg_file[7493] <= 8'h85;
            reg_file[7494] <= 8'hE5;
            reg_file[7495] <= 8'h41;
            reg_file[7496] <= 8'h33;
            reg_file[7497] <= 8'hD8;
            reg_file[7498] <= 8'hA7;
            reg_file[7499] <= 8'h00;
            reg_file[7500] <= 8'hB3;
            reg_file[7501] <= 8'h16;
            reg_file[7502] <= 8'hB4;
            reg_file[7503] <= 8'h00;
            reg_file[7504] <= 8'hB3;
            reg_file[7505] <= 8'h97;
            reg_file[7506] <= 8'hB7;
            reg_file[7507] <= 8'h00;
            reg_file[7508] <= 8'hB3;
            reg_file[7509] <= 8'hE6;
            reg_file[7510] <= 8'h06;
            reg_file[7511] <= 8'h01;
            reg_file[7512] <= 8'hB3;
            reg_file[7513] <= 8'h37;
            reg_file[7514] <= 8'hF0;
            reg_file[7515] <= 8'h00;
            reg_file[7516] <= 8'hB3;
            reg_file[7517] <= 8'hE7;
            reg_file[7518] <= 8'hF6;
            reg_file[7519] <= 8'h00;
            reg_file[7520] <= 8'h33;
            reg_file[7521] <= 8'h55;
            reg_file[7522] <= 8'hA4;
            reg_file[7523] <= 8'h00;
            reg_file[7524] <= 8'h93;
            reg_file[7525] <= 8'hF6;
            reg_file[7526] <= 8'h77;
            reg_file[7527] <= 8'h00;
            reg_file[7528] <= 8'h63;
            reg_file[7529] <= 8'h80;
            reg_file[7530] <= 8'h06;
            reg_file[7531] <= 8'h08;
            reg_file[7532] <= 8'h93;
            reg_file[7533] <= 8'h06;
            reg_file[7534] <= 8'h20;
            reg_file[7535] <= 8'h00;
            reg_file[7536] <= 8'h93;
            reg_file[7537] <= 8'hE4;
            reg_file[7538] <= 8'h14;
            reg_file[7539] <= 8'h00;
            reg_file[7540] <= 8'h63;
            reg_file[7541] <= 8'h08;
            reg_file[7542] <= 8'hD9;
            reg_file[7543] <= 8'h06;
            reg_file[7544] <= 8'h93;
            reg_file[7545] <= 8'h06;
            reg_file[7546] <= 8'h30;
            reg_file[7547] <= 8'h00;
            reg_file[7548] <= 8'h63;
            reg_file[7549] <= 8'h0E;
            reg_file[7550] <= 8'hD9;
            reg_file[7551] <= 8'h04;
            reg_file[7552] <= 8'h63;
            reg_file[7553] <= 8'h14;
            reg_file[7554] <= 8'h09;
            reg_file[7555] <= 8'h06;
            reg_file[7556] <= 8'h93;
            reg_file[7557] <= 8'hF6;
            reg_file[7558] <= 8'hF7;
            reg_file[7559] <= 8'h00;
            reg_file[7560] <= 8'h93;
            reg_file[7561] <= 8'h05;
            reg_file[7562] <= 8'h40;
            reg_file[7563] <= 8'h00;
            reg_file[7564] <= 8'h63;
            reg_file[7565] <= 8'h8E;
            reg_file[7566] <= 8'hB6;
            reg_file[7567] <= 8'h04;
            reg_file[7568] <= 8'h93;
            reg_file[7569] <= 8'h86;
            reg_file[7570] <= 8'h47;
            reg_file[7571] <= 8'h00;
            reg_file[7572] <= 8'hB3;
            reg_file[7573] <= 8'hB7;
            reg_file[7574] <= 8'hF6;
            reg_file[7575] <= 8'h00;
            reg_file[7576] <= 8'h33;
            reg_file[7577] <= 8'h05;
            reg_file[7578] <= 8'hF5;
            reg_file[7579] <= 8'h00;
            reg_file[7580] <= 8'h93;
            reg_file[7581] <= 8'h87;
            reg_file[7582] <= 8'h06;
            reg_file[7583] <= 8'h00;
            reg_file[7584] <= 8'h6F;
            reg_file[7585] <= 8'h00;
            reg_file[7586] <= 8'h80;
            reg_file[7587] <= 8'h04;
            reg_file[7588] <= 8'h93;
            reg_file[7589] <= 8'h06;
            reg_file[7590] <= 8'h10;
            reg_file[7591] <= 8'hFE;
            reg_file[7592] <= 8'hB3;
            reg_file[7593] <= 8'h86;
            reg_file[7594] <= 8'h06;
            reg_file[7595] <= 8'h41;
            reg_file[7596] <= 8'h93;
            reg_file[7597] <= 8'h08;
            reg_file[7598] <= 8'h00;
            reg_file[7599] <= 8'h02;
            reg_file[7600] <= 8'hB3;
            reg_file[7601] <= 8'h56;
            reg_file[7602] <= 8'hD4;
            reg_file[7603] <= 8'h00;
            reg_file[7604] <= 8'h13;
            reg_file[7605] <= 8'h08;
            reg_file[7606] <= 8'h00;
            reg_file[7607] <= 8'h00;
            reg_file[7608] <= 8'h63;
            reg_file[7609] <= 8'h06;
            reg_file[7610] <= 8'h15;
            reg_file[7611] <= 8'h01;
            reg_file[7612] <= 8'h93;
            reg_file[7613] <= 8'h85;
            reg_file[7614] <= 8'hE5;
            reg_file[7615] <= 8'h43;
            reg_file[7616] <= 8'h33;
            reg_file[7617] <= 8'h18;
            reg_file[7618] <= 8'hB4;
            reg_file[7619] <= 8'h00;
            reg_file[7620] <= 8'hB3;
            reg_file[7621] <= 8'h67;
            reg_file[7622] <= 8'hF8;
            reg_file[7623] <= 8'h00;
            reg_file[7624] <= 8'hB3;
            reg_file[7625] <= 8'h37;
            reg_file[7626] <= 8'hF0;
            reg_file[7627] <= 8'h00;
            reg_file[7628] <= 8'hB3;
            reg_file[7629] <= 8'hE7;
            reg_file[7630] <= 8'hF6;
            reg_file[7631] <= 8'h00;
            reg_file[7632] <= 8'h13;
            reg_file[7633] <= 8'h05;
            reg_file[7634] <= 8'h00;
            reg_file[7635] <= 8'h00;
            reg_file[7636] <= 8'h6F;
            reg_file[7637] <= 8'hF0;
            reg_file[7638] <= 8'h1F;
            reg_file[7639] <= 8'hF9;
            reg_file[7640] <= 8'h63;
            reg_file[7641] <= 8'h18;
            reg_file[7642] <= 8'h06;
            reg_file[7643] <= 8'h00;
            reg_file[7644] <= 8'h93;
            reg_file[7645] <= 8'h86;
            reg_file[7646] <= 8'h87;
            reg_file[7647] <= 8'h00;
            reg_file[7648] <= 8'h6F;
            reg_file[7649] <= 8'hF0;
            reg_file[7650] <= 8'h5F;
            reg_file[7651] <= 8'hFB;
            reg_file[7652] <= 8'hE3;
            reg_file[7653] <= 8'h1C;
            reg_file[7654] <= 8'h06;
            reg_file[7655] <= 8'hFE;
            reg_file[7656] <= 8'h93;
            reg_file[7657] <= 8'h16;
            reg_file[7658] <= 8'h85;
            reg_file[7659] <= 8'h00;
            reg_file[7660] <= 8'h63;
            reg_file[7661] <= 8'hDE;
            reg_file[7662] <= 8'h06;
            reg_file[7663] <= 8'h00;
            reg_file[7664] <= 8'h93;
            reg_file[7665] <= 8'hE4;
            reg_file[7666] <= 8'h14;
            reg_file[7667] <= 8'h00;
            reg_file[7668] <= 8'h13;
            reg_file[7669] <= 8'h05;
            reg_file[7670] <= 8'h00;
            reg_file[7671] <= 8'h00;
            reg_file[7672] <= 8'h93;
            reg_file[7673] <= 8'h07;
            reg_file[7674] <= 8'h00;
            reg_file[7675] <= 8'h00;
            reg_file[7676] <= 8'h63;
            reg_file[7677] <= 8'h16;
            reg_file[7678] <= 8'h07;
            reg_file[7679] <= 8'h02;
            reg_file[7680] <= 8'h13;
            reg_file[7681] <= 8'h07;
            reg_file[7682] <= 8'h10;
            reg_file[7683] <= 8'h00;
            reg_file[7684] <= 8'h6F;
            reg_file[7685] <= 8'hF0;
            reg_file[7686] <= 8'h5F;
            reg_file[7687] <= 8'hE1;
            reg_file[7688] <= 8'h93;
            reg_file[7689] <= 8'hD6;
            reg_file[7690] <= 8'h37;
            reg_file[7691] <= 8'h00;
            reg_file[7692] <= 8'h93;
            reg_file[7693] <= 8'h17;
            reg_file[7694] <= 8'hD5;
            reg_file[7695] <= 8'h01;
            reg_file[7696] <= 8'hB3;
            reg_file[7697] <= 8'hE7;
            reg_file[7698] <= 8'hD7;
            reg_file[7699] <= 8'h00;
            reg_file[7700] <= 8'h13;
            reg_file[7701] <= 8'h55;
            reg_file[7702] <= 8'h35;
            reg_file[7703] <= 8'h00;
            reg_file[7704] <= 8'hE3;
            reg_file[7705] <= 8'h00;
            reg_file[7706] <= 8'h07;
            reg_file[7707] <= 8'hE0;
            reg_file[7708] <= 8'h13;
            reg_file[7709] <= 8'hF7;
            reg_file[7710] <= 8'h14;
            reg_file[7711] <= 8'h00;
            reg_file[7712] <= 8'hE3;
            reg_file[7713] <= 8'h0C;
            reg_file[7714] <= 8'h07;
            reg_file[7715] <= 8'hDE;
            reg_file[7716] <= 8'h13;
            reg_file[7717] <= 8'h07;
            reg_file[7718] <= 8'h00;
            reg_file[7719] <= 8'h00;
            reg_file[7720] <= 8'h93;
            reg_file[7721] <= 8'hE4;
            reg_file[7722] <= 8'h24;
            reg_file[7723] <= 8'h00;
            reg_file[7724] <= 8'h6F;
            reg_file[7725] <= 8'hF0;
            reg_file[7726] <= 8'hDF;
            reg_file[7727] <= 8'hDE;
            reg_file[7728] <= 8'hB3;
            reg_file[7729] <= 8'hE7;
            reg_file[7730] <= 8'h87;
            reg_file[7731] <= 8'h00;
            reg_file[7732] <= 8'h63;
            reg_file[7733] <= 8'h84;
            reg_file[7734] <= 8'h07;
            reg_file[7735] <= 8'h02;
            reg_file[7736] <= 8'h93;
            reg_file[7737] <= 8'h07;
            reg_file[7738] <= 8'h20;
            reg_file[7739] <= 8'h00;
            reg_file[7740] <= 8'h93;
            reg_file[7741] <= 8'hE4;
            reg_file[7742] <= 8'h14;
            reg_file[7743] <= 8'h00;
            reg_file[7744] <= 8'h63;
            reg_file[7745] <= 8'h0E;
            reg_file[7746] <= 8'hF9;
            reg_file[7747] <= 8'h02;
            reg_file[7748] <= 8'h93;
            reg_file[7749] <= 8'h07;
            reg_file[7750] <= 8'h30;
            reg_file[7751] <= 8'h00;
            reg_file[7752] <= 8'h63;
            reg_file[7753] <= 8'h02;
            reg_file[7754] <= 8'hF9;
            reg_file[7755] <= 8'h02;
            reg_file[7756] <= 8'h93;
            reg_file[7757] <= 8'h07;
            reg_file[7758] <= 8'h10;
            reg_file[7759] <= 8'h00;
            reg_file[7760] <= 8'h63;
            reg_file[7761] <= 8'h14;
            reg_file[7762] <= 8'h09;
            reg_file[7763] <= 8'h00;
            reg_file[7764] <= 8'h93;
            reg_file[7765] <= 8'h07;
            reg_file[7766] <= 8'h50;
            reg_file[7767] <= 8'h00;
            reg_file[7768] <= 8'h93;
            reg_file[7769] <= 8'hD7;
            reg_file[7770] <= 8'h37;
            reg_file[7771] <= 8'h00;
            reg_file[7772] <= 8'h93;
            reg_file[7773] <= 8'hE4;
            reg_file[7774] <= 8'h24;
            reg_file[7775] <= 8'h00;
            reg_file[7776] <= 8'h13;
            reg_file[7777] <= 8'h05;
            reg_file[7778] <= 8'h00;
            reg_file[7779] <= 8'h00;
            reg_file[7780] <= 8'h13;
            reg_file[7781] <= 8'h07;
            reg_file[7782] <= 8'h00;
            reg_file[7783] <= 8'h00;
            reg_file[7784] <= 8'h6F;
            reg_file[7785] <= 8'hF0;
            reg_file[7786] <= 8'h1F;
            reg_file[7787] <= 8'hDB;
            reg_file[7788] <= 8'h93;
            reg_file[7789] <= 8'h07;
            reg_file[7790] <= 8'h90;
            reg_file[7791] <= 8'h00;
            reg_file[7792] <= 8'hE3;
            reg_file[7793] <= 8'h04;
            reg_file[7794] <= 8'h06;
            reg_file[7795] <= 8'hFE;
            reg_file[7796] <= 8'h93;
            reg_file[7797] <= 8'h07;
            reg_file[7798] <= 8'h10;
            reg_file[7799] <= 8'h00;
            reg_file[7800] <= 8'h6F;
            reg_file[7801] <= 8'hF0;
            reg_file[7802] <= 8'h1F;
            reg_file[7803] <= 8'hFE;
            reg_file[7804] <= 8'h93;
            reg_file[7805] <= 8'h07;
            reg_file[7806] <= 8'h90;
            reg_file[7807] <= 8'h00;
            reg_file[7808] <= 8'hE3;
            reg_file[7809] <= 8'h1C;
            reg_file[7810] <= 8'h06;
            reg_file[7811] <= 8'hFC;
            reg_file[7812] <= 8'h6F;
            reg_file[7813] <= 8'hF0;
            reg_file[7814] <= 8'h1F;
            reg_file[7815] <= 8'hFF;
            reg_file[7816] <= 8'h37;
            reg_file[7817] <= 8'h05;
            reg_file[7818] <= 8'h08;
            reg_file[7819] <= 8'h00;
            reg_file[7820] <= 8'h93;
            reg_file[7821] <= 8'h07;
            reg_file[7822] <= 8'h00;
            reg_file[7823] <= 8'h00;
            reg_file[7824] <= 8'h13;
            reg_file[7825] <= 8'h07;
            reg_file[7826] <= 8'hF0;
            reg_file[7827] <= 8'h7F;
            reg_file[7828] <= 8'h13;
            reg_file[7829] <= 8'h06;
            reg_file[7830] <= 8'h00;
            reg_file[7831] <= 8'h00;
            reg_file[7832] <= 8'h93;
            reg_file[7833] <= 8'h04;
            reg_file[7834] <= 8'h00;
            reg_file[7835] <= 8'h01;
            reg_file[7836] <= 8'h6F;
            reg_file[7837] <= 8'hF0;
            reg_file[7838] <= 8'hDF;
            reg_file[7839] <= 8'hD7;
            reg_file[7840] <= 8'h13;
            reg_file[7841] <= 8'h05;
            reg_file[7842] <= 8'h00;
            reg_file[7843] <= 8'h00;
            reg_file[7844] <= 8'h93;
            reg_file[7845] <= 8'h07;
            reg_file[7846] <= 8'h00;
            reg_file[7847] <= 8'h00;
            reg_file[7848] <= 8'h6F;
            reg_file[7849] <= 8'hF0;
            reg_file[7850] <= 8'hDF;
            reg_file[7851] <= 8'hFB;
            reg_file[7852] <= 8'h37;
            reg_file[7853] <= 8'h05;
            reg_file[7854] <= 8'h08;
            reg_file[7855] <= 8'h00;
            reg_file[7856] <= 8'h93;
            reg_file[7857] <= 8'h07;
            reg_file[7858] <= 8'h00;
            reg_file[7859] <= 8'h00;
            reg_file[7860] <= 8'h13;
            reg_file[7861] <= 8'h07;
            reg_file[7862] <= 8'hF0;
            reg_file[7863] <= 8'h7F;
            reg_file[7864] <= 8'h13;
            reg_file[7865] <= 8'h06;
            reg_file[7866] <= 8'h00;
            reg_file[7867] <= 8'h00;
            reg_file[7868] <= 8'h6F;
            reg_file[7869] <= 8'hF0;
            reg_file[7870] <= 8'hDF;
            reg_file[7871] <= 8'hD5;
            reg_file[7872] <= 8'h93;
            reg_file[7873] <= 8'h86;
            reg_file[7874] <= 8'h07;
            reg_file[7875] <= 8'h00;
            reg_file[7876] <= 8'h93;
            reg_file[7877] <= 8'h87;
            reg_file[7878] <= 8'h06;
            reg_file[7879] <= 8'h00;
            reg_file[7880] <= 8'h6F;
            reg_file[7881] <= 8'hF0;
            reg_file[7882] <= 8'h9F;
            reg_file[7883] <= 8'hC5;
            reg_file[7884] <= 8'h13;
            reg_file[7885] <= 8'h01;
            reg_file[7886] <= 8'h01;
            reg_file[7887] <= 8'hFD;
            reg_file[7888] <= 8'h23;
            reg_file[7889] <= 8'h24;
            reg_file[7890] <= 8'h81;
            reg_file[7891] <= 8'h02;
            reg_file[7892] <= 8'h23;
            reg_file[7893] <= 8'h28;
            reg_file[7894] <= 8'h61;
            reg_file[7895] <= 8'h01;
            reg_file[7896] <= 8'h23;
            reg_file[7897] <= 8'h22;
            reg_file[7898] <= 8'h91;
            reg_file[7899] <= 8'h01;
            reg_file[7900] <= 8'h23;
            reg_file[7901] <= 8'h26;
            reg_file[7902] <= 8'h11;
            reg_file[7903] <= 8'h02;
            reg_file[7904] <= 8'h23;
            reg_file[7905] <= 8'h22;
            reg_file[7906] <= 8'h91;
            reg_file[7907] <= 8'h02;
            reg_file[7908] <= 8'h23;
            reg_file[7909] <= 8'h20;
            reg_file[7910] <= 8'h21;
            reg_file[7911] <= 8'h03;
            reg_file[7912] <= 8'h23;
            reg_file[7913] <= 8'h2E;
            reg_file[7914] <= 8'h31;
            reg_file[7915] <= 8'h01;
            reg_file[7916] <= 8'h23;
            reg_file[7917] <= 8'h2C;
            reg_file[7918] <= 8'h41;
            reg_file[7919] <= 8'h01;
            reg_file[7920] <= 8'h23;
            reg_file[7921] <= 8'h2A;
            reg_file[7922] <= 8'h51;
            reg_file[7923] <= 8'h01;
            reg_file[7924] <= 8'h23;
            reg_file[7925] <= 8'h26;
            reg_file[7926] <= 8'h71;
            reg_file[7927] <= 8'h01;
            reg_file[7928] <= 8'h23;
            reg_file[7929] <= 8'h24;
            reg_file[7930] <= 8'h81;
            reg_file[7931] <= 8'h01;
            reg_file[7932] <= 8'h13;
            reg_file[7933] <= 8'h04;
            reg_file[7934] <= 8'h05;
            reg_file[7935] <= 8'h00;
            reg_file[7936] <= 8'h93;
            reg_file[7937] <= 8'h0C;
            reg_file[7938] <= 8'h06;
            reg_file[7939] <= 8'h00;
            reg_file[7940] <= 8'h13;
            reg_file[7941] <= 8'h8B;
            reg_file[7942] <= 8'h06;
            reg_file[7943] <= 8'h00;
            reg_file[7944] <= 8'h73;
            reg_file[7945] <= 8'h29;
            reg_file[7946] <= 8'h20;
            reg_file[7947] <= 8'h00;
            reg_file[7948] <= 8'h93;
            reg_file[7949] <= 8'hD7;
            reg_file[7950] <= 8'h45;
            reg_file[7951] <= 8'h01;
            reg_file[7952] <= 8'h93;
            reg_file[7953] <= 8'h99;
            reg_file[7954] <= 8'hC5;
            reg_file[7955] <= 8'h00;
            reg_file[7956] <= 8'h13;
            reg_file[7957] <= 8'h97;
            reg_file[7958] <= 8'h57;
            reg_file[7959] <= 8'h01;
            reg_file[7960] <= 8'h93;
            reg_file[7961] <= 8'hD9;
            reg_file[7962] <= 8'hC9;
            reg_file[7963] <= 8'h00;
            reg_file[7964] <= 8'h93;
            reg_file[7965] <= 8'hDA;
            reg_file[7966] <= 8'hF5;
            reg_file[7967] <= 8'h01;
            reg_file[7968] <= 8'h63;
            reg_file[7969] <= 8'h0C;
            reg_file[7970] <= 8'h07;
            reg_file[7971] <= 8'h02;
            reg_file[7972] <= 8'h93;
            reg_file[7973] <= 8'hFB;
            reg_file[7974] <= 8'hF7;
            reg_file[7975] <= 8'h7F;
            reg_file[7976] <= 8'h93;
            reg_file[7977] <= 8'h07;
            reg_file[7978] <= 8'hF0;
            reg_file[7979] <= 8'h7F;
            reg_file[7980] <= 8'h63;
            reg_file[7981] <= 8'h88;
            reg_file[7982] <= 8'hFB;
            reg_file[7983] <= 8'h08;
            reg_file[7984] <= 8'h93;
            reg_file[7985] <= 8'h57;
            reg_file[7986] <= 8'hD5;
            reg_file[7987] <= 8'h01;
            reg_file[7988] <= 8'h93;
            reg_file[7989] <= 8'h99;
            reg_file[7990] <= 8'h39;
            reg_file[7991] <= 8'h00;
            reg_file[7992] <= 8'hB3;
            reg_file[7993] <= 8'hE9;
            reg_file[7994] <= 8'h37;
            reg_file[7995] <= 8'h01;
            reg_file[7996] <= 8'hB7;
            reg_file[7997] <= 8'h07;
            reg_file[7998] <= 8'h80;
            reg_file[7999] <= 8'h00;
            reg_file[8000] <= 8'hB3;
            reg_file[8001] <= 8'hE9;
            reg_file[8002] <= 8'hF9;
            reg_file[8003] <= 8'h00;
            reg_file[8004] <= 8'h13;
            reg_file[8005] <= 8'h1A;
            reg_file[8006] <= 8'h35;
            reg_file[8007] <= 8'h00;
            reg_file[8008] <= 8'h93;
            reg_file[8009] <= 8'h8B;
            reg_file[8010] <= 8'h1B;
            reg_file[8011] <= 8'hC0;
            reg_file[8012] <= 8'h13;
            reg_file[8013] <= 8'h0C;
            reg_file[8014] <= 8'h00;
            reg_file[8015] <= 8'h00;
            reg_file[8016] <= 8'h93;
            reg_file[8017] <= 8'h04;
            reg_file[8018] <= 8'h00;
            reg_file[8019] <= 8'h00;
            reg_file[8020] <= 8'h6F;
            reg_file[8021] <= 8'h00;
            reg_file[8022] <= 8'h80;
            reg_file[8023] <= 8'h08;
            reg_file[8024] <= 8'hB3;
            reg_file[8025] <= 8'hE7;
            reg_file[8026] <= 8'hA9;
            reg_file[8027] <= 8'h00;
            reg_file[8028] <= 8'h63;
            reg_file[8029] <= 8'h80;
            reg_file[8030] <= 8'h07;
            reg_file[8031] <= 8'h10;
            reg_file[8032] <= 8'h63;
            reg_file[8033] <= 8'h80;
            reg_file[8034] <= 8'h09;
            reg_file[8035] <= 8'h04;
            reg_file[8036] <= 8'h13;
            reg_file[8037] <= 8'h85;
            reg_file[8038] <= 8'h09;
            reg_file[8039] <= 8'h00;
            reg_file[8040] <= 8'hEF;
            reg_file[8041] <= 8'h10;
            reg_file[8042] <= 8'h80;
            reg_file[8043] <= 8'h28;
            reg_file[8044] <= 8'h13;
            reg_file[8045] <= 8'h07;
            reg_file[8046] <= 8'h55;
            reg_file[8047] <= 8'hFF;
            reg_file[8048] <= 8'h93;
            reg_file[8049] <= 8'h07;
            reg_file[8050] <= 8'hC0;
            reg_file[8051] <= 8'h01;
            reg_file[8052] <= 8'h63;
            reg_file[8053] <= 8'hCC;
            reg_file[8054] <= 8'hE7;
            reg_file[8055] <= 8'h02;
            reg_file[8056] <= 8'h93;
            reg_file[8057] <= 8'h07;
            reg_file[8058] <= 8'hD0;
            reg_file[8059] <= 8'h01;
            reg_file[8060] <= 8'h13;
            reg_file[8061] <= 8'h0A;
            reg_file[8062] <= 8'h85;
            reg_file[8063] <= 8'hFF;
            reg_file[8064] <= 8'hB3;
            reg_file[8065] <= 8'h87;
            reg_file[8066] <= 8'hE7;
            reg_file[8067] <= 8'h40;
            reg_file[8068] <= 8'hB3;
            reg_file[8069] <= 8'h99;
            reg_file[8070] <= 8'h49;
            reg_file[8071] <= 8'h01;
            reg_file[8072] <= 8'hB3;
            reg_file[8073] <= 8'h57;
            reg_file[8074] <= 8'hF4;
            reg_file[8075] <= 8'h00;
            reg_file[8076] <= 8'hB3;
            reg_file[8077] <= 8'hE9;
            reg_file[8078] <= 8'h37;
            reg_file[8079] <= 8'h01;
            reg_file[8080] <= 8'h33;
            reg_file[8081] <= 8'h1A;
            reg_file[8082] <= 8'h44;
            reg_file[8083] <= 8'h01;
            reg_file[8084] <= 8'h93;
            reg_file[8085] <= 8'h0B;
            reg_file[8086] <= 8'hD0;
            reg_file[8087] <= 8'hC0;
            reg_file[8088] <= 8'hB3;
            reg_file[8089] <= 8'h8B;
            reg_file[8090] <= 8'hAB;
            reg_file[8091] <= 8'h40;
            reg_file[8092] <= 8'h6F;
            reg_file[8093] <= 8'hF0;
            reg_file[8094] <= 8'h1F;
            reg_file[8095] <= 8'hFB;
            reg_file[8096] <= 8'hEF;
            reg_file[8097] <= 8'h10;
            reg_file[8098] <= 8'h00;
            reg_file[8099] <= 8'h25;
            reg_file[8100] <= 8'h13;
            reg_file[8101] <= 8'h05;
            reg_file[8102] <= 8'h05;
            reg_file[8103] <= 8'h02;
            reg_file[8104] <= 8'h6F;
            reg_file[8105] <= 8'hF0;
            reg_file[8106] <= 8'h5F;
            reg_file[8107] <= 8'hFC;
            reg_file[8108] <= 8'h93;
            reg_file[8109] <= 8'h09;
            reg_file[8110] <= 8'h85;
            reg_file[8111] <= 8'hFD;
            reg_file[8112] <= 8'hB3;
            reg_file[8113] <= 8'h19;
            reg_file[8114] <= 8'h34;
            reg_file[8115] <= 8'h01;
            reg_file[8116] <= 8'h13;
            reg_file[8117] <= 8'h0A;
            reg_file[8118] <= 8'h00;
            reg_file[8119] <= 8'h00;
            reg_file[8120] <= 8'h6F;
            reg_file[8121] <= 8'hF0;
            reg_file[8122] <= 8'hDF;
            reg_file[8123] <= 8'hFD;
            reg_file[8124] <= 8'h33;
            reg_file[8125] <= 8'hE4;
            reg_file[8126] <= 8'hA9;
            reg_file[8127] <= 8'h00;
            reg_file[8128] <= 8'h63;
            reg_file[8129] <= 8'h08;
            reg_file[8130] <= 8'h04;
            reg_file[8131] <= 8'h0A;
            reg_file[8132] <= 8'h93;
            reg_file[8133] <= 8'h97;
            reg_file[8134] <= 8'hC9;
            reg_file[8135] <= 8'h00;
            reg_file[8136] <= 8'h13;
            reg_file[8137] <= 8'h0A;
            reg_file[8138] <= 8'h05;
            reg_file[8139] <= 8'h00;
            reg_file[8140] <= 8'h93;
            reg_file[8141] <= 8'h0B;
            reg_file[8142] <= 8'hF0;
            reg_file[8143] <= 8'h7F;
            reg_file[8144] <= 8'h13;
            reg_file[8145] <= 8'h0C;
            reg_file[8146] <= 8'h30;
            reg_file[8147] <= 8'h00;
            reg_file[8148] <= 8'h93;
            reg_file[8149] <= 8'h04;
            reg_file[8150] <= 8'h00;
            reg_file[8151] <= 8'h01;
            reg_file[8152] <= 8'hE3;
            reg_file[8153] <= 8'hCC;
            reg_file[8154] <= 8'h07;
            reg_file[8155] <= 8'hF6;
            reg_file[8156] <= 8'h13;
            reg_file[8157] <= 8'h57;
            reg_file[8158] <= 8'h4B;
            reg_file[8159] <= 8'h01;
            reg_file[8160] <= 8'h13;
            reg_file[8161] <= 8'h14;
            reg_file[8162] <= 8'hCB;
            reg_file[8163] <= 8'h00;
            reg_file[8164] <= 8'h93;
            reg_file[8165] <= 8'h16;
            reg_file[8166] <= 8'h57;
            reg_file[8167] <= 8'h01;
            reg_file[8168] <= 8'h93;
            reg_file[8169] <= 8'h87;
            reg_file[8170] <= 8'h0C;
            reg_file[8171] <= 8'h00;
            reg_file[8172] <= 8'h13;
            reg_file[8173] <= 8'h54;
            reg_file[8174] <= 8'hC4;
            reg_file[8175] <= 8'h00;
            reg_file[8176] <= 8'h13;
            reg_file[8177] <= 8'h75;
            reg_file[8178] <= 8'hF7;
            reg_file[8179] <= 8'h7F;
            reg_file[8180] <= 8'h13;
            reg_file[8181] <= 8'h5B;
            reg_file[8182] <= 8'hFB;
            reg_file[8183] <= 8'h01;
            reg_file[8184] <= 8'h63;
            reg_file[8185] <= 8'h86;
            reg_file[8186] <= 8'h06;
            reg_file[8187] <= 8'h08;
            reg_file[8188] <= 8'h13;
            reg_file[8189] <= 8'h07;
            reg_file[8190] <= 8'hF0;
            reg_file[8191] <= 8'h7F;
            reg_file[8192] <= 8'h63;
            reg_file[8193] <= 8'h06;
            reg_file[8194] <= 8'hE5;
            reg_file[8195] <= 8'h0E;
            reg_file[8196] <= 8'h93;
            reg_file[8197] <= 8'hD7;
            reg_file[8198] <= 8'hDC;
            reg_file[8199] <= 8'h01;
            reg_file[8200] <= 8'h13;
            reg_file[8201] <= 8'h14;
            reg_file[8202] <= 8'h34;
            reg_file[8203] <= 8'h00;
            reg_file[8204] <= 8'h33;
            reg_file[8205] <= 8'hE4;
            reg_file[8206] <= 8'h87;
            reg_file[8207] <= 8'h00;
            reg_file[8208] <= 8'hB7;
            reg_file[8209] <= 8'h07;
            reg_file[8210] <= 8'h80;
            reg_file[8211] <= 8'h00;
            reg_file[8212] <= 8'h33;
            reg_file[8213] <= 8'h64;
            reg_file[8214] <= 8'hF4;
            reg_file[8215] <= 8'h00;
            reg_file[8216] <= 8'h13;
            reg_file[8217] <= 8'h05;
            reg_file[8218] <= 8'h15;
            reg_file[8219] <= 8'hC0;
            reg_file[8220] <= 8'h93;
            reg_file[8221] <= 8'h97;
            reg_file[8222] <= 8'h3C;
            reg_file[8223] <= 8'h00;
            reg_file[8224] <= 8'h13;
            reg_file[8225] <= 8'h07;
            reg_file[8226] <= 8'h00;
            reg_file[8227] <= 8'h00;
            reg_file[8228] <= 8'h93;
            reg_file[8229] <= 8'h16;
            reg_file[8230] <= 8'h2C;
            reg_file[8231] <= 8'h00;
            reg_file[8232] <= 8'hB3;
            reg_file[8233] <= 8'hE6;
            reg_file[8234] <= 8'hE6;
            reg_file[8235] <= 8'h00;
            reg_file[8236] <= 8'hB3;
            reg_file[8237] <= 8'h8B;
            reg_file[8238] <= 8'hAB;
            reg_file[8239] <= 8'h00;
            reg_file[8240] <= 8'h93;
            reg_file[8241] <= 8'h86;
            reg_file[8242] <= 8'hF6;
            reg_file[8243] <= 8'hFF;
            reg_file[8244] <= 8'h13;
            reg_file[8245] <= 8'h06;
            reg_file[8246] <= 8'hE0;
            reg_file[8247] <= 8'h00;
            reg_file[8248] <= 8'hB3;
            reg_file[8249] <= 8'hC5;
            reg_file[8250] <= 8'h6A;
            reg_file[8251] <= 8'h01;
            reg_file[8252] <= 8'h13;
            reg_file[8253] <= 8'h85;
            reg_file[8254] <= 8'h1B;
            reg_file[8255] <= 8'h00;
            reg_file[8256] <= 8'h63;
            reg_file[8257] <= 8'h6A;
            reg_file[8258] <= 8'hD6;
            reg_file[8259] <= 8'h16;
            reg_file[8260] <= 8'h37;
            reg_file[8261] <= 8'h36;
            reg_file[8262] <= 8'h00;
            reg_file[8263] <= 8'h80;
            reg_file[8264] <= 8'h93;
            reg_file[8265] <= 8'h96;
            reg_file[8266] <= 8'h26;
            reg_file[8267] <= 8'h00;
            reg_file[8268] <= 8'h13;
            reg_file[8269] <= 8'h06;
            reg_file[8270] <= 8'h86;
            reg_file[8271] <= 8'h67;
            reg_file[8272] <= 8'hB3;
            reg_file[8273] <= 8'h86;
            reg_file[8274] <= 8'hC6;
            reg_file[8275] <= 8'h00;
            reg_file[8276] <= 8'h83;
            reg_file[8277] <= 8'hA6;
            reg_file[8278] <= 8'h06;
            reg_file[8279] <= 8'h00;
            reg_file[8280] <= 8'h67;
            reg_file[8281] <= 8'h80;
            reg_file[8282] <= 8'h06;
            reg_file[8283] <= 8'h00;
            reg_file[8284] <= 8'h93;
            reg_file[8285] <= 8'h09;
            reg_file[8286] <= 8'h00;
            reg_file[8287] <= 8'h00;
            reg_file[8288] <= 8'h13;
            reg_file[8289] <= 8'h0A;
            reg_file[8290] <= 8'h00;
            reg_file[8291] <= 8'h00;
            reg_file[8292] <= 8'h93;
            reg_file[8293] <= 8'h0B;
            reg_file[8294] <= 8'h00;
            reg_file[8295] <= 8'h00;
            reg_file[8296] <= 8'h13;
            reg_file[8297] <= 8'h0C;
            reg_file[8298] <= 8'h10;
            reg_file[8299] <= 8'h00;
            reg_file[8300] <= 8'h6F;
            reg_file[8301] <= 8'hF0;
            reg_file[8302] <= 8'h5F;
            reg_file[8303] <= 8'hEE;
            reg_file[8304] <= 8'h93;
            reg_file[8305] <= 8'h09;
            reg_file[8306] <= 8'h00;
            reg_file[8307] <= 8'h00;
            reg_file[8308] <= 8'h13;
            reg_file[8309] <= 8'h0A;
            reg_file[8310] <= 8'h00;
            reg_file[8311] <= 8'h00;
            reg_file[8312] <= 8'h93;
            reg_file[8313] <= 8'h0B;
            reg_file[8314] <= 8'hF0;
            reg_file[8315] <= 8'h7F;
            reg_file[8316] <= 8'h13;
            reg_file[8317] <= 8'h0C;
            reg_file[8318] <= 8'h20;
            reg_file[8319] <= 8'h00;
            reg_file[8320] <= 8'h6F;
            reg_file[8321] <= 8'hF0;
            reg_file[8322] <= 8'h1F;
            reg_file[8323] <= 8'hED;
            reg_file[8324] <= 8'hB3;
            reg_file[8325] <= 8'h67;
            reg_file[8326] <= 8'h94;
            reg_file[8327] <= 8'h01;
            reg_file[8328] <= 8'h63;
            reg_file[8329] <= 8'h82;
            reg_file[8330] <= 8'h07;
            reg_file[8331] <= 8'h08;
            reg_file[8332] <= 8'h63;
            reg_file[8333] <= 8'h00;
            reg_file[8334] <= 8'h04;
            reg_file[8335] <= 8'h04;
            reg_file[8336] <= 8'h13;
            reg_file[8337] <= 8'h05;
            reg_file[8338] <= 8'h04;
            reg_file[8339] <= 8'h00;
            reg_file[8340] <= 8'hEF;
            reg_file[8341] <= 8'h10;
            reg_file[8342] <= 8'hC0;
            reg_file[8343] <= 8'h15;
            reg_file[8344] <= 8'h93;
            reg_file[8345] <= 8'h06;
            reg_file[8346] <= 8'h55;
            reg_file[8347] <= 8'hFF;
            reg_file[8348] <= 8'h93;
            reg_file[8349] <= 8'h07;
            reg_file[8350] <= 8'hC0;
            reg_file[8351] <= 8'h01;
            reg_file[8352] <= 8'h63;
            reg_file[8353] <= 8'hCE;
            reg_file[8354] <= 8'hD7;
            reg_file[8355] <= 8'h02;
            reg_file[8356] <= 8'h13;
            reg_file[8357] <= 8'h07;
            reg_file[8358] <= 8'hD0;
            reg_file[8359] <= 8'h01;
            reg_file[8360] <= 8'h93;
            reg_file[8361] <= 8'h07;
            reg_file[8362] <= 8'h85;
            reg_file[8363] <= 8'hFF;
            reg_file[8364] <= 8'h33;
            reg_file[8365] <= 8'h07;
            reg_file[8366] <= 8'hD7;
            reg_file[8367] <= 8'h40;
            reg_file[8368] <= 8'h33;
            reg_file[8369] <= 8'h14;
            reg_file[8370] <= 8'hF4;
            reg_file[8371] <= 8'h00;
            reg_file[8372] <= 8'h33;
            reg_file[8373] <= 8'hD7;
            reg_file[8374] <= 8'hEC;
            reg_file[8375] <= 8'h00;
            reg_file[8376] <= 8'h33;
            reg_file[8377] <= 8'h64;
            reg_file[8378] <= 8'h87;
            reg_file[8379] <= 8'h00;
            reg_file[8380] <= 8'hB3;
            reg_file[8381] <= 8'h97;
            reg_file[8382] <= 8'hFC;
            reg_file[8383] <= 8'h00;
            reg_file[8384] <= 8'h13;
            reg_file[8385] <= 8'h07;
            reg_file[8386] <= 8'hD0;
            reg_file[8387] <= 8'hC0;
            reg_file[8388] <= 8'h33;
            reg_file[8389] <= 8'h05;
            reg_file[8390] <= 8'hA7;
            reg_file[8391] <= 8'h40;
            reg_file[8392] <= 8'h6F;
            reg_file[8393] <= 8'hF0;
            reg_file[8394] <= 8'h9F;
            reg_file[8395] <= 8'hF5;
            reg_file[8396] <= 8'h13;
            reg_file[8397] <= 8'h85;
            reg_file[8398] <= 8'h0C;
            reg_file[8399] <= 8'h00;
            reg_file[8400] <= 8'hEF;
            reg_file[8401] <= 8'h10;
            reg_file[8402] <= 8'h00;
            reg_file[8403] <= 8'h12;
            reg_file[8404] <= 8'h13;
            reg_file[8405] <= 8'h05;
            reg_file[8406] <= 8'h05;
            reg_file[8407] <= 8'h02;
            reg_file[8408] <= 8'h6F;
            reg_file[8409] <= 8'hF0;
            reg_file[8410] <= 8'h1F;
            reg_file[8411] <= 8'hFC;
            reg_file[8412] <= 8'h13;
            reg_file[8413] <= 8'h04;
            reg_file[8414] <= 8'h85;
            reg_file[8415] <= 8'hFD;
            reg_file[8416] <= 8'h33;
            reg_file[8417] <= 8'h94;
            reg_file[8418] <= 8'h8C;
            reg_file[8419] <= 8'h00;
            reg_file[8420] <= 8'h93;
            reg_file[8421] <= 8'h07;
            reg_file[8422] <= 8'h00;
            reg_file[8423] <= 8'h00;
            reg_file[8424] <= 8'h6F;
            reg_file[8425] <= 8'hF0;
            reg_file[8426] <= 8'h9F;
            reg_file[8427] <= 8'hFD;
            reg_file[8428] <= 8'h33;
            reg_file[8429] <= 8'h66;
            reg_file[8430] <= 8'h94;
            reg_file[8431] <= 8'h01;
            reg_file[8432] <= 8'h63;
            reg_file[8433] <= 8'h08;
            reg_file[8434] <= 8'h06;
            reg_file[8435] <= 8'h02;
            reg_file[8436] <= 8'h13;
            reg_file[8437] <= 8'h17;
            reg_file[8438] <= 8'hC4;
            reg_file[8439] <= 8'h00;
            reg_file[8440] <= 8'h13;
            reg_file[8441] <= 8'h05;
            reg_file[8442] <= 8'hF0;
            reg_file[8443] <= 8'h7F;
            reg_file[8444] <= 8'h63;
            reg_file[8445] <= 8'h4C;
            reg_file[8446] <= 8'h07;
            reg_file[8447] <= 8'h02;
            reg_file[8448] <= 8'h13;
            reg_file[8449] <= 8'h07;
            reg_file[8450] <= 8'h30;
            reg_file[8451] <= 8'h00;
            reg_file[8452] <= 8'h93;
            reg_file[8453] <= 8'h04;
            reg_file[8454] <= 8'h00;
            reg_file[8455] <= 8'h01;
            reg_file[8456] <= 8'h6F;
            reg_file[8457] <= 8'hF0;
            reg_file[8458] <= 8'hDF;
            reg_file[8459] <= 8'hF1;
            reg_file[8460] <= 8'h13;
            reg_file[8461] <= 8'h04;
            reg_file[8462] <= 8'h00;
            reg_file[8463] <= 8'h00;
            reg_file[8464] <= 8'h93;
            reg_file[8465] <= 8'h07;
            reg_file[8466] <= 8'h00;
            reg_file[8467] <= 8'h00;
            reg_file[8468] <= 8'h13;
            reg_file[8469] <= 8'h05;
            reg_file[8470] <= 8'h00;
            reg_file[8471] <= 8'h00;
            reg_file[8472] <= 8'h13;
            reg_file[8473] <= 8'h07;
            reg_file[8474] <= 8'h10;
            reg_file[8475] <= 8'h00;
            reg_file[8476] <= 8'h6F;
            reg_file[8477] <= 8'hF0;
            reg_file[8478] <= 8'h9F;
            reg_file[8479] <= 8'hF0;
            reg_file[8480] <= 8'h13;
            reg_file[8481] <= 8'h04;
            reg_file[8482] <= 8'h00;
            reg_file[8483] <= 8'h00;
            reg_file[8484] <= 8'h93;
            reg_file[8485] <= 8'h07;
            reg_file[8486] <= 8'h00;
            reg_file[8487] <= 8'h00;
            reg_file[8488] <= 8'h13;
            reg_file[8489] <= 8'h05;
            reg_file[8490] <= 8'hF0;
            reg_file[8491] <= 8'h7F;
            reg_file[8492] <= 8'h13;
            reg_file[8493] <= 8'h07;
            reg_file[8494] <= 8'h20;
            reg_file[8495] <= 8'h00;
            reg_file[8496] <= 8'h6F;
            reg_file[8497] <= 8'hF0;
            reg_file[8498] <= 8'h5F;
            reg_file[8499] <= 8'hEF;
            reg_file[8500] <= 8'h13;
            reg_file[8501] <= 8'h07;
            reg_file[8502] <= 8'h30;
            reg_file[8503] <= 8'h00;
            reg_file[8504] <= 8'h6F;
            reg_file[8505] <= 8'hF0;
            reg_file[8506] <= 8'hDF;
            reg_file[8507] <= 8'hEE;
            reg_file[8508] <= 8'h37;
            reg_file[8509] <= 8'h04;
            reg_file[8510] <= 8'h08;
            reg_file[8511] <= 8'h00;
            reg_file[8512] <= 8'h93;
            reg_file[8513] <= 8'h07;
            reg_file[8514] <= 8'h00;
            reg_file[8515] <= 8'h00;
            reg_file[8516] <= 8'h13;
            reg_file[8517] <= 8'h07;
            reg_file[8518] <= 8'hF0;
            reg_file[8519] <= 8'h7F;
            reg_file[8520] <= 8'h93;
            reg_file[8521] <= 8'h05;
            reg_file[8522] <= 8'h00;
            reg_file[8523] <= 8'h00;
            reg_file[8524] <= 8'h93;
            reg_file[8525] <= 8'h04;
            reg_file[8526] <= 8'h00;
            reg_file[8527] <= 8'h01;
            reg_file[8528] <= 8'h13;
            reg_file[8529] <= 8'h17;
            reg_file[8530] <= 8'h47;
            reg_file[8531] <= 8'h01;
            reg_file[8532] <= 8'hB7;
            reg_file[8533] <= 8'h06;
            reg_file[8534] <= 8'hF0;
            reg_file[8535] <= 8'h7F;
            reg_file[8536] <= 8'h13;
            reg_file[8537] <= 8'h14;
            reg_file[8538] <= 8'hC4;
            reg_file[8539] <= 8'h00;
            reg_file[8540] <= 8'h33;
            reg_file[8541] <= 8'h77;
            reg_file[8542] <= 8'hD7;
            reg_file[8543] <= 8'h00;
            reg_file[8544] <= 8'h13;
            reg_file[8545] <= 8'h54;
            reg_file[8546] <= 8'hC4;
            reg_file[8547] <= 8'h00;
            reg_file[8548] <= 8'h93;
            reg_file[8549] <= 8'h95;
            reg_file[8550] <= 8'hF5;
            reg_file[8551] <= 8'h01;
            reg_file[8552] <= 8'h33;
            reg_file[8553] <= 8'h64;
            reg_file[8554] <= 8'h87;
            reg_file[8555] <= 8'h00;
            reg_file[8556] <= 8'h33;
            reg_file[8557] <= 8'h67;
            reg_file[8558] <= 8'hB4;
            reg_file[8559] <= 8'h00;
            reg_file[8560] <= 8'h13;
            reg_file[8561] <= 8'h85;
            reg_file[8562] <= 8'h07;
            reg_file[8563] <= 8'h00;
            reg_file[8564] <= 8'h93;
            reg_file[8565] <= 8'h05;
            reg_file[8566] <= 8'h07;
            reg_file[8567] <= 8'h00;
            reg_file[8568] <= 8'h63;
            reg_file[8569] <= 8'h84;
            reg_file[8570] <= 8'h04;
            reg_file[8571] <= 8'h00;
            reg_file[8572] <= 8'h73;
            reg_file[8573] <= 8'hA0;
            reg_file[8574] <= 8'h14;
            reg_file[8575] <= 8'h00;
            reg_file[8576] <= 8'h83;
            reg_file[8577] <= 8'h20;
            reg_file[8578] <= 8'hC1;
            reg_file[8579] <= 8'h02;
            reg_file[8580] <= 8'h03;
            reg_file[8581] <= 8'h24;
            reg_file[8582] <= 8'h81;
            reg_file[8583] <= 8'h02;
            reg_file[8584] <= 8'h83;
            reg_file[8585] <= 8'h24;
            reg_file[8586] <= 8'h41;
            reg_file[8587] <= 8'h02;
            reg_file[8588] <= 8'h03;
            reg_file[8589] <= 8'h29;
            reg_file[8590] <= 8'h01;
            reg_file[8591] <= 8'h02;
            reg_file[8592] <= 8'h83;
            reg_file[8593] <= 8'h29;
            reg_file[8594] <= 8'hC1;
            reg_file[8595] <= 8'h01;
            reg_file[8596] <= 8'h03;
            reg_file[8597] <= 8'h2A;
            reg_file[8598] <= 8'h81;
            reg_file[8599] <= 8'h01;
            reg_file[8600] <= 8'h83;
            reg_file[8601] <= 8'h2A;
            reg_file[8602] <= 8'h41;
            reg_file[8603] <= 8'h01;
            reg_file[8604] <= 8'h03;
            reg_file[8605] <= 8'h2B;
            reg_file[8606] <= 8'h01;
            reg_file[8607] <= 8'h01;
            reg_file[8608] <= 8'h83;
            reg_file[8609] <= 8'h2B;
            reg_file[8610] <= 8'hC1;
            reg_file[8611] <= 8'h00;
            reg_file[8612] <= 8'h03;
            reg_file[8613] <= 8'h2C;
            reg_file[8614] <= 8'h81;
            reg_file[8615] <= 8'h00;
            reg_file[8616] <= 8'h83;
            reg_file[8617] <= 8'h2C;
            reg_file[8618] <= 8'h41;
            reg_file[8619] <= 8'h00;
            reg_file[8620] <= 8'h13;
            reg_file[8621] <= 8'h01;
            reg_file[8622] <= 8'h01;
            reg_file[8623] <= 8'h03;
            reg_file[8624] <= 8'h67;
            reg_file[8625] <= 8'h80;
            reg_file[8626] <= 8'h00;
            reg_file[8627] <= 8'h00;
            reg_file[8628] <= 8'h37;
            reg_file[8629] <= 8'h06;
            reg_file[8630] <= 8'h01;
            reg_file[8631] <= 8'h00;
            reg_file[8632] <= 8'h13;
            reg_file[8633] <= 8'h07;
            reg_file[8634] <= 8'hF6;
            reg_file[8635] <= 8'hFF;
            reg_file[8636] <= 8'h93;
            reg_file[8637] <= 8'h56;
            reg_file[8638] <= 8'h0A;
            reg_file[8639] <= 8'h01;
            reg_file[8640] <= 8'h13;
            reg_file[8641] <= 8'hDE;
            reg_file[8642] <= 8'h07;
            reg_file[8643] <= 8'h01;
            reg_file[8644] <= 8'h33;
            reg_file[8645] <= 8'h7A;
            reg_file[8646] <= 8'hEA;
            reg_file[8647] <= 8'h00;
            reg_file[8648] <= 8'hB3;
            reg_file[8649] <= 8'hF7;
            reg_file[8650] <= 8'hE7;
            reg_file[8651] <= 8'h00;
            reg_file[8652] <= 8'h33;
            reg_file[8653] <= 8'h03;
            reg_file[8654] <= 8'h4E;
            reg_file[8655] <= 8'h03;
            reg_file[8656] <= 8'hB3;
            reg_file[8657] <= 8'h8E;
            reg_file[8658] <= 8'h47;
            reg_file[8659] <= 8'h03;
            reg_file[8660] <= 8'h33;
            reg_file[8661] <= 8'h8F;
            reg_file[8662] <= 8'hF6;
            reg_file[8663] <= 8'h02;
            reg_file[8664] <= 8'h33;
            reg_file[8665] <= 8'h08;
            reg_file[8666] <= 8'hE3;
            reg_file[8667] <= 8'h01;
            reg_file[8668] <= 8'h13;
            reg_file[8669] <= 8'hD3;
            reg_file[8670] <= 8'h0E;
            reg_file[8671] <= 8'h01;
            reg_file[8672] <= 8'h33;
            reg_file[8673] <= 8'h03;
            reg_file[8674] <= 8'h03;
            reg_file[8675] <= 8'h01;
            reg_file[8676] <= 8'hB3;
            reg_file[8677] <= 8'h88;
            reg_file[8678] <= 8'hC6;
            reg_file[8679] <= 8'h03;
            reg_file[8680] <= 8'h63;
            reg_file[8681] <= 8'h74;
            reg_file[8682] <= 8'hE3;
            reg_file[8683] <= 8'h01;
            reg_file[8684] <= 8'hB3;
            reg_file[8685] <= 8'h88;
            reg_file[8686] <= 8'hC8;
            reg_file[8687] <= 8'h00;
            reg_file[8688] <= 8'h33;
            reg_file[8689] <= 8'h78;
            reg_file[8690] <= 8'hE3;
            reg_file[8691] <= 8'h00;
            reg_file[8692] <= 8'hB3;
            reg_file[8693] <= 8'hFE;
            reg_file[8694] <= 8'hEE;
            reg_file[8695] <= 8'h00;
            reg_file[8696] <= 8'h13;
            reg_file[8697] <= 8'h56;
            reg_file[8698] <= 8'h03;
            reg_file[8699] <= 8'h01;
            reg_file[8700] <= 8'h13;
            reg_file[8701] <= 8'h18;
            reg_file[8702] <= 8'h08;
            reg_file[8703] <= 8'h01;
            reg_file[8704] <= 8'h13;
            reg_file[8705] <= 8'h53;
            reg_file[8706] <= 8'h04;
            reg_file[8707] <= 8'h01;
            reg_file[8708] <= 8'h33;
            reg_file[8709] <= 8'h74;
            reg_file[8710] <= 8'hE4;
            reg_file[8711] <= 8'h00;
            reg_file[8712] <= 8'h33;
            reg_file[8713] <= 8'h08;
            reg_file[8714] <= 8'hD8;
            reg_file[8715] <= 8'h01;
            reg_file[8716] <= 8'h33;
            reg_file[8717] <= 8'h0F;
            reg_file[8718] <= 8'h8A;
            reg_file[8719] <= 8'h02;
            reg_file[8720] <= 8'hB3;
            reg_file[8721] <= 8'h8E;
            reg_file[8722] <= 8'h86;
            reg_file[8723] <= 8'h02;
            reg_file[8724] <= 8'h33;
            reg_file[8725] <= 8'h0A;
            reg_file[8726] <= 8'h43;
            reg_file[8727] <= 8'h03;
            reg_file[8728] <= 8'h33;
            reg_file[8729] <= 8'h07;
            reg_file[8730] <= 8'hDA;
            reg_file[8731] <= 8'h01;
            reg_file[8732] <= 8'h13;
            reg_file[8733] <= 8'h5A;
            reg_file[8734] <= 8'h0F;
            reg_file[8735] <= 8'h01;
            reg_file[8736] <= 8'h33;
            reg_file[8737] <= 8'h0A;
            reg_file[8738] <= 8'hEA;
            reg_file[8739] <= 8'h00;
            reg_file[8740] <= 8'hB3;
            reg_file[8741] <= 8'h86;
            reg_file[8742] <= 8'h66;
            reg_file[8743] <= 8'h02;
            reg_file[8744] <= 8'h63;
            reg_file[8745] <= 8'h76;
            reg_file[8746] <= 8'hDA;
            reg_file[8747] <= 8'h01;
            reg_file[8748] <= 8'h37;
            reg_file[8749] <= 8'h07;
            reg_file[8750] <= 8'h01;
            reg_file[8751] <= 8'h00;
            reg_file[8752] <= 8'hB3;
            reg_file[8753] <= 8'h86;
            reg_file[8754] <= 8'hE6;
            reg_file[8755] <= 8'h00;
            reg_file[8756] <= 8'h93;
            reg_file[8757] <= 8'h5E;
            reg_file[8758] <= 8'h0A;
            reg_file[8759] <= 8'h01;
            reg_file[8760] <= 8'hB3;
            reg_file[8761] <= 8'h8E;
            reg_file[8762] <= 8'hDE;
            reg_file[8763] <= 8'h00;
            reg_file[8764] <= 8'hB7;
            reg_file[8765] <= 8'h06;
            reg_file[8766] <= 8'h01;
            reg_file[8767] <= 8'h00;
            reg_file[8768] <= 8'h93;
            reg_file[8769] <= 8'h82;
            reg_file[8770] <= 8'hF6;
            reg_file[8771] <= 8'hFF;
            reg_file[8772] <= 8'h33;
            reg_file[8773] <= 8'h7A;
            reg_file[8774] <= 8'h5A;
            reg_file[8775] <= 8'h00;
            reg_file[8776] <= 8'h33;
            reg_file[8777] <= 8'h7F;
            reg_file[8778] <= 8'h5F;
            reg_file[8779] <= 8'h00;
            reg_file[8780] <= 8'h13;
            reg_file[8781] <= 8'hD7;
            reg_file[8782] <= 8'h09;
            reg_file[8783] <= 8'h01;
            reg_file[8784] <= 8'h13;
            reg_file[8785] <= 8'h1A;
            reg_file[8786] <= 8'h0A;
            reg_file[8787] <= 8'h01;
            reg_file[8788] <= 8'hB3;
            reg_file[8789] <= 8'hF9;
            reg_file[8790] <= 8'h59;
            reg_file[8791] <= 8'h00;
            reg_file[8792] <= 8'h33;
            reg_file[8793] <= 8'h0A;
            reg_file[8794] <= 8'hEA;
            reg_file[8795] <= 8'h01;
            reg_file[8796] <= 8'hB3;
            reg_file[8797] <= 8'h02;
            reg_file[8798] <= 8'hEE;
            reg_file[8799] <= 8'h02;
            reg_file[8800] <= 8'hB3;
            reg_file[8801] <= 8'h0F;
            reg_file[8802] <= 8'h46;
            reg_file[8803] <= 8'h01;
            reg_file[8804] <= 8'h33;
            reg_file[8805] <= 8'h8F;
            reg_file[8806] <= 8'h37;
            reg_file[8807] <= 8'h03;
            reg_file[8808] <= 8'h33;
            reg_file[8809] <= 8'h0E;
            reg_file[8810] <= 8'h3E;
            reg_file[8811] <= 8'h03;
            reg_file[8812] <= 8'h13;
            reg_file[8813] <= 8'h56;
            reg_file[8814] <= 8'h0F;
            reg_file[8815] <= 8'h01;
            reg_file[8816] <= 8'hB3;
            reg_file[8817] <= 8'h07;
            reg_file[8818] <= 8'hF7;
            reg_file[8819] <= 8'h02;
            reg_file[8820] <= 8'h33;
            reg_file[8821] <= 8'h0E;
            reg_file[8822] <= 8'hFE;
            reg_file[8823] <= 8'h00;
            reg_file[8824] <= 8'h33;
            reg_file[8825] <= 8'h06;
            reg_file[8826] <= 8'hC6;
            reg_file[8827] <= 8'h01;
            reg_file[8828] <= 8'h63;
            reg_file[8829] <= 8'h74;
            reg_file[8830] <= 8'hF6;
            reg_file[8831] <= 8'h00;
            reg_file[8832] <= 8'hB3;
            reg_file[8833] <= 8'h82;
            reg_file[8834] <= 8'hD2;
            reg_file[8835] <= 8'h00;
            reg_file[8836] <= 8'hB7;
            reg_file[8837] <= 8'h06;
            reg_file[8838] <= 8'h01;
            reg_file[8839] <= 8'h00;
            reg_file[8840] <= 8'h93;
            reg_file[8841] <= 8'h87;
            reg_file[8842] <= 8'hF6;
            reg_file[8843] <= 8'hFF;
            reg_file[8844] <= 8'h13;
            reg_file[8845] <= 8'h5E;
            reg_file[8846] <= 8'h06;
            reg_file[8847] <= 8'h01;
            reg_file[8848] <= 8'h33;
            reg_file[8849] <= 8'h76;
            reg_file[8850] <= 8'hF6;
            reg_file[8851] <= 8'h00;
            reg_file[8852] <= 8'h33;
            reg_file[8853] <= 8'h7F;
            reg_file[8854] <= 8'hFF;
            reg_file[8855] <= 8'h00;
            reg_file[8856] <= 8'h13;
            reg_file[8857] <= 8'h16;
            reg_file[8858] <= 8'h06;
            reg_file[8859] <= 8'h01;
            reg_file[8860] <= 8'hB3;
            reg_file[8861] <= 8'h87;
            reg_file[8862] <= 8'h89;
            reg_file[8863] <= 8'h02;
            reg_file[8864] <= 8'h33;
            reg_file[8865] <= 8'h06;
            reg_file[8866] <= 8'hE6;
            reg_file[8867] <= 8'h01;
            reg_file[8868] <= 8'h33;
            reg_file[8869] <= 8'h0E;
            reg_file[8870] <= 8'h5E;
            reg_file[8871] <= 8'h00;
            reg_file[8872] <= 8'h33;
            reg_file[8873] <= 8'h04;
            reg_file[8874] <= 8'h87;
            reg_file[8875] <= 8'h02;
            reg_file[8876] <= 8'h33;
            reg_file[8877] <= 8'h0F;
            reg_file[8878] <= 8'hE3;
            reg_file[8879] <= 8'h02;
            reg_file[8880] <= 8'h13;
            reg_file[8881] <= 8'hD7;
            reg_file[8882] <= 8'h07;
            reg_file[8883] <= 8'h01;
            reg_file[8884] <= 8'h33;
            reg_file[8885] <= 8'h03;
            reg_file[8886] <= 8'h33;
            reg_file[8887] <= 8'h03;
            reg_file[8888] <= 8'h33;
            reg_file[8889] <= 8'h03;
            reg_file[8890] <= 8'h83;
            reg_file[8891] <= 8'h00;
            reg_file[8892] <= 8'h33;
            reg_file[8893] <= 8'h03;
            reg_file[8894] <= 8'h67;
            reg_file[8895] <= 8'h00;
            reg_file[8896] <= 8'h63;
            reg_file[8897] <= 8'h74;
            reg_file[8898] <= 8'h83;
            reg_file[8899] <= 8'h00;
            reg_file[8900] <= 8'h33;
            reg_file[8901] <= 8'h0F;
            reg_file[8902] <= 8'hDF;
            reg_file[8903] <= 8'h00;
            reg_file[8904] <= 8'h37;
            reg_file[8905] <= 8'h07;
            reg_file[8906] <= 8'h01;
            reg_file[8907] <= 8'h00;
            reg_file[8908] <= 8'h13;
            reg_file[8909] <= 8'h07;
            reg_file[8910] <= 8'hF7;
            reg_file[8911] <= 8'hFF;
            reg_file[8912] <= 8'hB3;
            reg_file[8913] <= 8'h76;
            reg_file[8914] <= 8'hE3;
            reg_file[8915] <= 8'h00;
            reg_file[8916] <= 8'hB3;
            reg_file[8917] <= 8'hF7;
            reg_file[8918] <= 8'hE7;
            reg_file[8919] <= 8'h00;
            reg_file[8920] <= 8'h93;
            reg_file[8921] <= 8'h96;
            reg_file[8922] <= 8'h06;
            reg_file[8923] <= 8'h01;
            reg_file[8924] <= 8'hB3;
            reg_file[8925] <= 8'h88;
            reg_file[8926] <= 8'hF8;
            reg_file[8927] <= 8'h01;
            reg_file[8928] <= 8'hB3;
            reg_file[8929] <= 8'h86;
            reg_file[8930] <= 8'hF6;
            reg_file[8931] <= 8'h00;
            reg_file[8932] <= 8'h33;
            reg_file[8933] <= 8'hBA;
            reg_file[8934] <= 8'h48;
            reg_file[8935] <= 8'h01;
            reg_file[8936] <= 8'hB3;
            reg_file[8937] <= 8'h86;
            reg_file[8938] <= 8'hD6;
            reg_file[8939] <= 8'h01;
            reg_file[8940] <= 8'h33;
            reg_file[8941] <= 8'h87;
            reg_file[8942] <= 8'h46;
            reg_file[8943] <= 8'h01;
            reg_file[8944] <= 8'hB3;
            reg_file[8945] <= 8'h88;
            reg_file[8946] <= 8'hC8;
            reg_file[8947] <= 8'h00;
            reg_file[8948] <= 8'h33;
            reg_file[8949] <= 8'hB6;
            reg_file[8950] <= 8'hC8;
            reg_file[8951] <= 8'h00;
            reg_file[8952] <= 8'hB3;
            reg_file[8953] <= 8'h0F;
            reg_file[8954] <= 8'hC7;
            reg_file[8955] <= 8'h01;
            reg_file[8956] <= 8'hB3;
            reg_file[8957] <= 8'h82;
            reg_file[8958] <= 8'hCF;
            reg_file[8959] <= 8'h00;
            reg_file[8960] <= 8'hB3;
            reg_file[8961] <= 8'hB6;
            reg_file[8962] <= 8'hD6;
            reg_file[8963] <= 8'h01;
            reg_file[8964] <= 8'h33;
            reg_file[8965] <= 8'h37;
            reg_file[8966] <= 8'h47;
            reg_file[8967] <= 8'h01;
            reg_file[8968] <= 8'h33;
            reg_file[8969] <= 8'hE7;
            reg_file[8970] <= 8'hE6;
            reg_file[8971] <= 8'h00;
            reg_file[8972] <= 8'h33;
            reg_file[8973] <= 8'hB6;
            reg_file[8974] <= 8'hC2;
            reg_file[8975] <= 8'h00;
            reg_file[8976] <= 8'h13;
            reg_file[8977] <= 8'h53;
            reg_file[8978] <= 8'h03;
            reg_file[8979] <= 8'h01;
            reg_file[8980] <= 8'h33;
            reg_file[8981] <= 8'hBE;
            reg_file[8982] <= 8'hCF;
            reg_file[8983] <= 8'h01;
            reg_file[8984] <= 8'h33;
            reg_file[8985] <= 8'h07;
            reg_file[8986] <= 8'h67;
            reg_file[8987] <= 8'h00;
            reg_file[8988] <= 8'h33;
            reg_file[8989] <= 8'h66;
            reg_file[8990] <= 8'hCE;
            reg_file[8991] <= 8'h00;
            reg_file[8992] <= 8'h93;
            reg_file[8993] <= 8'h97;
            reg_file[8994] <= 8'h98;
            reg_file[8995] <= 8'h00;
            reg_file[8996] <= 8'h33;
            reg_file[8997] <= 8'h07;
            reg_file[8998] <= 8'hC7;
            reg_file[8999] <= 8'h00;
            reg_file[9000] <= 8'h33;
            reg_file[9001] <= 8'h07;
            reg_file[9002] <= 8'hE7;
            reg_file[9003] <= 8'h01;
            reg_file[9004] <= 8'hB3;
            reg_file[9005] <= 8'hE7;
            reg_file[9006] <= 8'h07;
            reg_file[9007] <= 8'h01;
            reg_file[9008] <= 8'h13;
            reg_file[9009] <= 8'h17;
            reg_file[9010] <= 8'h97;
            reg_file[9011] <= 8'h00;
            reg_file[9012] <= 8'hB3;
            reg_file[9013] <= 8'h37;
            reg_file[9014] <= 8'hF0;
            reg_file[9015] <= 8'h00;
            reg_file[9016] <= 8'h93;
            reg_file[9017] <= 8'hD8;
            reg_file[9018] <= 8'h78;
            reg_file[9019] <= 8'h01;
            reg_file[9020] <= 8'h13;
            reg_file[9021] <= 8'hD4;
            reg_file[9022] <= 8'h72;
            reg_file[9023] <= 8'h01;
            reg_file[9024] <= 8'hB3;
            reg_file[9025] <= 8'hE7;
            reg_file[9026] <= 8'h17;
            reg_file[9027] <= 8'h01;
            reg_file[9028] <= 8'h93;
            reg_file[9029] <= 8'h92;
            reg_file[9030] <= 8'h92;
            reg_file[9031] <= 8'h00;
            reg_file[9032] <= 8'h93;
            reg_file[9033] <= 8'h16;
            reg_file[9034] <= 8'h77;
            reg_file[9035] <= 8'h00;
            reg_file[9036] <= 8'h33;
            reg_file[9037] <= 8'h64;
            reg_file[9038] <= 8'h87;
            reg_file[9039] <= 8'h00;
            reg_file[9040] <= 8'hB3;
            reg_file[9041] <= 8'hE7;
            reg_file[9042] <= 8'h57;
            reg_file[9043] <= 8'h00;
            reg_file[9044] <= 8'h63;
            reg_file[9045] <= 8'hD0;
            reg_file[9046] <= 8'h06;
            reg_file[9047] <= 8'h0A;
            reg_file[9048] <= 8'h13;
            reg_file[9049] <= 8'hD7;
            reg_file[9050] <= 8'h17;
            reg_file[9051] <= 8'h00;
            reg_file[9052] <= 8'h93;
            reg_file[9053] <= 8'hF7;
            reg_file[9054] <= 8'h17;
            reg_file[9055] <= 8'h00;
            reg_file[9056] <= 8'hB3;
            reg_file[9057] <= 8'h67;
            reg_file[9058] <= 8'hF7;
            reg_file[9059] <= 8'h00;
            reg_file[9060] <= 8'h13;
            reg_file[9061] <= 8'h17;
            reg_file[9062] <= 8'hF4;
            reg_file[9063] <= 8'h01;
            reg_file[9064] <= 8'hB3;
            reg_file[9065] <= 8'hE7;
            reg_file[9066] <= 8'hE7;
            reg_file[9067] <= 8'h00;
            reg_file[9068] <= 8'h13;
            reg_file[9069] <= 8'h54;
            reg_file[9070] <= 8'h14;
            reg_file[9071] <= 8'h00;
            reg_file[9072] <= 8'h13;
            reg_file[9073] <= 8'h08;
            reg_file[9074] <= 8'hF5;
            reg_file[9075] <= 8'h3F;
            reg_file[9076] <= 8'h63;
            reg_file[9077] <= 8'h58;
            reg_file[9078] <= 8'h00;
            reg_file[9079] <= 8'h11;
            reg_file[9080] <= 8'h13;
            reg_file[9081] <= 8'hF7;
            reg_file[9082] <= 8'h77;
            reg_file[9083] <= 8'h00;
            reg_file[9084] <= 8'h63;
            reg_file[9085] <= 8'h08;
            reg_file[9086] <= 8'h07;
            reg_file[9087] <= 8'h08;
            reg_file[9088] <= 8'h13;
            reg_file[9089] <= 8'h07;
            reg_file[9090] <= 8'h20;
            reg_file[9091] <= 8'h00;
            reg_file[9092] <= 8'h93;
            reg_file[9093] <= 8'hE4;
            reg_file[9094] <= 8'h14;
            reg_file[9095] <= 8'h00;
            reg_file[9096] <= 8'h63;
            reg_file[9097] <= 8'h00;
            reg_file[9098] <= 8'hE9;
            reg_file[9099] <= 8'h08;
            reg_file[9100] <= 8'h13;
            reg_file[9101] <= 8'h07;
            reg_file[9102] <= 8'h30;
            reg_file[9103] <= 8'h00;
            reg_file[9104] <= 8'h63;
            reg_file[9105] <= 8'h06;
            reg_file[9106] <= 8'hE9;
            reg_file[9107] <= 8'h06;
            reg_file[9108] <= 8'h63;
            reg_file[9109] <= 8'h1C;
            reg_file[9110] <= 8'h09;
            reg_file[9111] <= 8'h06;
            reg_file[9112] <= 8'h13;
            reg_file[9113] <= 8'hF7;
            reg_file[9114] <= 8'hF7;
            reg_file[9115] <= 8'h00;
            reg_file[9116] <= 8'h93;
            reg_file[9117] <= 8'h06;
            reg_file[9118] <= 8'h40;
            reg_file[9119] <= 8'h00;
            reg_file[9120] <= 8'h63;
            reg_file[9121] <= 8'h06;
            reg_file[9122] <= 8'hD7;
            reg_file[9123] <= 8'h06;
            reg_file[9124] <= 8'h13;
            reg_file[9125] <= 8'h87;
            reg_file[9126] <= 8'h47;
            reg_file[9127] <= 8'h00;
            reg_file[9128] <= 8'hB3;
            reg_file[9129] <= 8'h37;
            reg_file[9130] <= 8'hF7;
            reg_file[9131] <= 8'h00;
            reg_file[9132] <= 8'h33;
            reg_file[9133] <= 8'h04;
            reg_file[9134] <= 8'hF4;
            reg_file[9135] <= 8'h00;
            reg_file[9136] <= 8'h93;
            reg_file[9137] <= 8'h07;
            reg_file[9138] <= 8'h07;
            reg_file[9139] <= 8'h00;
            reg_file[9140] <= 8'h6F;
            reg_file[9141] <= 8'h00;
            reg_file[9142] <= 8'h80;
            reg_file[9143] <= 8'h05;
            reg_file[9144] <= 8'h93;
            reg_file[9145] <= 8'h85;
            reg_file[9146] <= 8'h0A;
            reg_file[9147] <= 8'h00;
            reg_file[9148] <= 8'h13;
            reg_file[9149] <= 8'h84;
            reg_file[9150] <= 8'h09;
            reg_file[9151] <= 8'h00;
            reg_file[9152] <= 8'h93;
            reg_file[9153] <= 8'h07;
            reg_file[9154] <= 8'h0A;
            reg_file[9155] <= 8'h00;
            reg_file[9156] <= 8'h13;
            reg_file[9157] <= 8'h07;
            reg_file[9158] <= 8'h0C;
            reg_file[9159] <= 8'h00;
            reg_file[9160] <= 8'h93;
            reg_file[9161] <= 8'h06;
            reg_file[9162] <= 8'h20;
            reg_file[9163] <= 8'h00;
            reg_file[9164] <= 8'h63;
            reg_file[9165] <= 8'h02;
            reg_file[9166] <= 8'hD7;
            reg_file[9167] <= 8'h28;
            reg_file[9168] <= 8'h93;
            reg_file[9169] <= 8'h06;
            reg_file[9170] <= 8'h30;
            reg_file[9171] <= 8'h00;
            reg_file[9172] <= 8'h63;
            reg_file[9173] <= 8'h06;
            reg_file[9174] <= 8'hD7;
            reg_file[9175] <= 8'h28;
            reg_file[9176] <= 8'h93;
            reg_file[9177] <= 8'h06;
            reg_file[9178] <= 8'h10;
            reg_file[9179] <= 8'h00;
            reg_file[9180] <= 8'hE3;
            reg_file[9181] <= 8'h1A;
            reg_file[9182] <= 8'hD7;
            reg_file[9183] <= 8'hF8;
            reg_file[9184] <= 8'h13;
            reg_file[9185] <= 8'h04;
            reg_file[9186] <= 8'h00;
            reg_file[9187] <= 8'h00;
            reg_file[9188] <= 8'h93;
            reg_file[9189] <= 8'h07;
            reg_file[9190] <= 8'h00;
            reg_file[9191] <= 8'h00;
            reg_file[9192] <= 8'h6F;
            reg_file[9193] <= 8'h00;
            reg_file[9194] <= 8'h40;
            reg_file[9195] <= 8'h24;
            reg_file[9196] <= 8'h93;
            reg_file[9197] <= 8'h05;
            reg_file[9198] <= 8'h0B;
            reg_file[9199] <= 8'h00;
            reg_file[9200] <= 8'h6F;
            reg_file[9201] <= 8'hF0;
            reg_file[9202] <= 8'h9F;
            reg_file[9203] <= 8'hFD;
            reg_file[9204] <= 8'h13;
            reg_file[9205] <= 8'h85;
            reg_file[9206] <= 8'h0B;
            reg_file[9207] <= 8'h00;
            reg_file[9208] <= 8'h6F;
            reg_file[9209] <= 8'hF0;
            reg_file[9210] <= 8'h9F;
            reg_file[9211] <= 8'hF7;
            reg_file[9212] <= 8'h63;
            reg_file[9213] <= 8'h98;
            reg_file[9214] <= 8'h05;
            reg_file[9215] <= 8'h00;
            reg_file[9216] <= 8'h13;
            reg_file[9217] <= 8'h87;
            reg_file[9218] <= 8'h87;
            reg_file[9219] <= 8'h00;
            reg_file[9220] <= 8'h6F;
            reg_file[9221] <= 8'hF0;
            reg_file[9222] <= 8'h5F;
            reg_file[9223] <= 8'hFA;
            reg_file[9224] <= 8'hE3;
            reg_file[9225] <= 8'h9C;
            reg_file[9226] <= 8'h05;
            reg_file[9227] <= 8'hFE;
            reg_file[9228] <= 8'h13;
            reg_file[9229] <= 8'h17;
            reg_file[9230] <= 8'h74;
            reg_file[9231] <= 8'h00;
            reg_file[9232] <= 8'h63;
            reg_file[9233] <= 8'h5A;
            reg_file[9234] <= 8'h07;
            reg_file[9235] <= 8'h00;
            reg_file[9236] <= 8'h37;
            reg_file[9237] <= 8'h07;
            reg_file[9238] <= 8'h00;
            reg_file[9239] <= 8'hFF;
            reg_file[9240] <= 8'h13;
            reg_file[9241] <= 8'h07;
            reg_file[9242] <= 8'hF7;
            reg_file[9243] <= 8'hFF;
            reg_file[9244] <= 8'h33;
            reg_file[9245] <= 8'h74;
            reg_file[9246] <= 8'hE4;
            reg_file[9247] <= 8'h00;
            reg_file[9248] <= 8'h13;
            reg_file[9249] <= 8'h08;
            reg_file[9250] <= 8'h05;
            reg_file[9251] <= 8'h40;
            reg_file[9252] <= 8'h13;
            reg_file[9253] <= 8'h07;
            reg_file[9254] <= 8'hE0;
            reg_file[9255] <= 8'h7F;
            reg_file[9256] <= 8'h63;
            reg_file[9257] <= 8'h4E;
            reg_file[9258] <= 8'h07;
            reg_file[9259] <= 8'h01;
            reg_file[9260] <= 8'h13;
            reg_file[9261] <= 8'hD7;
            reg_file[9262] <= 8'h37;
            reg_file[9263] <= 8'h00;
            reg_file[9264] <= 8'h93;
            reg_file[9265] <= 8'h17;
            reg_file[9266] <= 8'hD4;
            reg_file[9267] <= 8'h01;
            reg_file[9268] <= 8'hB3;
            reg_file[9269] <= 8'hE7;
            reg_file[9270] <= 8'hE7;
            reg_file[9271] <= 8'h00;
            reg_file[9272] <= 8'h13;
            reg_file[9273] <= 8'h54;
            reg_file[9274] <= 8'h34;
            reg_file[9275] <= 8'h00;
            reg_file[9276] <= 8'h13;
            reg_file[9277] <= 8'h07;
            reg_file[9278] <= 8'h08;
            reg_file[9279] <= 8'h00;
            reg_file[9280] <= 8'h6F;
            reg_file[9281] <= 8'hF0;
            reg_file[9282] <= 8'h1F;
            reg_file[9283] <= 8'hD1;
            reg_file[9284] <= 8'h93;
            reg_file[9285] <= 8'h07;
            reg_file[9286] <= 8'h20;
            reg_file[9287] <= 8'h00;
            reg_file[9288] <= 8'h63;
            reg_file[9289] <= 8'h0A;
            reg_file[9290] <= 8'hF9;
            reg_file[9291] <= 8'h02;
            reg_file[9292] <= 8'h93;
            reg_file[9293] <= 8'h07;
            reg_file[9294] <= 8'h30;
            reg_file[9295] <= 8'h00;
            reg_file[9296] <= 8'h63;
            reg_file[9297] <= 8'h0A;
            reg_file[9298] <= 8'hF9;
            reg_file[9299] <= 8'h00;
            reg_file[9300] <= 8'h63;
            reg_file[9301] <= 8'h1A;
            reg_file[9302] <= 8'h09;
            reg_file[9303] <= 8'h00;
            reg_file[9304] <= 8'h93;
            reg_file[9305] <= 8'h07;
            reg_file[9306] <= 8'h00;
            reg_file[9307] <= 8'h00;
            reg_file[9308] <= 8'h13;
            reg_file[9309] <= 8'h07;
            reg_file[9310] <= 8'hF0;
            reg_file[9311] <= 8'h7F;
            reg_file[9312] <= 8'h6F;
            reg_file[9313] <= 8'h00;
            reg_file[9314] <= 8'h00;
            reg_file[9315] <= 8'h01;
            reg_file[9316] <= 8'hE3;
            reg_file[9317] <= 8'h8A;
            reg_file[9318] <= 8'h05;
            reg_file[9319] <= 8'hFE;
            reg_file[9320] <= 8'h93;
            reg_file[9321] <= 8'h07;
            reg_file[9322] <= 8'hF0;
            reg_file[9323] <= 8'hFF;
            reg_file[9324] <= 8'h13;
            reg_file[9325] <= 8'h07;
            reg_file[9326] <= 8'hE0;
            reg_file[9327] <= 8'h7F;
            reg_file[9328] <= 8'h93;
            reg_file[9329] <= 8'hE4;
            reg_file[9330] <= 8'h54;
            reg_file[9331] <= 8'h00;
            reg_file[9332] <= 8'h13;
            reg_file[9333] <= 8'h84;
            reg_file[9334] <= 8'h07;
            reg_file[9335] <= 8'h00;
            reg_file[9336] <= 8'h6F;
            reg_file[9337] <= 8'hF0;
            reg_file[9338] <= 8'h9F;
            reg_file[9339] <= 8'hCD;
            reg_file[9340] <= 8'hE3;
            reg_file[9341] <= 8'h9E;
            reg_file[9342] <= 8'h05;
            reg_file[9343] <= 8'hFC;
            reg_file[9344] <= 8'h6F;
            reg_file[9345] <= 8'hF0;
            reg_file[9346] <= 8'h9F;
            reg_file[9347] <= 8'hFE;
            reg_file[9348] <= 8'h13;
            reg_file[9349] <= 8'h07;
            reg_file[9350] <= 8'h10;
            reg_file[9351] <= 8'h00;
            reg_file[9352] <= 8'h63;
            reg_file[9353] <= 8'h16;
            reg_file[9354] <= 8'h08;
            reg_file[9355] <= 8'h06;
            reg_file[9356] <= 8'h93;
            reg_file[9357] <= 8'hF6;
            reg_file[9358] <= 8'h77;
            reg_file[9359] <= 8'h00;
            reg_file[9360] <= 8'h13;
            reg_file[9361] <= 8'h07;
            reg_file[9362] <= 8'h04;
            reg_file[9363] <= 8'h00;
            reg_file[9364] <= 8'h63;
            reg_file[9365] <= 8'h8A;
            reg_file[9366] <= 8'h06;
            reg_file[9367] <= 8'h04;
            reg_file[9368] <= 8'h13;
            reg_file[9369] <= 8'h07;
            reg_file[9370] <= 8'h20;
            reg_file[9371] <= 8'h00;
            reg_file[9372] <= 8'h93;
            reg_file[9373] <= 8'hE4;
            reg_file[9374] <= 8'h14;
            reg_file[9375] <= 8'h00;
            reg_file[9376] <= 8'h63;
            reg_file[9377] <= 8'h00;
            reg_file[9378] <= 8'hE9;
            reg_file[9379] <= 8'h04;
            reg_file[9380] <= 8'h13;
            reg_file[9381] <= 8'h07;
            reg_file[9382] <= 8'h30;
            reg_file[9383] <= 8'h00;
            reg_file[9384] <= 8'h63;
            reg_file[9385] <= 8'h04;
            reg_file[9386] <= 8'hE9;
            reg_file[9387] <= 8'h02;
            reg_file[9388] <= 8'h13;
            reg_file[9389] <= 8'h07;
            reg_file[9390] <= 8'h04;
            reg_file[9391] <= 8'h00;
            reg_file[9392] <= 8'h63;
            reg_file[9393] <= 8'h1C;
            reg_file[9394] <= 8'h09;
            reg_file[9395] <= 8'h02;
            reg_file[9396] <= 8'h93;
            reg_file[9397] <= 8'hF6;
            reg_file[9398] <= 8'hF7;
            reg_file[9399] <= 8'h00;
            reg_file[9400] <= 8'h13;
            reg_file[9401] <= 8'h06;
            reg_file[9402] <= 8'h40;
            reg_file[9403] <= 8'h00;
            reg_file[9404] <= 8'h63;
            reg_file[9405] <= 8'h86;
            reg_file[9406] <= 8'hC6;
            reg_file[9407] <= 8'h02;
            reg_file[9408] <= 8'h13;
            reg_file[9409] <= 8'hB7;
            reg_file[9410] <= 8'hC7;
            reg_file[9411] <= 8'hFF;
            reg_file[9412] <= 8'h13;
            reg_file[9413] <= 8'h47;
            reg_file[9414] <= 8'h17;
            reg_file[9415] <= 8'h00;
            reg_file[9416] <= 8'h33;
            reg_file[9417] <= 8'h07;
            reg_file[9418] <= 8'h87;
            reg_file[9419] <= 8'h00;
            reg_file[9420] <= 8'h6F;
            reg_file[9421] <= 8'h00;
            reg_file[9422] <= 8'hC0;
            reg_file[9423] <= 8'h01;
            reg_file[9424] <= 8'h13;
            reg_file[9425] <= 8'h07;
            reg_file[9426] <= 8'h04;
            reg_file[9427] <= 8'h00;
            reg_file[9428] <= 8'h63;
            reg_file[9429] <= 8'h9A;
            reg_file[9430] <= 8'h05;
            reg_file[9431] <= 8'h00;
            reg_file[9432] <= 8'h13;
            reg_file[9433] <= 8'hB7;
            reg_file[9434] <= 8'h87;
            reg_file[9435] <= 8'hFF;
            reg_file[9436] <= 8'h6F;
            reg_file[9437] <= 8'hF0;
            reg_file[9438] <= 8'h9F;
            reg_file[9439] <= 8'hFE;
            reg_file[9440] <= 8'h13;
            reg_file[9441] <= 8'h07;
            reg_file[9442] <= 8'h04;
            reg_file[9443] <= 8'h00;
            reg_file[9444] <= 8'hE3;
            reg_file[9445] <= 8'h9A;
            reg_file[9446] <= 8'h05;
            reg_file[9447] <= 8'hFE;
            reg_file[9448] <= 8'h13;
            reg_file[9449] <= 8'h57;
            reg_file[9450] <= 8'h87;
            reg_file[9451] <= 8'h01;
            reg_file[9452] <= 8'h13;
            reg_file[9453] <= 8'h47;
            reg_file[9454] <= 8'h17;
            reg_file[9455] <= 8'h00;
            reg_file[9456] <= 8'h13;
            reg_file[9457] <= 8'h77;
            reg_file[9458] <= 8'h17;
            reg_file[9459] <= 8'h00;
            reg_file[9460] <= 8'h93;
            reg_file[9461] <= 8'h06;
            reg_file[9462] <= 8'h10;
            reg_file[9463] <= 8'h00;
            reg_file[9464] <= 8'hB3;
            reg_file[9465] <= 8'h86;
            reg_file[9466] <= 8'h06;
            reg_file[9467] <= 8'h41;
            reg_file[9468] <= 8'h13;
            reg_file[9469] <= 8'h06;
            reg_file[9470] <= 8'h80;
            reg_file[9471] <= 8'h03;
            reg_file[9472] <= 8'h63;
            reg_file[9473] <= 8'h4C;
            reg_file[9474] <= 8'hD6;
            reg_file[9475] <= 8'h0E;
            reg_file[9476] <= 8'h13;
            reg_file[9477] <= 8'h06;
            reg_file[9478] <= 8'hF0;
            reg_file[9479] <= 8'h01;
            reg_file[9480] <= 8'h63;
            reg_file[9481] <= 8'h42;
            reg_file[9482] <= 8'hD6;
            reg_file[9483] <= 8'h06;
            reg_file[9484] <= 8'h13;
            reg_file[9485] <= 8'h05;
            reg_file[9486] <= 8'hE5;
            reg_file[9487] <= 8'h41;
            reg_file[9488] <= 8'h33;
            reg_file[9489] <= 8'h16;
            reg_file[9490] <= 8'hA4;
            reg_file[9491] <= 8'h00;
            reg_file[9492] <= 8'h33;
            reg_file[9493] <= 8'hD8;
            reg_file[9494] <= 8'hD7;
            reg_file[9495] <= 8'h00;
            reg_file[9496] <= 8'hB3;
            reg_file[9497] <= 8'h97;
            reg_file[9498] <= 8'hA7;
            reg_file[9499] <= 8'h00;
            reg_file[9500] <= 8'h33;
            reg_file[9501] <= 8'h66;
            reg_file[9502] <= 8'h06;
            reg_file[9503] <= 8'h01;
            reg_file[9504] <= 8'hB3;
            reg_file[9505] <= 8'h37;
            reg_file[9506] <= 8'hF0;
            reg_file[9507] <= 8'h00;
            reg_file[9508] <= 8'hB3;
            reg_file[9509] <= 8'h67;
            reg_file[9510] <= 8'hF6;
            reg_file[9511] <= 8'h00;
            reg_file[9512] <= 8'h33;
            reg_file[9513] <= 8'h54;
            reg_file[9514] <= 8'hD4;
            reg_file[9515] <= 8'h00;
            reg_file[9516] <= 8'h93;
            reg_file[9517] <= 8'hF6;
            reg_file[9518] <= 8'h77;
            reg_file[9519] <= 8'h00;
            reg_file[9520] <= 8'h63;
            reg_file[9521] <= 8'h80;
            reg_file[9522] <= 8'h06;
            reg_file[9523] <= 8'h08;
            reg_file[9524] <= 8'h93;
            reg_file[9525] <= 8'h06;
            reg_file[9526] <= 8'h20;
            reg_file[9527] <= 8'h00;
            reg_file[9528] <= 8'h93;
            reg_file[9529] <= 8'hE4;
            reg_file[9530] <= 8'h14;
            reg_file[9531] <= 8'h00;
            reg_file[9532] <= 8'h63;
            reg_file[9533] <= 8'h08;
            reg_file[9534] <= 8'hD9;
            reg_file[9535] <= 8'h06;
            reg_file[9536] <= 8'h93;
            reg_file[9537] <= 8'h06;
            reg_file[9538] <= 8'h30;
            reg_file[9539] <= 8'h00;
            reg_file[9540] <= 8'h63;
            reg_file[9541] <= 8'h0E;
            reg_file[9542] <= 8'hD9;
            reg_file[9543] <= 8'h04;
            reg_file[9544] <= 8'h63;
            reg_file[9545] <= 8'h14;
            reg_file[9546] <= 8'h09;
            reg_file[9547] <= 8'h06;
            reg_file[9548] <= 8'h93;
            reg_file[9549] <= 8'hF6;
            reg_file[9550] <= 8'hF7;
            reg_file[9551] <= 8'h00;
            reg_file[9552] <= 8'h13;
            reg_file[9553] <= 8'h06;
            reg_file[9554] <= 8'h40;
            reg_file[9555] <= 8'h00;
            reg_file[9556] <= 8'h63;
            reg_file[9557] <= 8'h8E;
            reg_file[9558] <= 8'hC6;
            reg_file[9559] <= 8'h04;
            reg_file[9560] <= 8'h93;
            reg_file[9561] <= 8'h86;
            reg_file[9562] <= 8'h47;
            reg_file[9563] <= 8'h00;
            reg_file[9564] <= 8'hB3;
            reg_file[9565] <= 8'hB7;
            reg_file[9566] <= 8'hF6;
            reg_file[9567] <= 8'h00;
            reg_file[9568] <= 8'h33;
            reg_file[9569] <= 8'h04;
            reg_file[9570] <= 8'hF4;
            reg_file[9571] <= 8'h00;
            reg_file[9572] <= 8'h93;
            reg_file[9573] <= 8'h87;
            reg_file[9574] <= 8'h06;
            reg_file[9575] <= 8'h00;
            reg_file[9576] <= 8'h6F;
            reg_file[9577] <= 8'h00;
            reg_file[9578] <= 8'h80;
            reg_file[9579] <= 8'h04;
            reg_file[9580] <= 8'h13;
            reg_file[9581] <= 8'h06;
            reg_file[9582] <= 8'h10;
            reg_file[9583] <= 8'hFE;
            reg_file[9584] <= 8'h33;
            reg_file[9585] <= 8'h06;
            reg_file[9586] <= 8'h06;
            reg_file[9587] <= 8'h41;
            reg_file[9588] <= 8'h93;
            reg_file[9589] <= 8'h08;
            reg_file[9590] <= 8'h00;
            reg_file[9591] <= 8'h02;
            reg_file[9592] <= 8'h33;
            reg_file[9593] <= 8'h56;
            reg_file[9594] <= 8'hC4;
            reg_file[9595] <= 8'h00;
            reg_file[9596] <= 8'h13;
            reg_file[9597] <= 8'h08;
            reg_file[9598] <= 8'h00;
            reg_file[9599] <= 8'h00;
            reg_file[9600] <= 8'h63;
            reg_file[9601] <= 8'h86;
            reg_file[9602] <= 8'h16;
            reg_file[9603] <= 8'h01;
            reg_file[9604] <= 8'h13;
            reg_file[9605] <= 8'h05;
            reg_file[9606] <= 8'hE5;
            reg_file[9607] <= 8'h43;
            reg_file[9608] <= 8'h33;
            reg_file[9609] <= 8'h18;
            reg_file[9610] <= 8'hA4;
            reg_file[9611] <= 8'h00;
            reg_file[9612] <= 8'hB3;
            reg_file[9613] <= 8'h67;
            reg_file[9614] <= 8'hF8;
            reg_file[9615] <= 8'h00;
            reg_file[9616] <= 8'hB3;
            reg_file[9617] <= 8'h37;
            reg_file[9618] <= 8'hF0;
            reg_file[9619] <= 8'h00;
            reg_file[9620] <= 8'hB3;
            reg_file[9621] <= 8'h67;
            reg_file[9622] <= 8'hF6;
            reg_file[9623] <= 8'h00;
            reg_file[9624] <= 8'h13;
            reg_file[9625] <= 8'h04;
            reg_file[9626] <= 8'h00;
            reg_file[9627] <= 8'h00;
            reg_file[9628] <= 8'h6F;
            reg_file[9629] <= 8'hF0;
            reg_file[9630] <= 8'h1F;
            reg_file[9631] <= 8'hF9;
            reg_file[9632] <= 8'h63;
            reg_file[9633] <= 8'h98;
            reg_file[9634] <= 8'h05;
            reg_file[9635] <= 8'h00;
            reg_file[9636] <= 8'h93;
            reg_file[9637] <= 8'h86;
            reg_file[9638] <= 8'h87;
            reg_file[9639] <= 8'h00;
            reg_file[9640] <= 8'h6F;
            reg_file[9641] <= 8'hF0;
            reg_file[9642] <= 8'h5F;
            reg_file[9643] <= 8'hFB;
            reg_file[9644] <= 8'hE3;
            reg_file[9645] <= 8'h9C;
            reg_file[9646] <= 8'h05;
            reg_file[9647] <= 8'hFE;
            reg_file[9648] <= 8'h93;
            reg_file[9649] <= 8'h16;
            reg_file[9650] <= 8'h84;
            reg_file[9651] <= 8'h00;
            reg_file[9652] <= 8'h63;
            reg_file[9653] <= 8'hDE;
            reg_file[9654] <= 8'h06;
            reg_file[9655] <= 8'h00;
            reg_file[9656] <= 8'h93;
            reg_file[9657] <= 8'hE4;
            reg_file[9658] <= 8'h14;
            reg_file[9659] <= 8'h00;
            reg_file[9660] <= 8'h13;
            reg_file[9661] <= 8'h04;
            reg_file[9662] <= 8'h00;
            reg_file[9663] <= 8'h00;
            reg_file[9664] <= 8'h93;
            reg_file[9665] <= 8'h07;
            reg_file[9666] <= 8'h00;
            reg_file[9667] <= 8'h00;
            reg_file[9668] <= 8'h63;
            reg_file[9669] <= 8'h16;
            reg_file[9670] <= 8'h07;
            reg_file[9671] <= 8'h02;
            reg_file[9672] <= 8'h13;
            reg_file[9673] <= 8'h07;
            reg_file[9674] <= 8'h10;
            reg_file[9675] <= 8'h00;
            reg_file[9676] <= 8'h6F;
            reg_file[9677] <= 8'hF0;
            reg_file[9678] <= 8'h5F;
            reg_file[9679] <= 8'hB8;
            reg_file[9680] <= 8'h93;
            reg_file[9681] <= 8'hD6;
            reg_file[9682] <= 8'h37;
            reg_file[9683] <= 8'h00;
            reg_file[9684] <= 8'h93;
            reg_file[9685] <= 8'h17;
            reg_file[9686] <= 8'hD4;
            reg_file[9687] <= 8'h01;
            reg_file[9688] <= 8'hB3;
            reg_file[9689] <= 8'hE7;
            reg_file[9690] <= 8'hD7;
            reg_file[9691] <= 8'h00;
            reg_file[9692] <= 8'h13;
            reg_file[9693] <= 8'h54;
            reg_file[9694] <= 8'h34;
            reg_file[9695] <= 8'h00;
            reg_file[9696] <= 8'hE3;
            reg_file[9697] <= 8'h08;
            reg_file[9698] <= 8'h07;
            reg_file[9699] <= 8'hB6;
            reg_file[9700] <= 8'h13;
            reg_file[9701] <= 8'hF7;
            reg_file[9702] <= 8'h14;
            reg_file[9703] <= 8'h00;
            reg_file[9704] <= 8'hE3;
            reg_file[9705] <= 8'h04;
            reg_file[9706] <= 8'h07;
            reg_file[9707] <= 8'hB6;
            reg_file[9708] <= 8'h13;
            reg_file[9709] <= 8'h07;
            reg_file[9710] <= 8'h00;
            reg_file[9711] <= 8'h00;
            reg_file[9712] <= 8'h93;
            reg_file[9713] <= 8'hE4;
            reg_file[9714] <= 8'h24;
            reg_file[9715] <= 8'h00;
            reg_file[9716] <= 8'h6F;
            reg_file[9717] <= 8'hF0;
            reg_file[9718] <= 8'hDF;
            reg_file[9719] <= 8'hB5;
            reg_file[9720] <= 8'hB3;
            reg_file[9721] <= 8'hE7;
            reg_file[9722] <= 8'h87;
            reg_file[9723] <= 8'h00;
            reg_file[9724] <= 8'h63;
            reg_file[9725] <= 8'h84;
            reg_file[9726] <= 8'h07;
            reg_file[9727] <= 8'h02;
            reg_file[9728] <= 8'h93;
            reg_file[9729] <= 8'h07;
            reg_file[9730] <= 8'h20;
            reg_file[9731] <= 8'h00;
            reg_file[9732] <= 8'h93;
            reg_file[9733] <= 8'hE4;
            reg_file[9734] <= 8'h14;
            reg_file[9735] <= 8'h00;
            reg_file[9736] <= 8'h63;
            reg_file[9737] <= 8'h0E;
            reg_file[9738] <= 8'hF9;
            reg_file[9739] <= 8'h02;
            reg_file[9740] <= 8'h93;
            reg_file[9741] <= 8'h07;
            reg_file[9742] <= 8'h30;
            reg_file[9743] <= 8'h00;
            reg_file[9744] <= 8'h63;
            reg_file[9745] <= 8'h02;
            reg_file[9746] <= 8'hF9;
            reg_file[9747] <= 8'h02;
            reg_file[9748] <= 8'h93;
            reg_file[9749] <= 8'h07;
            reg_file[9750] <= 8'h10;
            reg_file[9751] <= 8'h00;
            reg_file[9752] <= 8'h63;
            reg_file[9753] <= 8'h14;
            reg_file[9754] <= 8'h09;
            reg_file[9755] <= 8'h00;
            reg_file[9756] <= 8'h93;
            reg_file[9757] <= 8'h07;
            reg_file[9758] <= 8'h50;
            reg_file[9759] <= 8'h00;
            reg_file[9760] <= 8'h93;
            reg_file[9761] <= 8'hD7;
            reg_file[9762] <= 8'h37;
            reg_file[9763] <= 8'h00;
            reg_file[9764] <= 8'h93;
            reg_file[9765] <= 8'hE4;
            reg_file[9766] <= 8'h24;
            reg_file[9767] <= 8'h00;
            reg_file[9768] <= 8'h13;
            reg_file[9769] <= 8'h04;
            reg_file[9770] <= 8'h00;
            reg_file[9771] <= 8'h00;
            reg_file[9772] <= 8'h13;
            reg_file[9773] <= 8'h07;
            reg_file[9774] <= 8'h00;
            reg_file[9775] <= 8'h00;
            reg_file[9776] <= 8'h6F;
            reg_file[9777] <= 8'hF0;
            reg_file[9778] <= 8'h1F;
            reg_file[9779] <= 8'hB2;
            reg_file[9780] <= 8'h93;
            reg_file[9781] <= 8'h07;
            reg_file[9782] <= 8'h90;
            reg_file[9783] <= 8'h00;
            reg_file[9784] <= 8'hE3;
            reg_file[9785] <= 8'h84;
            reg_file[9786] <= 8'h05;
            reg_file[9787] <= 8'hFE;
            reg_file[9788] <= 8'h93;
            reg_file[9789] <= 8'h07;
            reg_file[9790] <= 8'h10;
            reg_file[9791] <= 8'h00;
            reg_file[9792] <= 8'h6F;
            reg_file[9793] <= 8'hF0;
            reg_file[9794] <= 8'h1F;
            reg_file[9795] <= 8'hFE;
            reg_file[9796] <= 8'h93;
            reg_file[9797] <= 8'h07;
            reg_file[9798] <= 8'h90;
            reg_file[9799] <= 8'h00;
            reg_file[9800] <= 8'hE3;
            reg_file[9801] <= 8'h9C;
            reg_file[9802] <= 8'h05;
            reg_file[9803] <= 8'hFC;
            reg_file[9804] <= 8'h6F;
            reg_file[9805] <= 8'hF0;
            reg_file[9806] <= 8'h1F;
            reg_file[9807] <= 8'hFF;
            reg_file[9808] <= 8'h13;
            reg_file[9809] <= 8'h04;
            reg_file[9810] <= 8'h00;
            reg_file[9811] <= 8'h00;
            reg_file[9812] <= 8'h93;
            reg_file[9813] <= 8'h07;
            reg_file[9814] <= 8'h00;
            reg_file[9815] <= 8'h00;
            reg_file[9816] <= 8'h13;
            reg_file[9817] <= 8'h07;
            reg_file[9818] <= 8'hF0;
            reg_file[9819] <= 8'h7F;
            reg_file[9820] <= 8'h6F;
            reg_file[9821] <= 8'hF0;
            reg_file[9822] <= 8'h5F;
            reg_file[9823] <= 8'hAF;
            reg_file[9824] <= 8'h37;
            reg_file[9825] <= 8'h04;
            reg_file[9826] <= 8'h08;
            reg_file[9827] <= 8'h00;
            reg_file[9828] <= 8'h93;
            reg_file[9829] <= 8'h07;
            reg_file[9830] <= 8'h00;
            reg_file[9831] <= 8'h00;
            reg_file[9832] <= 8'h13;
            reg_file[9833] <= 8'h07;
            reg_file[9834] <= 8'hF0;
            reg_file[9835] <= 8'h7F;
            reg_file[9836] <= 8'h93;
            reg_file[9837] <= 8'h05;
            reg_file[9838] <= 8'h00;
            reg_file[9839] <= 8'h00;
            reg_file[9840] <= 8'h6F;
            reg_file[9841] <= 8'hF0;
            reg_file[9842] <= 8'h1F;
            reg_file[9843] <= 8'hAE;
            reg_file[9844] <= 8'h13;
            reg_file[9845] <= 8'h01;
            reg_file[9846] <= 8'h01;
            reg_file[9847] <= 8'hFE;
            reg_file[9848] <= 8'h23;
            reg_file[9849] <= 8'h2E;
            reg_file[9850] <= 8'h11;
            reg_file[9851] <= 8'h00;
            reg_file[9852] <= 8'h23;
            reg_file[9853] <= 8'h2C;
            reg_file[9854] <= 8'h81;
            reg_file[9855] <= 8'h00;
            reg_file[9856] <= 8'h23;
            reg_file[9857] <= 8'h2A;
            reg_file[9858] <= 8'h91;
            reg_file[9859] <= 8'h00;
            reg_file[9860] <= 8'h23;
            reg_file[9861] <= 8'h28;
            reg_file[9862] <= 8'h21;
            reg_file[9863] <= 8'h01;
            reg_file[9864] <= 8'h23;
            reg_file[9865] <= 8'h26;
            reg_file[9866] <= 8'h31;
            reg_file[9867] <= 8'h01;
            reg_file[9868] <= 8'h23;
            reg_file[9869] <= 8'h24;
            reg_file[9870] <= 8'h41;
            reg_file[9871] <= 8'h01;
            reg_file[9872] <= 8'hF3;
            reg_file[9873] <= 8'h29;
            reg_file[9874] <= 8'h20;
            reg_file[9875] <= 8'h00;
            reg_file[9876] <= 8'hB7;
            reg_file[9877] <= 8'h08;
            reg_file[9878] <= 8'h10;
            reg_file[9879] <= 8'h00;
            reg_file[9880] <= 8'h93;
            reg_file[9881] <= 8'h88;
            reg_file[9882] <= 8'hF8;
            reg_file[9883] <= 8'hFF;
            reg_file[9884] <= 8'hB3;
            reg_file[9885] <= 8'hF7;
            reg_file[9886] <= 8'hB8;
            reg_file[9887] <= 8'h00;
            reg_file[9888] <= 8'h13;
            reg_file[9889] <= 8'h57;
            reg_file[9890] <= 8'hD5;
            reg_file[9891] <= 8'h01;
            reg_file[9892] <= 8'h13;
            reg_file[9893] <= 8'hD4;
            reg_file[9894] <= 8'h45;
            reg_file[9895] <= 8'h01;
            reg_file[9896] <= 8'h93;
            reg_file[9897] <= 8'hD4;
            reg_file[9898] <= 8'hF5;
            reg_file[9899] <= 8'h01;
            reg_file[9900] <= 8'h93;
            reg_file[9901] <= 8'h97;
            reg_file[9902] <= 8'h37;
            reg_file[9903] <= 8'h00;
            reg_file[9904] <= 8'hB3;
            reg_file[9905] <= 8'hF5;
            reg_file[9906] <= 8'hD8;
            reg_file[9907] <= 8'h00;
            reg_file[9908] <= 8'h93;
            reg_file[9909] <= 8'h95;
            reg_file[9910] <= 8'h35;
            reg_file[9911] <= 8'h00;
            reg_file[9912] <= 8'h93;
            reg_file[9913] <= 8'hD8;
            reg_file[9914] <= 8'h46;
            reg_file[9915] <= 8'h01;
            reg_file[9916] <= 8'hB3;
            reg_file[9917] <= 8'h67;
            reg_file[9918] <= 8'hF7;
            reg_file[9919] <= 8'h00;
            reg_file[9920] <= 8'h13;
            reg_file[9921] <= 8'h57;
            reg_file[9922] <= 8'hD6;
            reg_file[9923] <= 8'h01;
            reg_file[9924] <= 8'h33;
            reg_file[9925] <= 8'h67;
            reg_file[9926] <= 8'hB7;
            reg_file[9927] <= 8'h00;
            reg_file[9928] <= 8'h93;
            reg_file[9929] <= 8'hF8;
            reg_file[9930] <= 8'hF8;
            reg_file[9931] <= 8'h7F;
            reg_file[9932] <= 8'h93;
            reg_file[9933] <= 8'h05;
            reg_file[9934] <= 8'hF0;
            reg_file[9935] <= 8'h7F;
            reg_file[9936] <= 8'h13;
            reg_file[9937] <= 8'h74;
            reg_file[9938] <= 8'hF4;
            reg_file[9939] <= 8'h7F;
            reg_file[9940] <= 8'h13;
            reg_file[9941] <= 8'h15;
            reg_file[9942] <= 8'h35;
            reg_file[9943] <= 8'h00;
            reg_file[9944] <= 8'h93;
            reg_file[9945] <= 8'hD6;
            reg_file[9946] <= 8'hF6;
            reg_file[9947] <= 8'h01;
            reg_file[9948] <= 8'h13;
            reg_file[9949] <= 8'h16;
            reg_file[9950] <= 8'h36;
            reg_file[9951] <= 8'h00;
            reg_file[9952] <= 8'h63;
            reg_file[9953] <= 8'h96;
            reg_file[9954] <= 8'hB8;
            reg_file[9955] <= 8'h00;
            reg_file[9956] <= 8'hB3;
            reg_file[9957] <= 8'h65;
            reg_file[9958] <= 8'hC7;
            reg_file[9959] <= 8'h00;
            reg_file[9960] <= 8'h63;
            reg_file[9961] <= 8'h94;
            reg_file[9962] <= 8'h05;
            reg_file[9963] <= 8'h00;
            reg_file[9964] <= 8'h93;
            reg_file[9965] <= 8'hC6;
            reg_file[9966] <= 8'h16;
            reg_file[9967] <= 8'h00;
            reg_file[9968] <= 8'h33;
            reg_file[9969] <= 8'h08;
            reg_file[9970] <= 8'h14;
            reg_file[9971] <= 8'h41;
            reg_file[9972] <= 8'h63;
            reg_file[9973] <= 8'h9E;
            reg_file[9974] <= 8'h96;
            reg_file[9975] <= 8'h4E;
            reg_file[9976] <= 8'h63;
            reg_file[9977] <= 8'h54;
            reg_file[9978] <= 8'h00;
            reg_file[9979] <= 8'h17;
            reg_file[9980] <= 8'h63;
            reg_file[9981] <= 8'h9A;
            reg_file[9982] <= 8'h08;
            reg_file[9983] <= 8'h06;
            reg_file[9984] <= 8'hB3;
            reg_file[9985] <= 8'h66;
            reg_file[9986] <= 8'hC7;
            reg_file[9987] <= 8'h00;
            reg_file[9988] <= 8'h63;
            reg_file[9989] <= 8'h96;
            reg_file[9990] <= 8'h06;
            reg_file[9991] <= 8'h02;
            reg_file[9992] <= 8'h13;
            reg_file[9993] <= 8'h07;
            reg_file[9994] <= 8'hF0;
            reg_file[9995] <= 8'h7F;
            reg_file[9996] <= 8'h13;
            reg_file[9997] <= 8'h04;
            reg_file[9998] <= 8'h00;
            reg_file[9999] <= 8'h00;
            reg_file[10000] <= 8'h63;
            reg_file[10001] <= 8'h1E;
            reg_file[10002] <= 8'hE8;
            reg_file[10003] <= 8'h2C;
            reg_file[10004] <= 8'h33;
            reg_file[10005] <= 8'hE7;
            reg_file[10006] <= 8'hA7;
            reg_file[10007] <= 8'h00;
            reg_file[10008] <= 8'hE3;
            reg_file[10009] <= 8'h00;
            reg_file[10010] <= 8'h07;
            reg_file[10011] <= 8'h1E;
            reg_file[10012] <= 8'h37;
            reg_file[10013] <= 8'h04;
            reg_file[10014] <= 8'h40;
            reg_file[10015] <= 8'h00;
            reg_file[10016] <= 8'h33;
            reg_file[10017] <= 8'hF4;
            reg_file[10018] <= 8'h87;
            reg_file[10019] <= 8'h00;
            reg_file[10020] <= 8'h13;
            reg_file[10021] <= 8'h34;
            reg_file[10022] <= 8'h14;
            reg_file[10023] <= 8'h00;
            reg_file[10024] <= 8'h13;
            reg_file[10025] <= 8'h14;
            reg_file[10026] <= 8'h44;
            reg_file[10027] <= 8'h00;
            reg_file[10028] <= 8'h6F;
            reg_file[10029] <= 8'h00;
            reg_file[10030] <= 8'h00;
            reg_file[10031] <= 8'h2C;
            reg_file[10032] <= 8'h93;
            reg_file[10033] <= 8'h06;
            reg_file[10034] <= 8'hF8;
            reg_file[10035] <= 8'hFF;
            reg_file[10036] <= 8'h63;
            reg_file[10037] <= 8'h9E;
            reg_file[10038] <= 8'h06;
            reg_file[10039] <= 8'h00;
            reg_file[10040] <= 8'h33;
            reg_file[10041] <= 8'h06;
            reg_file[10042] <= 8'hA6;
            reg_file[10043] <= 8'h00;
            reg_file[10044] <= 8'hB3;
            reg_file[10045] <= 8'h87;
            reg_file[10046] <= 8'hE7;
            reg_file[10047] <= 8'h00;
            reg_file[10048] <= 8'hB3;
            reg_file[10049] <= 8'h36;
            reg_file[10050] <= 8'hA6;
            reg_file[10051] <= 8'h00;
            reg_file[10052] <= 8'h33;
            reg_file[10053] <= 8'h87;
            reg_file[10054] <= 8'hD7;
            reg_file[10055] <= 8'h00;
            reg_file[10056] <= 8'h13;
            reg_file[10057] <= 8'h08;
            reg_file[10058] <= 8'h10;
            reg_file[10059] <= 8'h00;
            reg_file[10060] <= 8'h6F;
            reg_file[10061] <= 8'h00;
            reg_file[10062] <= 8'h00;
            reg_file[10063] <= 8'h0A;
            reg_file[10064] <= 8'h93;
            reg_file[10065] <= 8'h05;
            reg_file[10066] <= 8'hF0;
            reg_file[10067] <= 8'h7F;
            reg_file[10068] <= 8'h63;
            reg_file[10069] <= 8'h18;
            reg_file[10070] <= 8'hB8;
            reg_file[10071] <= 8'h04;
            reg_file[10072] <= 8'h33;
            reg_file[10073] <= 8'hE7;
            reg_file[10074] <= 8'hA7;
            reg_file[10075] <= 8'h00;
            reg_file[10076] <= 8'hE3;
            reg_file[10077] <= 8'h10;
            reg_file[10078] <= 8'h07;
            reg_file[10079] <= 8'hFC;
            reg_file[10080] <= 8'h93;
            reg_file[10081] <= 8'h07;
            reg_file[10082] <= 8'h00;
            reg_file[10083] <= 8'h00;
            reg_file[10084] <= 8'h13;
            reg_file[10085] <= 8'h05;
            reg_file[10086] <= 8'h00;
            reg_file[10087] <= 8'h00;
            reg_file[10088] <= 8'h13;
            reg_file[10089] <= 8'h04;
            reg_file[10090] <= 8'h00;
            reg_file[10091] <= 8'h00;
            reg_file[10092] <= 8'h6F;
            reg_file[10093] <= 8'h00;
            reg_file[10094] <= 8'h40;
            reg_file[10095] <= 8'h31;
            reg_file[10096] <= 8'h93;
            reg_file[10097] <= 8'h06;
            reg_file[10098] <= 8'hF0;
            reg_file[10099] <= 8'h7F;
            reg_file[10100] <= 8'h63;
            reg_file[10101] <= 8'h12;
            reg_file[10102] <= 8'hD4;
            reg_file[10103] <= 8'h02;
            reg_file[10104] <= 8'h33;
            reg_file[10105] <= 8'hE7;
            reg_file[10106] <= 8'hA7;
            reg_file[10107] <= 8'h00;
            reg_file[10108] <= 8'hE3;
            reg_file[10109] <= 8'h04;
            reg_file[10110] <= 8'h07;
            reg_file[10111] <= 8'h18;
            reg_file[10112] <= 8'h13;
            reg_file[10113] <= 8'h97;
            reg_file[10114] <= 8'h97;
            reg_file[10115] <= 8'h00;
            reg_file[10116] <= 8'h13;
            reg_file[10117] <= 8'h08;
            reg_file[10118] <= 8'hF0;
            reg_file[10119] <= 8'h7F;
            reg_file[10120] <= 8'h93;
            reg_file[10121] <= 8'h08;
            reg_file[10122] <= 8'h00;
            reg_file[10123] <= 8'h00;
            reg_file[10124] <= 8'h63;
            reg_file[10125] <= 8'h4E;
            reg_file[10126] <= 8'h07;
            reg_file[10127] <= 8'h3A;
            reg_file[10128] <= 8'h13;
            reg_file[10129] <= 8'h04;
            reg_file[10130] <= 8'h00;
            reg_file[10131] <= 8'h01;
            reg_file[10132] <= 8'h6F;
            reg_file[10133] <= 8'h00;
            reg_file[10134] <= 8'h80;
            reg_file[10135] <= 8'h25;
            reg_file[10136] <= 8'hB7;
            reg_file[10137] <= 8'h06;
            reg_file[10138] <= 8'h80;
            reg_file[10139] <= 8'h00;
            reg_file[10140] <= 8'h33;
            reg_file[10141] <= 8'h67;
            reg_file[10142] <= 8'hD7;
            reg_file[10143] <= 8'h00;
            reg_file[10144] <= 8'h93;
            reg_file[10145] <= 8'h06;
            reg_file[10146] <= 8'h08;
            reg_file[10147] <= 8'h00;
            reg_file[10148] <= 8'h93;
            reg_file[10149] <= 8'h05;
            reg_file[10150] <= 8'h80;
            reg_file[10151] <= 8'h03;
            reg_file[10152] <= 8'h63;
            reg_file[10153] <= 8'hC6;
            reg_file[10154] <= 8'hD5;
            reg_file[10155] <= 8'h0A;
            reg_file[10156] <= 8'h93;
            reg_file[10157] <= 8'h05;
            reg_file[10158] <= 8'hF0;
            reg_file[10159] <= 8'h01;
            reg_file[10160] <= 8'h63;
            reg_file[10161] <= 8'hC8;
            reg_file[10162] <= 8'hD5;
            reg_file[10163] <= 8'h06;
            reg_file[10164] <= 8'h13;
            reg_file[10165] <= 8'h08;
            reg_file[10166] <= 8'h00;
            reg_file[10167] <= 8'h02;
            reg_file[10168] <= 8'h33;
            reg_file[10169] <= 8'h08;
            reg_file[10170] <= 8'hD8;
            reg_file[10171] <= 8'h40;
            reg_file[10172] <= 8'hB3;
            reg_file[10173] <= 8'h58;
            reg_file[10174] <= 8'hD6;
            reg_file[10175] <= 8'h00;
            reg_file[10176] <= 8'hB3;
            reg_file[10177] <= 8'h15;
            reg_file[10178] <= 8'h07;
            reg_file[10179] <= 8'h01;
            reg_file[10180] <= 8'h33;
            reg_file[10181] <= 8'h16;
            reg_file[10182] <= 8'h06;
            reg_file[10183] <= 8'h01;
            reg_file[10184] <= 8'hB3;
            reg_file[10185] <= 8'hE5;
            reg_file[10186] <= 8'h15;
            reg_file[10187] <= 8'h01;
            reg_file[10188] <= 8'h33;
            reg_file[10189] <= 8'h36;
            reg_file[10190] <= 8'hC0;
            reg_file[10191] <= 8'h00;
            reg_file[10192] <= 8'h33;
            reg_file[10193] <= 8'hE6;
            reg_file[10194] <= 8'hC5;
            reg_file[10195] <= 8'h00;
            reg_file[10196] <= 8'hB3;
            reg_file[10197] <= 8'h56;
            reg_file[10198] <= 8'hD7;
            reg_file[10199] <= 8'h00;
            reg_file[10200] <= 8'h33;
            reg_file[10201] <= 8'h06;
            reg_file[10202] <= 8'hA6;
            reg_file[10203] <= 8'h00;
            reg_file[10204] <= 8'hB3;
            reg_file[10205] <= 8'h86;
            reg_file[10206] <= 8'hF6;
            reg_file[10207] <= 8'h00;
            reg_file[10208] <= 8'hB3;
            reg_file[10209] <= 8'h37;
            reg_file[10210] <= 8'hA6;
            reg_file[10211] <= 8'h00;
            reg_file[10212] <= 8'h33;
            reg_file[10213] <= 8'h87;
            reg_file[10214] <= 8'hF6;
            reg_file[10215] <= 8'h00;
            reg_file[10216] <= 8'h13;
            reg_file[10217] <= 8'h08;
            reg_file[10218] <= 8'h04;
            reg_file[10219] <= 8'h00;
            reg_file[10220] <= 8'h93;
            reg_file[10221] <= 8'h17;
            reg_file[10222] <= 8'h87;
            reg_file[10223] <= 8'h00;
            reg_file[10224] <= 8'h63;
            reg_file[10225] <= 8'hD6;
            reg_file[10226] <= 8'h07;
            reg_file[10227] <= 8'h08;
            reg_file[10228] <= 8'h13;
            reg_file[10229] <= 8'h08;
            reg_file[10230] <= 8'h18;
            reg_file[10231] <= 8'h00;
            reg_file[10232] <= 8'h93;
            reg_file[10233] <= 8'h07;
            reg_file[10234] <= 8'hF0;
            reg_file[10235] <= 8'h7F;
            reg_file[10236] <= 8'h63;
            reg_file[10237] <= 8'h02;
            reg_file[10238] <= 8'hF8;
            reg_file[10239] <= 8'h3C;
            reg_file[10240] <= 8'hB7;
            reg_file[10241] <= 8'h07;
            reg_file[10242] <= 8'h80;
            reg_file[10243] <= 8'hFF;
            reg_file[10244] <= 8'h93;
            reg_file[10245] <= 8'h87;
            reg_file[10246] <= 8'hF7;
            reg_file[10247] <= 8'hFF;
            reg_file[10248] <= 8'h13;
            reg_file[10249] <= 8'h55;
            reg_file[10250] <= 8'h16;
            reg_file[10251] <= 8'h00;
            reg_file[10252] <= 8'hB3;
            reg_file[10253] <= 8'h77;
            reg_file[10254] <= 8'hF7;
            reg_file[10255] <= 8'h00;
            reg_file[10256] <= 8'h13;
            reg_file[10257] <= 8'h76;
            reg_file[10258] <= 8'h16;
            reg_file[10259] <= 8'h00;
            reg_file[10260] <= 8'h33;
            reg_file[10261] <= 8'h66;
            reg_file[10262] <= 8'hC5;
            reg_file[10263] <= 8'h00;
            reg_file[10264] <= 8'h13;
            reg_file[10265] <= 8'h95;
            reg_file[10266] <= 8'hF7;
            reg_file[10267] <= 8'h01;
            reg_file[10268] <= 8'h6F;
            reg_file[10269] <= 8'h00;
            reg_file[10270] <= 8'h00;
            reg_file[10271] <= 8'h32;
            reg_file[10272] <= 8'h93;
            reg_file[10273] <= 8'h85;
            reg_file[10274] <= 8'h06;
            reg_file[10275] <= 8'hFE;
            reg_file[10276] <= 8'h93;
            reg_file[10277] <= 8'h08;
            reg_file[10278] <= 8'h00;
            reg_file[10279] <= 8'h02;
            reg_file[10280] <= 8'hB3;
            reg_file[10281] <= 8'h55;
            reg_file[10282] <= 8'hB7;
            reg_file[10283] <= 8'h00;
            reg_file[10284] <= 8'h13;
            reg_file[10285] <= 8'h08;
            reg_file[10286] <= 8'h00;
            reg_file[10287] <= 8'h00;
            reg_file[10288] <= 8'h63;
            reg_file[10289] <= 8'h88;
            reg_file[10290] <= 8'h16;
            reg_file[10291] <= 8'h01;
            reg_file[10292] <= 8'h13;
            reg_file[10293] <= 8'h08;
            reg_file[10294] <= 8'h00;
            reg_file[10295] <= 8'h04;
            reg_file[10296] <= 8'hB3;
            reg_file[10297] <= 8'h06;
            reg_file[10298] <= 8'hD8;
            reg_file[10299] <= 8'h40;
            reg_file[10300] <= 8'h33;
            reg_file[10301] <= 8'h18;
            reg_file[10302] <= 8'hD7;
            reg_file[10303] <= 8'h00;
            reg_file[10304] <= 8'h33;
            reg_file[10305] <= 8'h66;
            reg_file[10306] <= 8'hC8;
            reg_file[10307] <= 8'h00;
            reg_file[10308] <= 8'h33;
            reg_file[10309] <= 8'h36;
            reg_file[10310] <= 8'hC0;
            reg_file[10311] <= 8'h00;
            reg_file[10312] <= 8'h33;
            reg_file[10313] <= 8'hE6;
            reg_file[10314] <= 8'hC5;
            reg_file[10315] <= 8'h00;
            reg_file[10316] <= 8'h93;
            reg_file[10317] <= 8'h06;
            reg_file[10318] <= 8'h00;
            reg_file[10319] <= 8'h00;
            reg_file[10320] <= 8'h6F;
            reg_file[10321] <= 8'hF0;
            reg_file[10322] <= 8'h9F;
            reg_file[10323] <= 8'hF8;
            reg_file[10324] <= 8'h33;
            reg_file[10325] <= 8'h66;
            reg_file[10326] <= 8'hC7;
            reg_file[10327] <= 8'h00;
            reg_file[10328] <= 8'h33;
            reg_file[10329] <= 8'h36;
            reg_file[10330] <= 8'hC0;
            reg_file[10331] <= 8'h00;
            reg_file[10332] <= 8'h6F;
            reg_file[10333] <= 8'hF0;
            reg_file[10334] <= 8'h1F;
            reg_file[10335] <= 8'hFF;
            reg_file[10336] <= 8'h63;
            reg_file[10337] <= 8'h0E;
            reg_file[10338] <= 8'h08;
            reg_file[10339] <= 8'h12;
            reg_file[10340] <= 8'h33;
            reg_file[10341] <= 8'h88;
            reg_file[10342] <= 8'h88;
            reg_file[10343] <= 8'h40;
            reg_file[10344] <= 8'h63;
            reg_file[10345] <= 8'h16;
            reg_file[10346] <= 8'h04;
            reg_file[10347] <= 8'h06;
            reg_file[10348] <= 8'hB3;
            reg_file[10349] <= 8'hE6;
            reg_file[10350] <= 8'hA7;
            reg_file[10351] <= 8'h00;
            reg_file[10352] <= 8'h63;
            reg_file[10353] <= 8'h9E;
            reg_file[10354] <= 8'h06;
            reg_file[10355] <= 8'h00;
            reg_file[10356] <= 8'h93;
            reg_file[10357] <= 8'h07;
            reg_file[10358] <= 8'hF0;
            reg_file[10359] <= 8'h7F;
            reg_file[10360] <= 8'h63;
            reg_file[10361] <= 8'h0E;
            reg_file[10362] <= 8'hF8;
            reg_file[10363] <= 8'h02;
            reg_file[10364] <= 8'h93;
            reg_file[10365] <= 8'h07;
            reg_file[10366] <= 8'h07;
            reg_file[10367] <= 8'h00;
            reg_file[10368] <= 8'h13;
            reg_file[10369] <= 8'h05;
            reg_file[10370] <= 8'h06;
            reg_file[10371] <= 8'h00;
            reg_file[10372] <= 8'h63;
            reg_file[10373] <= 8'h04;
            reg_file[10374] <= 8'h08;
            reg_file[10375] <= 8'h5C;
            reg_file[10376] <= 8'h6F;
            reg_file[10377] <= 8'h00;
            reg_file[10378] <= 8'hC0;
            reg_file[10379] <= 8'h2B;
            reg_file[10380] <= 8'h93;
            reg_file[10381] <= 8'h05;
            reg_file[10382] <= 8'hF8;
            reg_file[10383] <= 8'hFF;
            reg_file[10384] <= 8'h63;
            reg_file[10385] <= 8'h9E;
            reg_file[10386] <= 8'h05;
            reg_file[10387] <= 8'h00;
            reg_file[10388] <= 8'hB3;
            reg_file[10389] <= 8'h06;
            reg_file[10390] <= 8'hC5;
            reg_file[10391] <= 8'h00;
            reg_file[10392] <= 8'h33;
            reg_file[10393] <= 8'hB6;
            reg_file[10394] <= 8'hC6;
            reg_file[10395] <= 8'h00;
            reg_file[10396] <= 8'hB3;
            reg_file[10397] <= 8'h87;
            reg_file[10398] <= 8'hE7;
            reg_file[10399] <= 8'h00;
            reg_file[10400] <= 8'h33;
            reg_file[10401] <= 8'h87;
            reg_file[10402] <= 8'hC7;
            reg_file[10403] <= 8'h00;
            reg_file[10404] <= 8'h13;
            reg_file[10405] <= 8'h86;
            reg_file[10406] <= 8'h06;
            reg_file[10407] <= 8'h00;
            reg_file[10408] <= 8'h6F;
            reg_file[10409] <= 8'hF0;
            reg_file[10410] <= 8'h1F;
            reg_file[10411] <= 8'hEA;
            reg_file[10412] <= 8'h93;
            reg_file[10413] <= 8'h06;
            reg_file[10414] <= 8'hF0;
            reg_file[10415] <= 8'h7F;
            reg_file[10416] <= 8'h63;
            reg_file[10417] <= 8'h1E;
            reg_file[10418] <= 8'hD8;
            reg_file[10419] <= 8'h04;
            reg_file[10420] <= 8'h33;
            reg_file[10421] <= 8'h65;
            reg_file[10422] <= 8'hC7;
            reg_file[10423] <= 8'h00;
            reg_file[10424] <= 8'h93;
            reg_file[10425] <= 8'h07;
            reg_file[10426] <= 8'h00;
            reg_file[10427] <= 8'h00;
            reg_file[10428] <= 8'h63;
            reg_file[10429] <= 8'h02;
            reg_file[10430] <= 8'h05;
            reg_file[10431] <= 8'h1C;
            reg_file[10432] <= 8'h93;
            reg_file[10433] <= 8'h17;
            reg_file[10434] <= 8'h97;
            reg_file[10435] <= 8'h00;
            reg_file[10436] <= 8'hE3;
            reg_file[10437] <= 8'hC6;
            reg_file[10438] <= 8'h07;
            reg_file[10439] <= 8'h04;
            reg_file[10440] <= 8'h93;
            reg_file[10441] <= 8'h07;
            reg_file[10442] <= 8'h07;
            reg_file[10443] <= 8'h00;
            reg_file[10444] <= 8'h13;
            reg_file[10445] <= 8'h05;
            reg_file[10446] <= 8'h06;
            reg_file[10447] <= 8'h00;
            reg_file[10448] <= 8'h6F;
            reg_file[10449] <= 8'h00;
            reg_file[10450] <= 8'h80;
            reg_file[10451] <= 8'h02;
            reg_file[10452] <= 8'h93;
            reg_file[10453] <= 8'h06;
            reg_file[10454] <= 8'hF0;
            reg_file[10455] <= 8'h7F;
            reg_file[10456] <= 8'h63;
            reg_file[10457] <= 8'h94;
            reg_file[10458] <= 8'hD8;
            reg_file[10459] <= 8'h02;
            reg_file[10460] <= 8'h33;
            reg_file[10461] <= 8'h65;
            reg_file[10462] <= 8'hC7;
            reg_file[10463] <= 8'h00;
            reg_file[10464] <= 8'h63;
            reg_file[10465] <= 8'h04;
            reg_file[10466] <= 8'h05;
            reg_file[10467] <= 8'h7E;
            reg_file[10468] <= 8'h93;
            reg_file[10469] <= 8'h17;
            reg_file[10470] <= 8'h97;
            reg_file[10471] <= 8'h00;
            reg_file[10472] <= 8'h63;
            reg_file[10473] <= 8'hC6;
            reg_file[10474] <= 8'h07;
            reg_file[10475] <= 8'h7E;
            reg_file[10476] <= 8'h93;
            reg_file[10477] <= 8'h07;
            reg_file[10478] <= 8'h07;
            reg_file[10479] <= 8'h00;
            reg_file[10480] <= 8'h13;
            reg_file[10481] <= 8'h05;
            reg_file[10482] <= 8'h06;
            reg_file[10483] <= 8'h00;
            reg_file[10484] <= 8'h13;
            reg_file[10485] <= 8'h08;
            reg_file[10486] <= 8'hF0;
            reg_file[10487] <= 8'h7F;
            reg_file[10488] <= 8'h93;
            reg_file[10489] <= 8'h08;
            reg_file[10490] <= 8'h00;
            reg_file[10491] <= 8'h00;
            reg_file[10492] <= 8'h6F;
            reg_file[10493] <= 8'hF0;
            reg_file[10494] <= 8'h5F;
            reg_file[10495] <= 8'hE9;
            reg_file[10496] <= 8'hB7;
            reg_file[10497] <= 8'h06;
            reg_file[10498] <= 8'h80;
            reg_file[10499] <= 8'h00;
            reg_file[10500] <= 8'hB3;
            reg_file[10501] <= 8'hE7;
            reg_file[10502] <= 8'hD7;
            reg_file[10503] <= 8'h00;
            reg_file[10504] <= 8'h93;
            reg_file[10505] <= 8'h05;
            reg_file[10506] <= 8'h08;
            reg_file[10507] <= 8'h00;
            reg_file[10508] <= 8'h93;
            reg_file[10509] <= 8'h06;
            reg_file[10510] <= 8'h80;
            reg_file[10511] <= 8'h03;
            reg_file[10512] <= 8'h63;
            reg_file[10513] <= 8'hC0;
            reg_file[10514] <= 8'hB6;
            reg_file[10515] <= 8'h08;
            reg_file[10516] <= 8'h93;
            reg_file[10517] <= 8'h06;
            reg_file[10518] <= 8'hF0;
            reg_file[10519] <= 8'h01;
            reg_file[10520] <= 8'h63;
            reg_file[10521] <= 8'hC2;
            reg_file[10522] <= 8'hB6;
            reg_file[10523] <= 8'h04;
            reg_file[10524] <= 8'h13;
            reg_file[10525] <= 8'h08;
            reg_file[10526] <= 8'h00;
            reg_file[10527] <= 8'h02;
            reg_file[10528] <= 8'h33;
            reg_file[10529] <= 8'h08;
            reg_file[10530] <= 8'hB8;
            reg_file[10531] <= 8'h40;
            reg_file[10532] <= 8'hB3;
            reg_file[10533] <= 8'h96;
            reg_file[10534] <= 8'h07;
            reg_file[10535] <= 8'h01;
            reg_file[10536] <= 8'h33;
            reg_file[10537] <= 8'h53;
            reg_file[10538] <= 8'hB5;
            reg_file[10539] <= 8'h00;
            reg_file[10540] <= 8'h33;
            reg_file[10541] <= 8'h15;
            reg_file[10542] <= 8'h05;
            reg_file[10543] <= 8'h01;
            reg_file[10544] <= 8'hB3;
            reg_file[10545] <= 8'hE6;
            reg_file[10546] <= 8'h66;
            reg_file[10547] <= 8'h00;
            reg_file[10548] <= 8'h33;
            reg_file[10549] <= 8'h35;
            reg_file[10550] <= 8'hA0;
            reg_file[10551] <= 8'h00;
            reg_file[10552] <= 8'h33;
            reg_file[10553] <= 8'hE5;
            reg_file[10554] <= 8'hA6;
            reg_file[10555] <= 8'h00;
            reg_file[10556] <= 8'hB3;
            reg_file[10557] <= 8'hD7;
            reg_file[10558] <= 8'hB7;
            reg_file[10559] <= 8'h00;
            reg_file[10560] <= 8'hB3;
            reg_file[10561] <= 8'h06;
            reg_file[10562] <= 8'hC5;
            reg_file[10563] <= 8'h00;
            reg_file[10564] <= 8'hB3;
            reg_file[10565] <= 8'h87;
            reg_file[10566] <= 8'hE7;
            reg_file[10567] <= 8'h00;
            reg_file[10568] <= 8'h33;
            reg_file[10569] <= 8'hB7;
            reg_file[10570] <= 8'hC6;
            reg_file[10571] <= 8'h00;
            reg_file[10572] <= 8'h33;
            reg_file[10573] <= 8'h87;
            reg_file[10574] <= 8'hE7;
            reg_file[10575] <= 8'h00;
            reg_file[10576] <= 8'h13;
            reg_file[10577] <= 8'h86;
            reg_file[10578] <= 8'h06;
            reg_file[10579] <= 8'h00;
            reg_file[10580] <= 8'h13;
            reg_file[10581] <= 8'h88;
            reg_file[10582] <= 8'h08;
            reg_file[10583] <= 8'h00;
            reg_file[10584] <= 8'h6F;
            reg_file[10585] <= 8'hF0;
            reg_file[10586] <= 8'h5F;
            reg_file[10587] <= 8'hE9;
            reg_file[10588] <= 8'h93;
            reg_file[10589] <= 8'h86;
            reg_file[10590] <= 8'h05;
            reg_file[10591] <= 8'hFE;
            reg_file[10592] <= 8'h13;
            reg_file[10593] <= 8'h03;
            reg_file[10594] <= 8'h00;
            reg_file[10595] <= 8'h02;
            reg_file[10596] <= 8'hB3;
            reg_file[10597] <= 8'hD6;
            reg_file[10598] <= 8'hD7;
            reg_file[10599] <= 8'h00;
            reg_file[10600] <= 8'h13;
            reg_file[10601] <= 8'h08;
            reg_file[10602] <= 8'h00;
            reg_file[10603] <= 8'h00;
            reg_file[10604] <= 8'h63;
            reg_file[10605] <= 8'h88;
            reg_file[10606] <= 8'h65;
            reg_file[10607] <= 8'h00;
            reg_file[10608] <= 8'h13;
            reg_file[10609] <= 8'h08;
            reg_file[10610] <= 8'h00;
            reg_file[10611] <= 8'h04;
            reg_file[10612] <= 8'hB3;
            reg_file[10613] <= 8'h05;
            reg_file[10614] <= 8'hB8;
            reg_file[10615] <= 8'h40;
            reg_file[10616] <= 8'h33;
            reg_file[10617] <= 8'h98;
            reg_file[10618] <= 8'hB7;
            reg_file[10619] <= 8'h00;
            reg_file[10620] <= 8'h33;
            reg_file[10621] <= 8'h65;
            reg_file[10622] <= 8'hA8;
            reg_file[10623] <= 8'h00;
            reg_file[10624] <= 8'h33;
            reg_file[10625] <= 8'h35;
            reg_file[10626] <= 8'hA0;
            reg_file[10627] <= 8'h00;
            reg_file[10628] <= 8'h33;
            reg_file[10629] <= 8'hE5;
            reg_file[10630] <= 8'hA6;
            reg_file[10631] <= 8'h00;
            reg_file[10632] <= 8'h93;
            reg_file[10633] <= 8'h07;
            reg_file[10634] <= 8'h00;
            reg_file[10635] <= 8'h00;
            reg_file[10636] <= 8'h6F;
            reg_file[10637] <= 8'hF0;
            reg_file[10638] <= 8'h5F;
            reg_file[10639] <= 8'hFB;
            reg_file[10640] <= 8'h33;
            reg_file[10641] <= 8'hE5;
            reg_file[10642] <= 8'hA7;
            reg_file[10643] <= 8'h00;
            reg_file[10644] <= 8'h33;
            reg_file[10645] <= 8'h35;
            reg_file[10646] <= 8'hA0;
            reg_file[10647] <= 8'h00;
            reg_file[10648] <= 8'h6F;
            reg_file[10649] <= 8'hF0;
            reg_file[10650] <= 8'h1F;
            reg_file[10651] <= 8'hFF;
            reg_file[10652] <= 8'h13;
            reg_file[10653] <= 8'h08;
            reg_file[10654] <= 8'h14;
            reg_file[10655] <= 8'h00;
            reg_file[10656] <= 8'h93;
            reg_file[10657] <= 8'h76;
            reg_file[10658] <= 8'hE8;
            reg_file[10659] <= 8'h7F;
            reg_file[10660] <= 8'h63;
            reg_file[10661] <= 8'h9C;
            reg_file[10662] <= 8'h06;
            reg_file[10663] <= 8'h16;
            reg_file[10664] <= 8'hB3;
            reg_file[10665] <= 8'hE6;
            reg_file[10666] <= 8'hA7;
            reg_file[10667] <= 8'h00;
            reg_file[10668] <= 8'h63;
            reg_file[10669] <= 8'h1E;
            reg_file[10670] <= 8'h04;
            reg_file[10671] <= 8'h04;
            reg_file[10672] <= 8'h63;
            reg_file[10673] <= 8'h8E;
            reg_file[10674] <= 8'h06;
            reg_file[10675] <= 8'h6A;
            reg_file[10676] <= 8'hB3;
            reg_file[10677] <= 8'h66;
            reg_file[10678] <= 8'hC7;
            reg_file[10679] <= 8'h00;
            reg_file[10680] <= 8'h63;
            reg_file[10681] <= 8'h8A;
            reg_file[10682] <= 8'h06;
            reg_file[10683] <= 8'h48;
            reg_file[10684] <= 8'h33;
            reg_file[10685] <= 8'h06;
            reg_file[10686] <= 8'hC5;
            reg_file[10687] <= 8'h00;
            reg_file[10688] <= 8'hB3;
            reg_file[10689] <= 8'h87;
            reg_file[10690] <= 8'hE7;
            reg_file[10691] <= 8'h00;
            reg_file[10692] <= 8'h33;
            reg_file[10693] <= 8'h35;
            reg_file[10694] <= 8'hA6;
            reg_file[10695] <= 8'h00;
            reg_file[10696] <= 8'hB3;
            reg_file[10697] <= 8'h87;
            reg_file[10698] <= 8'hA7;
            reg_file[10699] <= 8'h00;
            reg_file[10700] <= 8'h13;
            reg_file[10701] <= 8'h97;
            reg_file[10702] <= 8'h87;
            reg_file[10703] <= 8'h00;
            reg_file[10704] <= 8'h63;
            reg_file[10705] <= 8'h50;
            reg_file[10706] <= 8'h07;
            reg_file[10707] <= 8'h6A;
            reg_file[10708] <= 8'h37;
            reg_file[10709] <= 8'h07;
            reg_file[10710] <= 8'h80;
            reg_file[10711] <= 8'hFF;
            reg_file[10712] <= 8'h13;
            reg_file[10713] <= 8'h07;
            reg_file[10714] <= 8'hF7;
            reg_file[10715] <= 8'hFF;
            reg_file[10716] <= 8'hB3;
            reg_file[10717] <= 8'hF7;
            reg_file[10718] <= 8'hE7;
            reg_file[10719] <= 8'h00;
            reg_file[10720] <= 8'h13;
            reg_file[10721] <= 8'h05;
            reg_file[10722] <= 8'h06;
            reg_file[10723] <= 8'h00;
            reg_file[10724] <= 8'h93;
            reg_file[10725] <= 8'h08;
            reg_file[10726] <= 8'h00;
            reg_file[10727] <= 8'h00;
            reg_file[10728] <= 8'h13;
            reg_file[10729] <= 8'h08;
            reg_file[10730] <= 8'h10;
            reg_file[10731] <= 8'h00;
            reg_file[10732] <= 8'h13;
            reg_file[10733] <= 8'h77;
            reg_file[10734] <= 8'h75;
            reg_file[10735] <= 8'h00;
            reg_file[10736] <= 8'h63;
            reg_file[10737] <= 8'h1C;
            reg_file[10738] <= 8'h07;
            reg_file[10739] <= 8'h18;
            reg_file[10740] <= 8'h63;
            reg_file[10741] <= 8'h86;
            reg_file[10742] <= 8'h08;
            reg_file[10743] <= 8'h08;
            reg_file[10744] <= 8'h13;
            reg_file[10745] <= 8'h77;
            reg_file[10746] <= 8'h14;
            reg_file[10747] <= 8'h00;
            reg_file[10748] <= 8'h63;
            reg_file[10749] <= 8'h02;
            reg_file[10750] <= 8'h07;
            reg_file[10751] <= 8'h08;
            reg_file[10752] <= 8'h13;
            reg_file[10753] <= 8'h64;
            reg_file[10754] <= 8'h24;
            reg_file[10755] <= 8'h00;
            reg_file[10756] <= 8'h6F;
            reg_file[10757] <= 8'h00;
            reg_file[10758] <= 8'hC0;
            reg_file[10759] <= 8'h07;
            reg_file[10760] <= 8'h93;
            reg_file[10761] <= 8'h05;
            reg_file[10762] <= 8'hF0;
            reg_file[10763] <= 8'h7F;
            reg_file[10764] <= 8'h63;
            reg_file[10765] <= 8'h1A;
            reg_file[10766] <= 8'hB4;
            reg_file[10767] <= 8'h02;
            reg_file[10768] <= 8'h63;
            reg_file[10769] <= 8'h8A;
            reg_file[10770] <= 8'h06;
            reg_file[10771] <= 8'h7C;
            reg_file[10772] <= 8'h37;
            reg_file[10773] <= 8'h04;
            reg_file[10774] <= 8'h40;
            reg_file[10775] <= 8'h00;
            reg_file[10776] <= 8'h33;
            reg_file[10777] <= 8'hF4;
            reg_file[10778] <= 8'h87;
            reg_file[10779] <= 8'h00;
            reg_file[10780] <= 8'h13;
            reg_file[10781] <= 8'h34;
            reg_file[10782] <= 8'h14;
            reg_file[10783] <= 8'h00;
            reg_file[10784] <= 8'h13;
            reg_file[10785] <= 8'h14;
            reg_file[10786] <= 8'h44;
            reg_file[10787] <= 8'h00;
            reg_file[10788] <= 8'h63;
            reg_file[10789] <= 8'h92;
            reg_file[10790] <= 8'hB8;
            reg_file[10791] <= 8'h04;
            reg_file[10792] <= 8'hB3;
            reg_file[10793] <= 8'h65;
            reg_file[10794] <= 8'hC7;
            reg_file[10795] <= 8'h00;
            reg_file[10796] <= 8'h63;
            reg_file[10797] <= 8'h8E;
            reg_file[10798] <= 8'h05;
            reg_file[10799] <= 8'h00;
            reg_file[10800] <= 8'h93;
            reg_file[10801] <= 8'h15;
            reg_file[10802] <= 8'h97;
            reg_file[10803] <= 8'h00;
            reg_file[10804] <= 8'h63;
            reg_file[10805] <= 8'hCA;
            reg_file[10806] <= 8'h05;
            reg_file[10807] <= 8'h00;
            reg_file[10808] <= 8'h13;
            reg_file[10809] <= 8'h04;
            reg_file[10810] <= 8'h00;
            reg_file[10811] <= 8'h01;
            reg_file[10812] <= 8'h6F;
            reg_file[10813] <= 8'h00;
            reg_file[10814] <= 8'hC0;
            reg_file[10815] <= 8'h00;
            reg_file[10816] <= 8'h13;
            reg_file[10817] <= 8'h04;
            reg_file[10818] <= 8'h00;
            reg_file[10819] <= 8'h00;
            reg_file[10820] <= 8'hE3;
            reg_file[10821] <= 8'h82;
            reg_file[10822] <= 8'hB8;
            reg_file[10823] <= 8'hFE;
            reg_file[10824] <= 8'h63;
            reg_file[10825] <= 8'h90;
            reg_file[10826] <= 8'h06;
            reg_file[10827] <= 8'h02;
            reg_file[10828] <= 8'h93;
            reg_file[10829] <= 8'h07;
            reg_file[10830] <= 8'h07;
            reg_file[10831] <= 8'h00;
            reg_file[10832] <= 8'h13;
            reg_file[10833] <= 8'h05;
            reg_file[10834] <= 8'h06;
            reg_file[10835] <= 8'h00;
            reg_file[10836] <= 8'h93;
            reg_file[10837] <= 8'h08;
            reg_file[10838] <= 8'h00;
            reg_file[10839] <= 8'h00;
            reg_file[10840] <= 8'h13;
            reg_file[10841] <= 8'h08;
            reg_file[10842] <= 8'hF0;
            reg_file[10843] <= 8'h7F;
            reg_file[10844] <= 8'h6F;
            reg_file[10845] <= 8'hF0;
            reg_file[10846] <= 8'h1F;
            reg_file[10847] <= 8'hF9;
            reg_file[10848] <= 8'h13;
            reg_file[10849] <= 8'h04;
            reg_file[10850] <= 8'h00;
            reg_file[10851] <= 8'h00;
            reg_file[10852] <= 8'h6F;
            reg_file[10853] <= 8'hF0;
            reg_file[10854] <= 8'h5F;
            reg_file[10855] <= 8'hFC;
            reg_file[10856] <= 8'h33;
            reg_file[10857] <= 8'h67;
            reg_file[10858] <= 8'hC7;
            reg_file[10859] <= 8'h00;
            reg_file[10860] <= 8'hE3;
            reg_file[10861] <= 8'h04;
            reg_file[10862] <= 8'h07;
            reg_file[10863] <= 8'hFE;
            reg_file[10864] <= 8'h93;
            reg_file[10865] <= 8'h04;
            reg_file[10866] <= 8'h00;
            reg_file[10867] <= 8'h00;
            reg_file[10868] <= 8'hB7;
            reg_file[10869] <= 8'h07;
            reg_file[10870] <= 8'h40;
            reg_file[10871] <= 8'h00;
            reg_file[10872] <= 8'h13;
            reg_file[10873] <= 8'h05;
            reg_file[10874] <= 8'h00;
            reg_file[10875] <= 8'h00;
            reg_file[10876] <= 8'h13;
            reg_file[10877] <= 8'h08;
            reg_file[10878] <= 8'hF0;
            reg_file[10879] <= 8'h7F;
            reg_file[10880] <= 8'h13;
            reg_file[10881] <= 8'h97;
            reg_file[10882] <= 8'h87;
            reg_file[10883] <= 8'h00;
            reg_file[10884] <= 8'h63;
            reg_file[10885] <= 8'h5E;
            reg_file[10886] <= 8'h07;
            reg_file[10887] <= 8'h00;
            reg_file[10888] <= 8'h13;
            reg_file[10889] <= 8'h08;
            reg_file[10890] <= 8'h18;
            reg_file[10891] <= 8'h00;
            reg_file[10892] <= 8'h13;
            reg_file[10893] <= 8'h07;
            reg_file[10894] <= 8'hF0;
            reg_file[10895] <= 8'h7F;
            reg_file[10896] <= 8'h63;
            reg_file[10897] <= 8'h08;
            reg_file[10898] <= 8'hE8;
            reg_file[10899] <= 8'h70;
            reg_file[10900] <= 8'h37;
            reg_file[10901] <= 8'h07;
            reg_file[10902] <= 8'h80;
            reg_file[10903] <= 8'hFF;
            reg_file[10904] <= 8'h13;
            reg_file[10905] <= 8'h07;
            reg_file[10906] <= 8'hF7;
            reg_file[10907] <= 8'hFF;
            reg_file[10908] <= 8'hB3;
            reg_file[10909] <= 8'hF7;
            reg_file[10910] <= 8'hE7;
            reg_file[10911] <= 8'h00;
            reg_file[10912] <= 8'h13;
            reg_file[10913] <= 8'h97;
            reg_file[10914] <= 8'hD7;
            reg_file[10915] <= 8'h01;
            reg_file[10916] <= 8'h13;
            reg_file[10917] <= 8'h55;
            reg_file[10918] <= 8'h35;
            reg_file[10919] <= 8'h00;
            reg_file[10920] <= 8'h33;
            reg_file[10921] <= 8'h65;
            reg_file[10922] <= 8'hA7;
            reg_file[10923] <= 8'h00;
            reg_file[10924] <= 8'h13;
            reg_file[10925] <= 8'h07;
            reg_file[10926] <= 8'hF0;
            reg_file[10927] <= 8'h7F;
            reg_file[10928] <= 8'h93;
            reg_file[10929] <= 8'hD7;
            reg_file[10930] <= 8'h37;
            reg_file[10931] <= 8'h00;
            reg_file[10932] <= 8'h63;
            reg_file[10933] <= 8'h1E;
            reg_file[10934] <= 8'hE8;
            reg_file[10935] <= 8'h00;
            reg_file[10936] <= 8'h33;
            reg_file[10937] <= 8'h65;
            reg_file[10938] <= 8'hF5;
            reg_file[10939] <= 8'h00;
            reg_file[10940] <= 8'h93;
            reg_file[10941] <= 8'h07;
            reg_file[10942] <= 8'h00;
            reg_file[10943] <= 8'h00;
            reg_file[10944] <= 8'h63;
            reg_file[10945] <= 8'h08;
            reg_file[10946] <= 8'h05;
            reg_file[10947] <= 8'h00;
            reg_file[10948] <= 8'hB7;
            reg_file[10949] <= 8'h07;
            reg_file[10950] <= 8'h08;
            reg_file[10951] <= 8'h00;
            reg_file[10952] <= 8'h13;
            reg_file[10953] <= 8'h05;
            reg_file[10954] <= 8'h00;
            reg_file[10955] <= 8'h00;
            reg_file[10956] <= 8'h93;
            reg_file[10957] <= 8'h04;
            reg_file[10958] <= 8'h00;
            reg_file[10959] <= 8'h00;
            reg_file[10960] <= 8'h37;
            reg_file[10961] <= 8'h07;
            reg_file[10962] <= 8'hF0;
            reg_file[10963] <= 8'h7F;
            reg_file[10964] <= 8'h13;
            reg_file[10965] <= 8'h18;
            reg_file[10966] <= 8'h48;
            reg_file[10967] <= 8'h01;
            reg_file[10968] <= 8'h93;
            reg_file[10969] <= 8'h97;
            reg_file[10970] <= 8'hC7;
            reg_file[10971] <= 8'h00;
            reg_file[10972] <= 8'h33;
            reg_file[10973] <= 8'h78;
            reg_file[10974] <= 8'hE8;
            reg_file[10975] <= 8'h00;
            reg_file[10976] <= 8'h93;
            reg_file[10977] <= 8'hD7;
            reg_file[10978] <= 8'hC7;
            reg_file[10979] <= 8'h00;
            reg_file[10980] <= 8'hB3;
            reg_file[10981] <= 8'h67;
            reg_file[10982] <= 8'hF8;
            reg_file[10983] <= 8'h00;
            reg_file[10984] <= 8'h93;
            reg_file[10985] <= 8'h94;
            reg_file[10986] <= 8'hF4;
            reg_file[10987] <= 8'h01;
            reg_file[10988] <= 8'h33;
            reg_file[10989] <= 8'hE7;
            reg_file[10990] <= 8'h97;
            reg_file[10991] <= 8'h00;
            reg_file[10992] <= 8'h93;
            reg_file[10993] <= 8'h05;
            reg_file[10994] <= 8'h07;
            reg_file[10995] <= 8'h00;
            reg_file[10996] <= 8'h63;
            reg_file[10997] <= 8'h04;
            reg_file[10998] <= 8'h04;
            reg_file[10999] <= 8'h00;
            reg_file[11000] <= 8'h73;
            reg_file[11001] <= 8'h20;
            reg_file[11002] <= 8'h14;
            reg_file[11003] <= 8'h00;
            reg_file[11004] <= 8'h83;
            reg_file[11005] <= 8'h20;
            reg_file[11006] <= 8'hC1;
            reg_file[11007] <= 8'h01;
            reg_file[11008] <= 8'h03;
            reg_file[11009] <= 8'h24;
            reg_file[11010] <= 8'h81;
            reg_file[11011] <= 8'h01;
            reg_file[11012] <= 8'h83;
            reg_file[11013] <= 8'h24;
            reg_file[11014] <= 8'h41;
            reg_file[11015] <= 8'h01;
            reg_file[11016] <= 8'h03;
            reg_file[11017] <= 8'h29;
            reg_file[11018] <= 8'h01;
            reg_file[11019] <= 8'h01;
            reg_file[11020] <= 8'h83;
            reg_file[11021] <= 8'h29;
            reg_file[11022] <= 8'hC1;
            reg_file[11023] <= 8'h00;
            reg_file[11024] <= 8'h03;
            reg_file[11025] <= 8'h2A;
            reg_file[11026] <= 8'h81;
            reg_file[11027] <= 8'h00;
            reg_file[11028] <= 8'h13;
            reg_file[11029] <= 8'h01;
            reg_file[11030] <= 8'h01;
            reg_file[11031] <= 8'h02;
            reg_file[11032] <= 8'h67;
            reg_file[11033] <= 8'h80;
            reg_file[11034] <= 8'h00;
            reg_file[11035] <= 8'h00;
            reg_file[11036] <= 8'h93;
            reg_file[11037] <= 8'h06;
            reg_file[11038] <= 8'hF0;
            reg_file[11039] <= 8'h7F;
            reg_file[11040] <= 8'h63;
            reg_file[11041] <= 8'h08;
            reg_file[11042] <= 8'hD8;
            reg_file[11043] <= 8'h02;
            reg_file[11044] <= 8'h33;
            reg_file[11045] <= 8'h06;
            reg_file[11046] <= 8'hC5;
            reg_file[11047] <= 8'h00;
            reg_file[11048] <= 8'h33;
            reg_file[11049] <= 8'h35;
            reg_file[11050] <= 8'hA6;
            reg_file[11051] <= 8'h00;
            reg_file[11052] <= 8'hB3;
            reg_file[11053] <= 8'h87;
            reg_file[11054] <= 8'hE7;
            reg_file[11055] <= 8'h00;
            reg_file[11056] <= 8'hB3;
            reg_file[11057] <= 8'h87;
            reg_file[11058] <= 8'hA7;
            reg_file[11059] <= 8'h00;
            reg_file[11060] <= 8'h13;
            reg_file[11061] <= 8'h95;
            reg_file[11062] <= 8'hF7;
            reg_file[11063] <= 8'h01;
            reg_file[11064] <= 8'h13;
            reg_file[11065] <= 8'h56;
            reg_file[11066] <= 8'h16;
            reg_file[11067] <= 8'h00;
            reg_file[11068] <= 8'h33;
            reg_file[11069] <= 8'h65;
            reg_file[11070] <= 8'hC5;
            reg_file[11071] <= 8'h00;
            reg_file[11072] <= 8'h93;
            reg_file[11073] <= 8'hD7;
            reg_file[11074] <= 8'h17;
            reg_file[11075] <= 8'h00;
            reg_file[11076] <= 8'h93;
            reg_file[11077] <= 8'h08;
            reg_file[11078] <= 8'h00;
            reg_file[11079] <= 8'h00;
            reg_file[11080] <= 8'h13;
            reg_file[11081] <= 8'h04;
            reg_file[11082] <= 8'h00;
            reg_file[11083] <= 8'h00;
            reg_file[11084] <= 8'h6F;
            reg_file[11085] <= 8'hF0;
            reg_file[11086] <= 8'h1F;
            reg_file[11087] <= 8'hEA;
            reg_file[11088] <= 8'h63;
            reg_file[11089] <= 8'h88;
            reg_file[11090] <= 8'h09;
            reg_file[11091] <= 8'h00;
            reg_file[11092] <= 8'h93;
            reg_file[11093] <= 8'h07;
            reg_file[11094] <= 8'h30;
            reg_file[11095] <= 8'h00;
            reg_file[11096] <= 8'h63;
            reg_file[11097] <= 8'h98;
            reg_file[11098] <= 8'hF9;
            reg_file[11099] <= 8'h00;
            reg_file[11100] <= 8'h63;
            reg_file[11101] <= 8'h9C;
            reg_file[11102] <= 8'h04;
            reg_file[11103] <= 8'h00;
            reg_file[11104] <= 8'h13;
            reg_file[11105] <= 8'h08;
            reg_file[11106] <= 8'hF0;
            reg_file[11107] <= 8'h7F;
            reg_file[11108] <= 8'h6F;
            reg_file[11109] <= 8'h00;
            reg_file[11110] <= 8'hC0;
            reg_file[11111] <= 8'h06;
            reg_file[11112] <= 8'h93;
            reg_file[11113] <= 8'h07;
            reg_file[11114] <= 8'h20;
            reg_file[11115] <= 8'h00;
            reg_file[11116] <= 8'h63;
            reg_file[11117] <= 8'h94;
            reg_file[11118] <= 8'hF9;
            reg_file[11119] <= 8'h00;
            reg_file[11120] <= 8'hE3;
            reg_file[11121] <= 8'h98;
            reg_file[11122] <= 8'h04;
            reg_file[11123] <= 8'hFE;
            reg_file[11124] <= 8'h93;
            reg_file[11125] <= 8'h08;
            reg_file[11126] <= 8'h00;
            reg_file[11127] <= 8'h00;
            reg_file[11128] <= 8'h93;
            reg_file[11129] <= 8'h07;
            reg_file[11130] <= 8'hF0;
            reg_file[11131] <= 8'hFF;
            reg_file[11132] <= 8'h13;
            reg_file[11133] <= 8'h05;
            reg_file[11134] <= 8'hF0;
            reg_file[11135] <= 8'hFF;
            reg_file[11136] <= 8'h13;
            reg_file[11137] <= 8'h08;
            reg_file[11138] <= 8'hE0;
            reg_file[11139] <= 8'h7F;
            reg_file[11140] <= 8'h13;
            reg_file[11141] <= 8'h04;
            reg_file[11142] <= 8'h50;
            reg_file[11143] <= 8'h00;
            reg_file[11144] <= 8'h13;
            reg_file[11145] <= 8'h07;
            reg_file[11146] <= 8'h20;
            reg_file[11147] <= 8'h00;
            reg_file[11148] <= 8'h13;
            reg_file[11149] <= 8'h64;
            reg_file[11150] <= 8'h14;
            reg_file[11151] <= 8'h00;
            reg_file[11152] <= 8'h63;
            reg_file[11153] <= 8'h82;
            reg_file[11154] <= 8'hE9;
            reg_file[11155] <= 8'h60;
            reg_file[11156] <= 8'h13;
            reg_file[11157] <= 8'h07;
            reg_file[11158] <= 8'h30;
            reg_file[11159] <= 8'h00;
            reg_file[11160] <= 8'h63;
            reg_file[11161] <= 8'h88;
            reg_file[11162] <= 8'hE9;
            reg_file[11163] <= 8'h5E;
            reg_file[11164] <= 8'h63;
            reg_file[11165] <= 8'h9E;
            reg_file[11166] <= 8'h09;
            reg_file[11167] <= 8'h5E;
            reg_file[11168] <= 8'h13;
            reg_file[11169] <= 8'h77;
            reg_file[11170] <= 8'hF5;
            reg_file[11171] <= 8'h00;
            reg_file[11172] <= 8'h93;
            reg_file[11173] <= 8'h06;
            reg_file[11174] <= 8'h40;
            reg_file[11175] <= 8'h00;
            reg_file[11176] <= 8'h63;
            reg_file[11177] <= 8'h08;
            reg_file[11178] <= 8'hD7;
            reg_file[11179] <= 8'h5E;
            reg_file[11180] <= 8'h13;
            reg_file[11181] <= 8'h07;
            reg_file[11182] <= 8'h45;
            reg_file[11183] <= 8'h00;
            reg_file[11184] <= 8'h33;
            reg_file[11185] <= 8'h35;
            reg_file[11186] <= 8'hA7;
            reg_file[11187] <= 8'h00;
            reg_file[11188] <= 8'hB3;
            reg_file[11189] <= 8'h87;
            reg_file[11190] <= 8'hA7;
            reg_file[11191] <= 8'h00;
            reg_file[11192] <= 8'h13;
            reg_file[11193] <= 8'h05;
            reg_file[11194] <= 8'h07;
            reg_file[11195] <= 8'h00;
            reg_file[11196] <= 8'h6F;
            reg_file[11197] <= 8'h00;
            reg_file[11198] <= 8'hC0;
            reg_file[11199] <= 8'h5D;
            reg_file[11200] <= 8'h63;
            reg_file[11201] <= 8'h88;
            reg_file[11202] <= 8'h09;
            reg_file[11203] <= 8'h00;
            reg_file[11204] <= 8'h93;
            reg_file[11205] <= 8'h07;
            reg_file[11206] <= 8'h30;
            reg_file[11207] <= 8'h00;
            reg_file[11208] <= 8'h63;
            reg_file[11209] <= 8'h9C;
            reg_file[11210] <= 8'hF9;
            reg_file[11211] <= 8'h00;
            reg_file[11212] <= 8'h63;
            reg_file[11213] <= 8'h9C;
            reg_file[11214] <= 8'h04;
            reg_file[11215] <= 8'h50;
            reg_file[11216] <= 8'h93;
            reg_file[11217] <= 8'h07;
            reg_file[11218] <= 8'h00;
            reg_file[11219] <= 8'h00;
            reg_file[11220] <= 8'h13;
            reg_file[11221] <= 8'h05;
            reg_file[11222] <= 8'h00;
            reg_file[11223] <= 8'h00;
            reg_file[11224] <= 8'h13;
            reg_file[11225] <= 8'h04;
            reg_file[11226] <= 8'h50;
            reg_file[11227] <= 8'h00;
            reg_file[11228] <= 8'h6F;
            reg_file[11229] <= 8'hF0;
            reg_file[11230] <= 8'h5F;
            reg_file[11231] <= 8'hEA;
            reg_file[11232] <= 8'h93;
            reg_file[11233] <= 8'h07;
            reg_file[11234] <= 8'h20;
            reg_file[11235] <= 8'h00;
            reg_file[11236] <= 8'h63;
            reg_file[11237] <= 8'h90;
            reg_file[11238] <= 8'hF9;
            reg_file[11239] <= 8'h50;
            reg_file[11240] <= 8'hE3;
            reg_file[11241] <= 8'h94;
            reg_file[11242] <= 8'h04;
            reg_file[11243] <= 8'hFE;
            reg_file[11244] <= 8'h6F;
            reg_file[11245] <= 8'hF0;
            reg_file[11246] <= 8'h9F;
            reg_file[11247] <= 8'hF8;
            reg_file[11248] <= 8'h63;
            reg_file[11249] <= 8'h5C;
            reg_file[11250] <= 8'h00;
            reg_file[11251] <= 8'h0F;
            reg_file[11252] <= 8'h63;
            reg_file[11253] <= 8'h9E;
            reg_file[11254] <= 8'h08;
            reg_file[11255] <= 8'h08;
            reg_file[11256] <= 8'hB3;
            reg_file[11257] <= 8'h66;
            reg_file[11258] <= 8'hC7;
            reg_file[11259] <= 8'h00;
            reg_file[11260] <= 8'hE3;
            reg_file[11261] <= 8'h86;
            reg_file[11262] <= 8'h06;
            reg_file[11263] <= 8'hB0;
            reg_file[11264] <= 8'h93;
            reg_file[11265] <= 8'h06;
            reg_file[11266] <= 8'hF8;
            reg_file[11267] <= 8'hFF;
            reg_file[11268] <= 8'h63;
            reg_file[11269] <= 8'h9E;
            reg_file[11270] <= 8'h06;
            reg_file[11271] <= 8'h00;
            reg_file[11272] <= 8'h33;
            reg_file[11273] <= 8'h06;
            reg_file[11274] <= 8'hC5;
            reg_file[11275] <= 8'h40;
            reg_file[11276] <= 8'hB3;
            reg_file[11277] <= 8'h87;
            reg_file[11278] <= 8'hE7;
            reg_file[11279] <= 8'h40;
            reg_file[11280] <= 8'hB3;
            reg_file[11281] <= 8'h36;
            reg_file[11282] <= 8'hC5;
            reg_file[11283] <= 8'h00;
            reg_file[11284] <= 8'h33;
            reg_file[11285] <= 8'h87;
            reg_file[11286] <= 8'hD7;
            reg_file[11287] <= 8'h40;
            reg_file[11288] <= 8'h13;
            reg_file[11289] <= 8'h08;
            reg_file[11290] <= 8'h10;
            reg_file[11291] <= 8'h00;
            reg_file[11292] <= 8'h6F;
            reg_file[11293] <= 8'h00;
            reg_file[11294] <= 8'h40;
            reg_file[11295] <= 8'h05;
            reg_file[11296] <= 8'h93;
            reg_file[11297] <= 8'h05;
            reg_file[11298] <= 8'hF0;
            reg_file[11299] <= 8'h7F;
            reg_file[11300] <= 8'hE3;
            reg_file[11301] <= 8'h0A;
            reg_file[11302] <= 8'hB8;
            reg_file[11303] <= 8'hB2;
            reg_file[11304] <= 8'h93;
            reg_file[11305] <= 8'h05;
            reg_file[11306] <= 8'h80;
            reg_file[11307] <= 8'h03;
            reg_file[11308] <= 8'h63;
            reg_file[11309] <= 8'hC8;
            reg_file[11310] <= 8'hD5;
            reg_file[11311] <= 8'h0A;
            reg_file[11312] <= 8'h93;
            reg_file[11313] <= 8'h05;
            reg_file[11314] <= 8'hF0;
            reg_file[11315] <= 8'h01;
            reg_file[11316] <= 8'h63;
            reg_file[11317] <= 8'hCA;
            reg_file[11318] <= 8'hD5;
            reg_file[11319] <= 8'h06;
            reg_file[11320] <= 8'h13;
            reg_file[11321] <= 8'h08;
            reg_file[11322] <= 8'h00;
            reg_file[11323] <= 8'h02;
            reg_file[11324] <= 8'h33;
            reg_file[11325] <= 8'h08;
            reg_file[11326] <= 8'hD8;
            reg_file[11327] <= 8'h40;
            reg_file[11328] <= 8'hB3;
            reg_file[11329] <= 8'h58;
            reg_file[11330] <= 8'hD6;
            reg_file[11331] <= 8'h00;
            reg_file[11332] <= 8'hB3;
            reg_file[11333] <= 8'h15;
            reg_file[11334] <= 8'h07;
            reg_file[11335] <= 8'h01;
            reg_file[11336] <= 8'h33;
            reg_file[11337] <= 8'h16;
            reg_file[11338] <= 8'h06;
            reg_file[11339] <= 8'h01;
            reg_file[11340] <= 8'hB3;
            reg_file[11341] <= 8'hE5;
            reg_file[11342] <= 8'h15;
            reg_file[11343] <= 8'h01;
            reg_file[11344] <= 8'h33;
            reg_file[11345] <= 8'h36;
            reg_file[11346] <= 8'hC0;
            reg_file[11347] <= 8'h00;
            reg_file[11348] <= 8'h33;
            reg_file[11349] <= 8'hE6;
            reg_file[11350] <= 8'hC5;
            reg_file[11351] <= 8'h00;
            reg_file[11352] <= 8'hB3;
            reg_file[11353] <= 8'h56;
            reg_file[11354] <= 8'hD7;
            reg_file[11355] <= 8'h00;
            reg_file[11356] <= 8'h33;
            reg_file[11357] <= 8'h06;
            reg_file[11358] <= 8'hC5;
            reg_file[11359] <= 8'h40;
            reg_file[11360] <= 8'hB3;
            reg_file[11361] <= 8'h86;
            reg_file[11362] <= 8'hD7;
            reg_file[11363] <= 8'h40;
            reg_file[11364] <= 8'hB3;
            reg_file[11365] <= 8'h37;
            reg_file[11366] <= 8'hC5;
            reg_file[11367] <= 8'h00;
            reg_file[11368] <= 8'h33;
            reg_file[11369] <= 8'h87;
            reg_file[11370] <= 8'hF6;
            reg_file[11371] <= 8'h40;
            reg_file[11372] <= 8'h13;
            reg_file[11373] <= 8'h08;
            reg_file[11374] <= 8'h04;
            reg_file[11375] <= 8'h00;
            reg_file[11376] <= 8'h93;
            reg_file[11377] <= 8'h17;
            reg_file[11378] <= 8'h87;
            reg_file[11379] <= 8'h00;
            reg_file[11380] <= 8'hE3;
            reg_file[11381] <= 8'hD4;
            reg_file[11382] <= 8'h07;
            reg_file[11383] <= 8'hC0;
            reg_file[11384] <= 8'h37;
            reg_file[11385] <= 8'h09;
            reg_file[11386] <= 8'h80;
            reg_file[11387] <= 8'h00;
            reg_file[11388] <= 8'h13;
            reg_file[11389] <= 8'h09;
            reg_file[11390] <= 8'hF9;
            reg_file[11391] <= 8'hFF;
            reg_file[11392] <= 8'h33;
            reg_file[11393] <= 8'h79;
            reg_file[11394] <= 8'h27;
            reg_file[11395] <= 8'h01;
            reg_file[11396] <= 8'h13;
            reg_file[11397] <= 8'h0A;
            reg_file[11398] <= 8'h06;
            reg_file[11399] <= 8'h00;
            reg_file[11400] <= 8'h13;
            reg_file[11401] <= 8'h04;
            reg_file[11402] <= 8'h08;
            reg_file[11403] <= 8'h00;
            reg_file[11404] <= 8'h6F;
            reg_file[11405] <= 8'h00;
            reg_file[11406] <= 8'h40;
            reg_file[11407] <= 8'h30;
            reg_file[11408] <= 8'h93;
            reg_file[11409] <= 8'h06;
            reg_file[11410] <= 8'hF0;
            reg_file[11411] <= 8'h7F;
            reg_file[11412] <= 8'hE3;
            reg_file[11413] <= 8'h02;
            reg_file[11414] <= 8'hD4;
            reg_file[11415] <= 8'hAE;
            reg_file[11416] <= 8'hB7;
            reg_file[11417] <= 8'h06;
            reg_file[11418] <= 8'h80;
            reg_file[11419] <= 8'h00;
            reg_file[11420] <= 8'h33;
            reg_file[11421] <= 8'h67;
            reg_file[11422] <= 8'hD7;
            reg_file[11423] <= 8'h00;
            reg_file[11424] <= 8'h93;
            reg_file[11425] <= 8'h06;
            reg_file[11426] <= 8'h08;
            reg_file[11427] <= 8'h00;
            reg_file[11428] <= 8'h6F;
            reg_file[11429] <= 8'hF0;
            reg_file[11430] <= 8'h5F;
            reg_file[11431] <= 8'hF8;
            reg_file[11432] <= 8'h93;
            reg_file[11433] <= 8'h85;
            reg_file[11434] <= 8'h06;
            reg_file[11435] <= 8'hFE;
            reg_file[11436] <= 8'h93;
            reg_file[11437] <= 8'h08;
            reg_file[11438] <= 8'h00;
            reg_file[11439] <= 8'h02;
            reg_file[11440] <= 8'hB3;
            reg_file[11441] <= 8'h55;
            reg_file[11442] <= 8'hB7;
            reg_file[11443] <= 8'h00;
            reg_file[11444] <= 8'h13;
            reg_file[11445] <= 8'h08;
            reg_file[11446] <= 8'h00;
            reg_file[11447] <= 8'h00;
            reg_file[11448] <= 8'h63;
            reg_file[11449] <= 8'h88;
            reg_file[11450] <= 8'h16;
            reg_file[11451] <= 8'h01;
            reg_file[11452] <= 8'h13;
            reg_file[11453] <= 8'h08;
            reg_file[11454] <= 8'h00;
            reg_file[11455] <= 8'h04;
            reg_file[11456] <= 8'hB3;
            reg_file[11457] <= 8'h06;
            reg_file[11458] <= 8'hD8;
            reg_file[11459] <= 8'h40;
            reg_file[11460] <= 8'h33;
            reg_file[11461] <= 8'h18;
            reg_file[11462] <= 8'hD7;
            reg_file[11463] <= 8'h00;
            reg_file[11464] <= 8'h33;
            reg_file[11465] <= 8'h66;
            reg_file[11466] <= 8'hC8;
            reg_file[11467] <= 8'h00;
            reg_file[11468] <= 8'h33;
            reg_file[11469] <= 8'h36;
            reg_file[11470] <= 8'hC0;
            reg_file[11471] <= 8'h00;
            reg_file[11472] <= 8'h33;
            reg_file[11473] <= 8'hE6;
            reg_file[11474] <= 8'hC5;
            reg_file[11475] <= 8'h00;
            reg_file[11476] <= 8'h93;
            reg_file[11477] <= 8'h06;
            reg_file[11478] <= 8'h00;
            reg_file[11479] <= 8'h00;
            reg_file[11480] <= 8'h6F;
            reg_file[11481] <= 8'hF0;
            reg_file[11482] <= 8'h5F;
            reg_file[11483] <= 8'hF8;
            reg_file[11484] <= 8'h33;
            reg_file[11485] <= 8'h66;
            reg_file[11486] <= 8'hC7;
            reg_file[11487] <= 8'h00;
            reg_file[11488] <= 8'h33;
            reg_file[11489] <= 8'h36;
            reg_file[11490] <= 8'hC0;
            reg_file[11491] <= 8'h00;
            reg_file[11492] <= 8'h6F;
            reg_file[11493] <= 8'hF0;
            reg_file[11494] <= 8'h1F;
            reg_file[11495] <= 8'hFF;
            reg_file[11496] <= 8'h63;
            reg_file[11497] <= 8'h0A;
            reg_file[11498] <= 8'h08;
            reg_file[11499] <= 8'h12;
            reg_file[11500] <= 8'h33;
            reg_file[11501] <= 8'h88;
            reg_file[11502] <= 8'h88;
            reg_file[11503] <= 8'h40;
            reg_file[11504] <= 8'h63;
            reg_file[11505] <= 8'h12;
            reg_file[11506] <= 8'h04;
            reg_file[11507] <= 8'h06;
            reg_file[11508] <= 8'hB3;
            reg_file[11509] <= 8'hE5;
            reg_file[11510] <= 8'hA7;
            reg_file[11511] <= 8'h00;
            reg_file[11512] <= 8'h63;
            reg_file[11513] <= 8'h98;
            reg_file[11514] <= 8'h05;
            reg_file[11515] <= 8'h00;
            reg_file[11516] <= 8'h93;
            reg_file[11517] <= 8'h07;
            reg_file[11518] <= 8'hF0;
            reg_file[11519] <= 8'h7F;
            reg_file[11520] <= 8'h93;
            reg_file[11521] <= 8'h84;
            reg_file[11522] <= 8'h06;
            reg_file[11523] <= 8'h00;
            reg_file[11524] <= 8'h6F;
            reg_file[11525] <= 8'hF0;
            reg_file[11526] <= 8'h5F;
            reg_file[11527] <= 8'hB7;
            reg_file[11528] <= 8'h13;
            reg_file[11529] <= 8'h03;
            reg_file[11530] <= 8'hF8;
            reg_file[11531] <= 8'hFF;
            reg_file[11532] <= 8'h63;
            reg_file[11533] <= 8'h10;
            reg_file[11534] <= 8'h03;
            reg_file[11535] <= 8'h02;
            reg_file[11536] <= 8'hB3;
            reg_file[11537] <= 8'h05;
            reg_file[11538] <= 8'hA6;
            reg_file[11539] <= 8'h40;
            reg_file[11540] <= 8'h33;
            reg_file[11541] <= 8'h36;
            reg_file[11542] <= 8'hB6;
            reg_file[11543] <= 8'h00;
            reg_file[11544] <= 8'hB3;
            reg_file[11545] <= 8'h07;
            reg_file[11546] <= 8'hF7;
            reg_file[11547] <= 8'h40;
            reg_file[11548] <= 8'h33;
            reg_file[11549] <= 8'h87;
            reg_file[11550] <= 8'hC7;
            reg_file[11551] <= 8'h40;
            reg_file[11552] <= 8'h93;
            reg_file[11553] <= 8'h84;
            reg_file[11554] <= 8'h06;
            reg_file[11555] <= 8'h00;
            reg_file[11556] <= 8'h13;
            reg_file[11557] <= 8'h86;
            reg_file[11558] <= 8'h05;
            reg_file[11559] <= 8'h00;
            reg_file[11560] <= 8'h6F;
            reg_file[11561] <= 8'hF0;
            reg_file[11562] <= 8'h1F;
            reg_file[11563] <= 8'hEF;
            reg_file[11564] <= 8'h93;
            reg_file[11565] <= 8'h05;
            reg_file[11566] <= 8'hF0;
            reg_file[11567] <= 8'h7F;
            reg_file[11568] <= 8'h63;
            reg_file[11569] <= 8'h1C;
            reg_file[11570] <= 8'hB8;
            reg_file[11571] <= 8'h04;
            reg_file[11572] <= 8'h33;
            reg_file[11573] <= 8'h65;
            reg_file[11574] <= 8'hC7;
            reg_file[11575] <= 8'h00;
            reg_file[11576] <= 8'h63;
            reg_file[11577] <= 8'h04;
            reg_file[11578] <= 8'h05;
            reg_file[11579] <= 8'h3E;
            reg_file[11580] <= 8'h93;
            reg_file[11581] <= 8'h17;
            reg_file[11582] <= 8'h97;
            reg_file[11583] <= 8'h00;
            reg_file[11584] <= 8'h63;
            reg_file[11585] <= 8'hC6;
            reg_file[11586] <= 8'h07;
            reg_file[11587] <= 8'h3E;
            reg_file[11588] <= 8'h93;
            reg_file[11589] <= 8'h07;
            reg_file[11590] <= 8'h07;
            reg_file[11591] <= 8'h00;
            reg_file[11592] <= 8'h13;
            reg_file[11593] <= 8'h05;
            reg_file[11594] <= 8'h06;
            reg_file[11595] <= 8'h00;
            reg_file[11596] <= 8'h93;
            reg_file[11597] <= 8'h84;
            reg_file[11598] <= 8'h06;
            reg_file[11599] <= 8'h00;
            reg_file[11600] <= 8'h6F;
            reg_file[11601] <= 8'hF0;
            reg_file[11602] <= 8'h9F;
            reg_file[11603] <= 8'hBA;
            reg_file[11604] <= 8'h93;
            reg_file[11605] <= 8'h05;
            reg_file[11606] <= 8'hF0;
            reg_file[11607] <= 8'h7F;
            reg_file[11608] <= 8'h63;
            reg_file[11609] <= 8'h92;
            reg_file[11610] <= 8'hB8;
            reg_file[11611] <= 8'h02;
            reg_file[11612] <= 8'h33;
            reg_file[11613] <= 8'h65;
            reg_file[11614] <= 8'hC7;
            reg_file[11615] <= 8'h00;
            reg_file[11616] <= 8'h63;
            reg_file[11617] <= 8'h0E;
            reg_file[11618] <= 8'h05;
            reg_file[11619] <= 8'h3C;
            reg_file[11620] <= 8'h93;
            reg_file[11621] <= 8'h17;
            reg_file[11622] <= 8'h97;
            reg_file[11623] <= 8'h00;
            reg_file[11624] <= 8'h63;
            reg_file[11625] <= 8'hC2;
            reg_file[11626] <= 8'h07;
            reg_file[11627] <= 8'h3E;
            reg_file[11628] <= 8'h93;
            reg_file[11629] <= 8'h07;
            reg_file[11630] <= 8'h07;
            reg_file[11631] <= 8'h00;
            reg_file[11632] <= 8'h13;
            reg_file[11633] <= 8'h05;
            reg_file[11634] <= 8'h06;
            reg_file[11635] <= 8'h00;
            reg_file[11636] <= 8'h13;
            reg_file[11637] <= 8'h08;
            reg_file[11638] <= 8'hF0;
            reg_file[11639] <= 8'h7F;
            reg_file[11640] <= 8'h6F;
            reg_file[11641] <= 8'hF0;
            reg_file[11642] <= 8'h5F;
            reg_file[11643] <= 8'hFD;
            reg_file[11644] <= 8'hB7;
            reg_file[11645] <= 8'h05;
            reg_file[11646] <= 8'h80;
            reg_file[11647] <= 8'h00;
            reg_file[11648] <= 8'hB3;
            reg_file[11649] <= 8'hE7;
            reg_file[11650] <= 8'hB7;
            reg_file[11651] <= 8'h00;
            reg_file[11652] <= 8'h13;
            reg_file[11653] <= 8'h03;
            reg_file[11654] <= 8'h08;
            reg_file[11655] <= 8'h00;
            reg_file[11656] <= 8'h93;
            reg_file[11657] <= 8'h05;
            reg_file[11658] <= 8'h80;
            reg_file[11659] <= 8'h03;
            reg_file[11660] <= 8'h63;
            reg_file[11661] <= 8'hC2;
            reg_file[11662] <= 8'h65;
            reg_file[11663] <= 8'h08;
            reg_file[11664] <= 8'h93;
            reg_file[11665] <= 8'h05;
            reg_file[11666] <= 8'hF0;
            reg_file[11667] <= 8'h01;
            reg_file[11668] <= 8'h63;
            reg_file[11669] <= 8'hC4;
            reg_file[11670] <= 8'h65;
            reg_file[11671] <= 8'h04;
            reg_file[11672] <= 8'h13;
            reg_file[11673] <= 8'h08;
            reg_file[11674] <= 8'h00;
            reg_file[11675] <= 8'h02;
            reg_file[11676] <= 8'h33;
            reg_file[11677] <= 8'h08;
            reg_file[11678] <= 8'h68;
            reg_file[11679] <= 8'h40;
            reg_file[11680] <= 8'hB3;
            reg_file[11681] <= 8'h95;
            reg_file[11682] <= 8'h07;
            reg_file[11683] <= 8'h01;
            reg_file[11684] <= 8'h33;
            reg_file[11685] <= 8'h5E;
            reg_file[11686] <= 8'h65;
            reg_file[11687] <= 8'h00;
            reg_file[11688] <= 8'h33;
            reg_file[11689] <= 8'h15;
            reg_file[11690] <= 8'h05;
            reg_file[11691] <= 8'h01;
            reg_file[11692] <= 8'hB3;
            reg_file[11693] <= 8'hE5;
            reg_file[11694] <= 8'hC5;
            reg_file[11695] <= 8'h01;
            reg_file[11696] <= 8'h33;
            reg_file[11697] <= 8'h35;
            reg_file[11698] <= 8'hA0;
            reg_file[11699] <= 8'h00;
            reg_file[11700] <= 8'h33;
            reg_file[11701] <= 8'hE5;
            reg_file[11702] <= 8'hA5;
            reg_file[11703] <= 8'h00;
            reg_file[11704] <= 8'hB3;
            reg_file[11705] <= 8'hD7;
            reg_file[11706] <= 8'h67;
            reg_file[11707] <= 8'h00;
            reg_file[11708] <= 8'hB3;
            reg_file[11709] <= 8'h05;
            reg_file[11710] <= 8'hA6;
            reg_file[11711] <= 8'h40;
            reg_file[11712] <= 8'hB3;
            reg_file[11713] <= 8'h07;
            reg_file[11714] <= 8'hF7;
            reg_file[11715] <= 8'h40;
            reg_file[11716] <= 8'h33;
            reg_file[11717] <= 8'h37;
            reg_file[11718] <= 8'hB6;
            reg_file[11719] <= 8'h00;
            reg_file[11720] <= 8'h33;
            reg_file[11721] <= 8'h87;
            reg_file[11722] <= 8'hE7;
            reg_file[11723] <= 8'h40;
            reg_file[11724] <= 8'h13;
            reg_file[11725] <= 8'h86;
            reg_file[11726] <= 8'h05;
            reg_file[11727] <= 8'h00;
            reg_file[11728] <= 8'h13;
            reg_file[11729] <= 8'h88;
            reg_file[11730] <= 8'h08;
            reg_file[11731] <= 8'h00;
            reg_file[11732] <= 8'h93;
            reg_file[11733] <= 8'h84;
            reg_file[11734] <= 8'h06;
            reg_file[11735] <= 8'h00;
            reg_file[11736] <= 8'h6F;
            reg_file[11737] <= 8'hF0;
            reg_file[11738] <= 8'h9F;
            reg_file[11739] <= 8'hE9;
            reg_file[11740] <= 8'h93;
            reg_file[11741] <= 8'h05;
            reg_file[11742] <= 8'h03;
            reg_file[11743] <= 8'hFE;
            reg_file[11744] <= 8'h13;
            reg_file[11745] <= 8'h0E;
            reg_file[11746] <= 8'h00;
            reg_file[11747] <= 8'h02;
            reg_file[11748] <= 8'hB3;
            reg_file[11749] <= 8'hD5;
            reg_file[11750] <= 8'hB7;
            reg_file[11751] <= 8'h00;
            reg_file[11752] <= 8'h13;
            reg_file[11753] <= 8'h08;
            reg_file[11754] <= 8'h00;
            reg_file[11755] <= 8'h00;
            reg_file[11756] <= 8'h63;
            reg_file[11757] <= 8'h08;
            reg_file[11758] <= 8'hC3;
            reg_file[11759] <= 8'h01;
            reg_file[11760] <= 8'h13;
            reg_file[11761] <= 8'h08;
            reg_file[11762] <= 8'h00;
            reg_file[11763] <= 8'h04;
            reg_file[11764] <= 8'h33;
            reg_file[11765] <= 8'h03;
            reg_file[11766] <= 8'h68;
            reg_file[11767] <= 8'h40;
            reg_file[11768] <= 8'h33;
            reg_file[11769] <= 8'h98;
            reg_file[11770] <= 8'h67;
            reg_file[11771] <= 8'h00;
            reg_file[11772] <= 8'h33;
            reg_file[11773] <= 8'h65;
            reg_file[11774] <= 8'hA8;
            reg_file[11775] <= 8'h00;
            reg_file[11776] <= 8'h33;
            reg_file[11777] <= 8'h35;
            reg_file[11778] <= 8'hA0;
            reg_file[11779] <= 8'h00;
            reg_file[11780] <= 8'h33;
            reg_file[11781] <= 8'hE5;
            reg_file[11782] <= 8'hA5;
            reg_file[11783] <= 8'h00;
            reg_file[11784] <= 8'h93;
            reg_file[11785] <= 8'h07;
            reg_file[11786] <= 8'h00;
            reg_file[11787] <= 8'h00;
            reg_file[11788] <= 8'h6F;
            reg_file[11789] <= 8'hF0;
            reg_file[11790] <= 8'h1F;
            reg_file[11791] <= 8'hFB;
            reg_file[11792] <= 8'h33;
            reg_file[11793] <= 8'hE5;
            reg_file[11794] <= 8'hA7;
            reg_file[11795] <= 8'h00;
            reg_file[11796] <= 8'h33;
            reg_file[11797] <= 8'h35;
            reg_file[11798] <= 8'hA0;
            reg_file[11799] <= 8'h00;
            reg_file[11800] <= 8'h6F;
            reg_file[11801] <= 8'hF0;
            reg_file[11802] <= 8'h1F;
            reg_file[11803] <= 8'hFF;
            reg_file[11804] <= 8'h93;
            reg_file[11805] <= 8'h05;
            reg_file[11806] <= 8'h14;
            reg_file[11807] <= 8'h00;
            reg_file[11808] <= 8'h93;
            reg_file[11809] <= 8'hF5;
            reg_file[11810] <= 8'hE5;
            reg_file[11811] <= 8'h7F;
            reg_file[11812] <= 8'h63;
            reg_file[11813] <= 8'h90;
            reg_file[11814] <= 8'h05;
            reg_file[11815] <= 8'h14;
            reg_file[11816] <= 8'h33;
            reg_file[11817] <= 8'hE3;
            reg_file[11818] <= 8'hA7;
            reg_file[11819] <= 8'h00;
            reg_file[11820] <= 8'hB3;
            reg_file[11821] <= 8'h65;
            reg_file[11822] <= 8'hC7;
            reg_file[11823] <= 8'h00;
            reg_file[11824] <= 8'h63;
            reg_file[11825] <= 8'h18;
            reg_file[11826] <= 8'h04;
            reg_file[11827] <= 8'h0C;
            reg_file[11828] <= 8'h63;
            reg_file[11829] <= 8'h10;
            reg_file[11830] <= 8'h03;
            reg_file[11831] <= 8'h08;
            reg_file[11832] <= 8'h63;
            reg_file[11833] <= 8'h90;
            reg_file[11834] <= 8'h05;
            reg_file[11835] <= 8'h24;
            reg_file[11836] <= 8'h93;
            reg_file[11837] <= 8'h84;
            reg_file[11838] <= 8'hE9;
            reg_file[11839] <= 8'hFF;
            reg_file[11840] <= 8'h93;
            reg_file[11841] <= 8'hB4;
            reg_file[11842] <= 8'h14;
            reg_file[11843] <= 8'h00;
            reg_file[11844] <= 8'h93;
            reg_file[11845] <= 8'h07;
            reg_file[11846] <= 8'h00;
            reg_file[11847] <= 8'h00;
            reg_file[11848] <= 8'h13;
            reg_file[11849] <= 8'h05;
            reg_file[11850] <= 8'h00;
            reg_file[11851] <= 8'h00;
            reg_file[11852] <= 8'h33;
            reg_file[11853] <= 8'h67;
            reg_file[11854] <= 8'hF5;
            reg_file[11855] <= 8'h00;
            reg_file[11856] <= 8'h63;
            reg_file[11857] <= 8'h04;
            reg_file[11858] <= 8'h07;
            reg_file[11859] <= 8'h32;
            reg_file[11860] <= 8'h13;
            reg_file[11861] <= 8'h57;
            reg_file[11862] <= 8'hF5;
            reg_file[11863] <= 8'h01;
            reg_file[11864] <= 8'h93;
            reg_file[11865] <= 8'h98;
            reg_file[11866] <= 8'h17;
            reg_file[11867] <= 8'h00;
            reg_file[11868] <= 8'hB3;
            reg_file[11869] <= 8'h88;
            reg_file[11870] <= 8'hE8;
            reg_file[11871] <= 8'h00;
            reg_file[11872] <= 8'h13;
            reg_file[11873] <= 8'h17;
            reg_file[11874] <= 8'h15;
            reg_file[11875] <= 8'h00;
            reg_file[11876] <= 8'h93;
            reg_file[11877] <= 8'h76;
            reg_file[11878] <= 8'h77;
            reg_file[11879] <= 8'h00;
            reg_file[11880] <= 8'h13;
            reg_file[11881] <= 8'h04;
            reg_file[11882] <= 8'h00;
            reg_file[11883] <= 8'h00;
            reg_file[11884] <= 8'h63;
            reg_file[11885] <= 8'h8A;
            reg_file[11886] <= 8'h06;
            reg_file[11887] <= 8'h02;
            reg_file[11888] <= 8'h93;
            reg_file[11889] <= 8'h06;
            reg_file[11890] <= 8'h20;
            reg_file[11891] <= 8'h00;
            reg_file[11892] <= 8'h63;
            reg_file[11893] <= 8'h8C;
            reg_file[11894] <= 8'hD9;
            reg_file[11895] <= 8'h22;
            reg_file[11896] <= 8'h93;
            reg_file[11897] <= 8'h06;
            reg_file[11898] <= 8'h30;
            reg_file[11899] <= 8'h00;
            reg_file[11900] <= 8'h63;
            reg_file[11901] <= 8'h8A;
            reg_file[11902] <= 8'hD9;
            reg_file[11903] <= 8'h20;
            reg_file[11904] <= 8'h13;
            reg_file[11905] <= 8'h04;
            reg_file[11906] <= 8'h10;
            reg_file[11907] <= 8'h00;
            reg_file[11908] <= 8'h63;
            reg_file[11909] <= 8'h9E;
            reg_file[11910] <= 8'h09;
            reg_file[11911] <= 8'h00;
            reg_file[11912] <= 8'h93;
            reg_file[11913] <= 8'h76;
            reg_file[11914] <= 8'hF7;
            reg_file[11915] <= 8'h00;
            reg_file[11916] <= 8'h13;
            reg_file[11917] <= 8'h06;
            reg_file[11918] <= 8'h40;
            reg_file[11919] <= 8'h00;
            reg_file[11920] <= 8'h63;
            reg_file[11921] <= 8'h88;
            reg_file[11922] <= 8'hC6;
            reg_file[11923] <= 8'h00;
            reg_file[11924] <= 8'h13;
            reg_file[11925] <= 8'h37;
            reg_file[11926] <= 8'hC7;
            reg_file[11927] <= 8'hFF;
            reg_file[11928] <= 8'h13;
            reg_file[11929] <= 8'h47;
            reg_file[11930] <= 8'h17;
            reg_file[11931] <= 8'h00;
            reg_file[11932] <= 8'hB3;
            reg_file[11933] <= 8'h88;
            reg_file[11934] <= 8'hE8;
            reg_file[11935] <= 8'h00;
            reg_file[11936] <= 8'h93;
            reg_file[11937] <= 8'hD8;
            reg_file[11938] <= 8'h88;
            reg_file[11939] <= 8'h01;
            reg_file[11940] <= 8'h93;
            reg_file[11941] <= 8'hC8;
            reg_file[11942] <= 8'h18;
            reg_file[11943] <= 8'h00;
            reg_file[11944] <= 8'h93;
            reg_file[11945] <= 8'hF8;
            reg_file[11946] <= 8'h18;
            reg_file[11947] <= 8'h00;
            reg_file[11948] <= 8'h13;
            reg_file[11949] <= 8'h08;
            reg_file[11950] <= 8'h00;
            reg_file[11951] <= 8'h00;
            reg_file[11952] <= 8'h6F;
            reg_file[11953] <= 8'hF0;
            reg_file[11954] <= 8'hDF;
            reg_file[11955] <= 8'hB3;
            reg_file[11956] <= 8'hE3;
            reg_file[11957] <= 8'h8C;
            reg_file[11958] <= 8'h05;
            reg_file[11959] <= 8'hF8;
            reg_file[11960] <= 8'h33;
            reg_file[11961] <= 8'h08;
            reg_file[11962] <= 8'hC5;
            reg_file[11963] <= 8'h40;
            reg_file[11964] <= 8'hB3;
            reg_file[11965] <= 8'h38;
            reg_file[11966] <= 8'h05;
            reg_file[11967] <= 8'h01;
            reg_file[11968] <= 8'hB3;
            reg_file[11969] <= 8'h85;
            reg_file[11970] <= 8'hE7;
            reg_file[11971] <= 8'h40;
            reg_file[11972] <= 8'hB3;
            reg_file[11973] <= 8'h85;
            reg_file[11974] <= 8'h15;
            reg_file[11975] <= 8'h41;
            reg_file[11976] <= 8'h93;
            reg_file[11977] <= 8'h98;
            reg_file[11978] <= 8'h85;
            reg_file[11979] <= 8'h00;
            reg_file[11980] <= 8'h63;
            reg_file[11981] <= 8'hDE;
            reg_file[11982] <= 8'h08;
            reg_file[11983] <= 8'h00;
            reg_file[11984] <= 8'h33;
            reg_file[11985] <= 8'h05;
            reg_file[11986] <= 8'hA6;
            reg_file[11987] <= 8'h40;
            reg_file[11988] <= 8'hB3;
            reg_file[11989] <= 8'h07;
            reg_file[11990] <= 8'hF7;
            reg_file[11991] <= 8'h40;
            reg_file[11992] <= 8'h33;
            reg_file[11993] <= 8'h36;
            reg_file[11994] <= 8'hA6;
            reg_file[11995] <= 8'h00;
            reg_file[11996] <= 8'hB3;
            reg_file[11997] <= 8'h87;
            reg_file[11998] <= 8'hC7;
            reg_file[11999] <= 8'h40;
            reg_file[12000] <= 8'h93;
            reg_file[12001] <= 8'h84;
            reg_file[12002] <= 8'h06;
            reg_file[12003] <= 8'h00;
            reg_file[12004] <= 8'h6F;
            reg_file[12005] <= 8'hF0;
            reg_file[12006] <= 8'h9F;
            reg_file[12007] <= 8'hF6;
            reg_file[12008] <= 8'h33;
            reg_file[12009] <= 8'h65;
            reg_file[12010] <= 8'hB8;
            reg_file[12011] <= 8'h00;
            reg_file[12012] <= 8'h63;
            reg_file[12013] <= 8'h1C;
            reg_file[12014] <= 8'h05;
            reg_file[12015] <= 8'h18;
            reg_file[12016] <= 8'h93;
            reg_file[12017] <= 8'h84;
            reg_file[12018] <= 8'hE9;
            reg_file[12019] <= 8'hFF;
            reg_file[12020] <= 8'h93;
            reg_file[12021] <= 8'hB4;
            reg_file[12022] <= 8'h14;
            reg_file[12023] <= 8'h00;
            reg_file[12024] <= 8'h93;
            reg_file[12025] <= 8'h07;
            reg_file[12026] <= 8'h00;
            reg_file[12027] <= 8'h00;
            reg_file[12028] <= 8'h6F;
            reg_file[12029] <= 8'hF0;
            reg_file[12030] <= 8'h1F;
            reg_file[12031] <= 8'hF5;
            reg_file[12032] <= 8'h13;
            reg_file[12033] <= 8'h0E;
            reg_file[12034] <= 8'hF0;
            reg_file[12035] <= 8'h7F;
            reg_file[12036] <= 8'h63;
            reg_file[12037] <= 8'h18;
            reg_file[12038] <= 8'hC4;
            reg_file[12039] <= 8'h03;
            reg_file[12040] <= 8'h63;
            reg_file[12041] <= 8'h08;
            reg_file[12042] <= 8'h03;
            reg_file[12043] <= 8'h2C;
            reg_file[12044] <= 8'h37;
            reg_file[12045] <= 8'h04;
            reg_file[12046] <= 8'h40;
            reg_file[12047] <= 8'h00;
            reg_file[12048] <= 8'h33;
            reg_file[12049] <= 8'hF4;
            reg_file[12050] <= 8'h87;
            reg_file[12051] <= 8'h00;
            reg_file[12052] <= 8'h13;
            reg_file[12053] <= 8'h34;
            reg_file[12054] <= 8'h14;
            reg_file[12055] <= 8'h00;
            reg_file[12056] <= 8'h13;
            reg_file[12057] <= 8'h14;
            reg_file[12058] <= 8'h44;
            reg_file[12059] <= 8'h00;
            reg_file[12060] <= 8'h63;
            reg_file[12061] <= 8'h90;
            reg_file[12062] <= 8'hC8;
            reg_file[12063] <= 8'h05;
            reg_file[12064] <= 8'h63;
            reg_file[12065] <= 8'h8E;
            reg_file[12066] <= 8'h05;
            reg_file[12067] <= 8'h00;
            reg_file[12068] <= 8'h13;
            reg_file[12069] <= 8'h18;
            reg_file[12070] <= 8'h97;
            reg_file[12071] <= 8'h00;
            reg_file[12072] <= 8'h63;
            reg_file[12073] <= 8'h4A;
            reg_file[12074] <= 8'h08;
            reg_file[12075] <= 8'h00;
            reg_file[12076] <= 8'h13;
            reg_file[12077] <= 8'h04;
            reg_file[12078] <= 8'h00;
            reg_file[12079] <= 8'h01;
            reg_file[12080] <= 8'h6F;
            reg_file[12081] <= 8'h00;
            reg_file[12082] <= 8'hC0;
            reg_file[12083] <= 8'h00;
            reg_file[12084] <= 8'h13;
            reg_file[12085] <= 8'h04;
            reg_file[12086] <= 8'h00;
            reg_file[12087] <= 8'h00;
            reg_file[12088] <= 8'hE3;
            reg_file[12089] <= 8'h84;
            reg_file[12090] <= 8'hC8;
            reg_file[12091] <= 8'hFF;
            reg_file[12092] <= 8'h63;
            reg_file[12093] <= 8'h10;
            reg_file[12094] <= 8'h03;
            reg_file[12095] <= 8'h02;
            reg_file[12096] <= 8'h63;
            reg_file[12097] <= 8'h80;
            reg_file[12098] <= 8'h05;
            reg_file[12099] <= 8'h22;
            reg_file[12100] <= 8'h93;
            reg_file[12101] <= 8'h07;
            reg_file[12102] <= 8'h07;
            reg_file[12103] <= 8'h00;
            reg_file[12104] <= 8'h13;
            reg_file[12105] <= 8'h05;
            reg_file[12106] <= 8'h06;
            reg_file[12107] <= 8'h00;
            reg_file[12108] <= 8'h93;
            reg_file[12109] <= 8'h84;
            reg_file[12110] <= 8'h06;
            reg_file[12111] <= 8'h00;
            reg_file[12112] <= 8'h6F;
            reg_file[12113] <= 8'hF0;
            reg_file[12114] <= 8'h5F;
            reg_file[12115] <= 8'hB0;
            reg_file[12116] <= 8'h13;
            reg_file[12117] <= 8'h04;
            reg_file[12118] <= 8'h00;
            reg_file[12119] <= 8'h00;
            reg_file[12120] <= 8'h6F;
            reg_file[12121] <= 8'hF0;
            reg_file[12122] <= 8'h9F;
            reg_file[12123] <= 8'hFC;
            reg_file[12124] <= 8'hE3;
            reg_file[12125] <= 8'h8C;
            reg_file[12126] <= 8'h05;
            reg_file[12127] <= 8'hAE;
            reg_file[12128] <= 8'h6F;
            reg_file[12129] <= 8'hF0;
            reg_file[12130] <= 8'h1F;
            reg_file[12131] <= 8'hB1;
            reg_file[12132] <= 8'h33;
            reg_file[12133] <= 8'h0A;
            reg_file[12134] <= 8'hC5;
            reg_file[12135] <= 8'h40;
            reg_file[12136] <= 8'hB3;
            reg_file[12137] <= 8'h35;
            reg_file[12138] <= 8'h45;
            reg_file[12139] <= 8'h01;
            reg_file[12140] <= 8'h33;
            reg_file[12141] <= 8'h89;
            reg_file[12142] <= 8'hE7;
            reg_file[12143] <= 8'h40;
            reg_file[12144] <= 8'h33;
            reg_file[12145] <= 8'h09;
            reg_file[12146] <= 8'hB9;
            reg_file[12147] <= 8'h40;
            reg_file[12148] <= 8'h93;
            reg_file[12149] <= 8'h15;
            reg_file[12150] <= 8'h89;
            reg_file[12151] <= 8'h00;
            reg_file[12152] <= 8'h63;
            reg_file[12153] <= 8'hD2;
            reg_file[12154] <= 8'h05;
            reg_file[12155] <= 8'h08;
            reg_file[12156] <= 8'h33;
            reg_file[12157] <= 8'h0A;
            reg_file[12158] <= 8'hA6;
            reg_file[12159] <= 8'h40;
            reg_file[12160] <= 8'hB3;
            reg_file[12161] <= 8'h07;
            reg_file[12162] <= 8'hF7;
            reg_file[12163] <= 8'h40;
            reg_file[12164] <= 8'h33;
            reg_file[12165] <= 8'h37;
            reg_file[12166] <= 8'h46;
            reg_file[12167] <= 8'h01;
            reg_file[12168] <= 8'h33;
            reg_file[12169] <= 8'h89;
            reg_file[12170] <= 8'hE7;
            reg_file[12171] <= 8'h40;
            reg_file[12172] <= 8'h93;
            reg_file[12173] <= 8'h84;
            reg_file[12174] <= 8'h06;
            reg_file[12175] <= 8'h00;
            reg_file[12176] <= 8'h63;
            reg_file[12177] <= 8'h0C;
            reg_file[12178] <= 8'h09;
            reg_file[12179] <= 8'h06;
            reg_file[12180] <= 8'h13;
            reg_file[12181] <= 8'h05;
            reg_file[12182] <= 8'h09;
            reg_file[12183] <= 8'h00;
            reg_file[12184] <= 8'hEF;
            reg_file[12185] <= 8'h00;
            reg_file[12186] <= 8'h80;
            reg_file[12187] <= 8'h25;
            reg_file[12188] <= 8'h13;
            reg_file[12189] <= 8'h08;
            reg_file[12190] <= 8'h85;
            reg_file[12191] <= 8'hFF;
            reg_file[12192] <= 8'h93;
            reg_file[12193] <= 8'h07;
            reg_file[12194] <= 8'hF0;
            reg_file[12195] <= 8'h01;
            reg_file[12196] <= 8'h63;
            reg_file[12197] <= 8'hCA;
            reg_file[12198] <= 8'h07;
            reg_file[12199] <= 8'h07;
            reg_file[12200] <= 8'h93;
            reg_file[12201] <= 8'h07;
            reg_file[12202] <= 8'h00;
            reg_file[12203] <= 8'h02;
            reg_file[12204] <= 8'hB3;
            reg_file[12205] <= 8'h87;
            reg_file[12206] <= 8'h07;
            reg_file[12207] <= 8'h41;
            reg_file[12208] <= 8'h33;
            reg_file[12209] <= 8'h17;
            reg_file[12210] <= 8'h09;
            reg_file[12211] <= 8'h01;
            reg_file[12212] <= 8'hB3;
            reg_file[12213] <= 8'h57;
            reg_file[12214] <= 8'hFA;
            reg_file[12215] <= 8'h00;
            reg_file[12216] <= 8'hB3;
            reg_file[12217] <= 8'hE7;
            reg_file[12218] <= 8'hE7;
            reg_file[12219] <= 8'h00;
            reg_file[12220] <= 8'h33;
            reg_file[12221] <= 8'h16;
            reg_file[12222] <= 8'h0A;
            reg_file[12223] <= 8'h01;
            reg_file[12224] <= 8'h63;
            reg_file[12225] <= 8'h4C;
            reg_file[12226] <= 8'h88;
            reg_file[12227] <= 8'h08;
            reg_file[12228] <= 8'h33;
            reg_file[12229] <= 8'h08;
            reg_file[12230] <= 8'h88;
            reg_file[12231] <= 8'h40;
            reg_file[12232] <= 8'h93;
            reg_file[12233] <= 8'h05;
            reg_file[12234] <= 8'h18;
            reg_file[12235] <= 8'h00;
            reg_file[12236] <= 8'h13;
            reg_file[12237] <= 8'h07;
            reg_file[12238] <= 8'hF0;
            reg_file[12239] <= 8'h01;
            reg_file[12240] <= 8'h63;
            reg_file[12241] <= 8'h4C;
            reg_file[12242] <= 8'hB7;
            reg_file[12243] <= 8'h04;
            reg_file[12244] <= 8'h93;
            reg_file[12245] <= 8'h06;
            reg_file[12246] <= 8'h00;
            reg_file[12247] <= 8'h02;
            reg_file[12248] <= 8'hB3;
            reg_file[12249] <= 8'h86;
            reg_file[12250] <= 8'hB6;
            reg_file[12251] <= 8'h40;
            reg_file[12252] <= 8'h33;
            reg_file[12253] <= 8'h95;
            reg_file[12254] <= 8'hD7;
            reg_file[12255] <= 8'h00;
            reg_file[12256] <= 8'h33;
            reg_file[12257] <= 8'h57;
            reg_file[12258] <= 8'hB6;
            reg_file[12259] <= 8'h00;
            reg_file[12260] <= 8'h33;
            reg_file[12261] <= 8'h16;
            reg_file[12262] <= 8'hD6;
            reg_file[12263] <= 8'h00;
            reg_file[12264] <= 8'h33;
            reg_file[12265] <= 8'h65;
            reg_file[12266] <= 8'hE5;
            reg_file[12267] <= 8'h00;
            reg_file[12268] <= 8'h33;
            reg_file[12269] <= 8'h36;
            reg_file[12270] <= 8'hC0;
            reg_file[12271] <= 8'h00;
            reg_file[12272] <= 8'h33;
            reg_file[12273] <= 8'h65;
            reg_file[12274] <= 8'hC5;
            reg_file[12275] <= 8'h00;
            reg_file[12276] <= 8'hB3;
            reg_file[12277] <= 8'hD7;
            reg_file[12278] <= 8'hB7;
            reg_file[12279] <= 8'h00;
            reg_file[12280] <= 8'h6F;
            reg_file[12281] <= 8'hF0;
            reg_file[12282] <= 8'h5F;
            reg_file[12283] <= 8'hE5;
            reg_file[12284] <= 8'h33;
            reg_file[12285] <= 8'h65;
            reg_file[12286] <= 8'h2A;
            reg_file[12287] <= 8'h01;
            reg_file[12288] <= 8'hE3;
            reg_file[12289] <= 8'h18;
            reg_file[12290] <= 8'h05;
            reg_file[12291] <= 8'hF8;
            reg_file[12292] <= 8'h6F;
            reg_file[12293] <= 8'hF0;
            reg_file[12294] <= 8'hDF;
            reg_file[12295] <= 8'hEE;
            reg_file[12296] <= 8'h13;
            reg_file[12297] <= 8'h05;
            reg_file[12298] <= 8'h0A;
            reg_file[12299] <= 8'h00;
            reg_file[12300] <= 8'hEF;
            reg_file[12301] <= 8'h00;
            reg_file[12302] <= 8'h40;
            reg_file[12303] <= 8'h1E;
            reg_file[12304] <= 8'h13;
            reg_file[12305] <= 8'h05;
            reg_file[12306] <= 8'h05;
            reg_file[12307] <= 8'h02;
            reg_file[12308] <= 8'h6F;
            reg_file[12309] <= 8'hF0;
            reg_file[12310] <= 8'h9F;
            reg_file[12311] <= 8'hF8;
            reg_file[12312] <= 8'h93;
            reg_file[12313] <= 8'h07;
            reg_file[12314] <= 8'h85;
            reg_file[12315] <= 8'hFD;
            reg_file[12316] <= 8'hB3;
            reg_file[12317] <= 8'h17;
            reg_file[12318] <= 8'hFA;
            reg_file[12319] <= 8'h00;
            reg_file[12320] <= 8'h13;
            reg_file[12321] <= 8'h06;
            reg_file[12322] <= 8'h00;
            reg_file[12323] <= 8'h00;
            reg_file[12324] <= 8'h6F;
            reg_file[12325] <= 8'hF0;
            reg_file[12326] <= 8'hDF;
            reg_file[12327] <= 8'hF9;
            reg_file[12328] <= 8'h13;
            reg_file[12329] <= 8'h08;
            reg_file[12330] <= 8'h18;
            reg_file[12331] <= 8'hFE;
            reg_file[12332] <= 8'h93;
            reg_file[12333] <= 8'h06;
            reg_file[12334] <= 8'h00;
            reg_file[12335] <= 8'h02;
            reg_file[12336] <= 8'h33;
            reg_file[12337] <= 8'hD8;
            reg_file[12338] <= 8'h07;
            reg_file[12339] <= 8'h01;
            reg_file[12340] <= 8'h13;
            reg_file[12341] <= 8'h07;
            reg_file[12342] <= 8'h00;
            reg_file[12343] <= 8'h00;
            reg_file[12344] <= 8'h63;
            reg_file[12345] <= 8'h88;
            reg_file[12346] <= 8'hD5;
            reg_file[12347] <= 8'h00;
            reg_file[12348] <= 8'h13;
            reg_file[12349] <= 8'h07;
            reg_file[12350] <= 8'h00;
            reg_file[12351] <= 8'h04;
            reg_file[12352] <= 8'h33;
            reg_file[12353] <= 8'h07;
            reg_file[12354] <= 8'hB7;
            reg_file[12355] <= 8'h40;
            reg_file[12356] <= 8'h33;
            reg_file[12357] <= 8'h97;
            reg_file[12358] <= 8'hE7;
            reg_file[12359] <= 8'h00;
            reg_file[12360] <= 8'h33;
            reg_file[12361] <= 8'h67;
            reg_file[12362] <= 8'hE6;
            reg_file[12363] <= 8'h00;
            reg_file[12364] <= 8'h33;
            reg_file[12365] <= 8'h35;
            reg_file[12366] <= 8'hE0;
            reg_file[12367] <= 8'h00;
            reg_file[12368] <= 8'h33;
            reg_file[12369] <= 8'h65;
            reg_file[12370] <= 8'hA8;
            reg_file[12371] <= 8'h00;
            reg_file[12372] <= 8'h6F;
            reg_file[12373] <= 8'hF0;
            reg_file[12374] <= 8'h5F;
            reg_file[12375] <= 8'hEA;
            reg_file[12376] <= 8'h37;
            reg_file[12377] <= 8'h07;
            reg_file[12378] <= 8'h80;
            reg_file[12379] <= 8'hFF;
            reg_file[12380] <= 8'h13;
            reg_file[12381] <= 8'h05;
            reg_file[12382] <= 8'hF7;
            reg_file[12383] <= 8'hFF;
            reg_file[12384] <= 8'h33;
            reg_file[12385] <= 8'h08;
            reg_file[12386] <= 8'h04;
            reg_file[12387] <= 8'h41;
            reg_file[12388] <= 8'h33;
            reg_file[12389] <= 8'hF7;
            reg_file[12390] <= 8'hA7;
            reg_file[12391] <= 8'h00;
            reg_file[12392] <= 8'h6F;
            reg_file[12393] <= 8'hF0;
            reg_file[12394] <= 8'h5F;
            reg_file[12395] <= 8'h81;
            reg_file[12396] <= 8'h93;
            reg_file[12397] <= 8'h07;
            reg_file[12398] <= 8'h07;
            reg_file[12399] <= 8'h00;
            reg_file[12400] <= 8'h13;
            reg_file[12401] <= 8'h05;
            reg_file[12402] <= 8'h06;
            reg_file[12403] <= 8'h00;
            reg_file[12404] <= 8'h6F;
            reg_file[12405] <= 8'hF0;
            reg_file[12406] <= 8'h9F;
            reg_file[12407] <= 8'hDD;
            reg_file[12408] <= 8'h93;
            reg_file[12409] <= 8'h07;
            reg_file[12410] <= 8'h07;
            reg_file[12411] <= 8'h00;
            reg_file[12412] <= 8'h13;
            reg_file[12413] <= 8'h05;
            reg_file[12414] <= 8'h06;
            reg_file[12415] <= 8'h00;
            reg_file[12416] <= 8'h6F;
            reg_file[12417] <= 8'hF0;
            reg_file[12418] <= 8'h1F;
            reg_file[12419] <= 8'hE6;
            reg_file[12420] <= 8'h93;
            reg_file[12421] <= 8'h87;
            reg_file[12422] <= 8'h05;
            reg_file[12423] <= 8'h00;
            reg_file[12424] <= 8'h13;
            reg_file[12425] <= 8'h05;
            reg_file[12426] <= 8'h08;
            reg_file[12427] <= 8'h00;
            reg_file[12428] <= 8'h6F;
            reg_file[12429] <= 8'hF0;
            reg_file[12430] <= 8'h1F;
            reg_file[12431] <= 8'hDC;
            reg_file[12432] <= 8'h13;
            reg_file[12433] <= 8'h84;
            reg_file[12434] <= 8'h04;
            reg_file[12435] <= 8'h00;
            reg_file[12436] <= 8'hE3;
            reg_file[12437] <= 8'h96;
            reg_file[12438] <= 8'h04;
            reg_file[12439] <= 8'hE0;
            reg_file[12440] <= 8'h13;
            reg_file[12441] <= 8'h37;
            reg_file[12442] <= 8'h87;
            reg_file[12443] <= 8'hFF;
            reg_file[12444] <= 8'h13;
            reg_file[12445] <= 8'h47;
            reg_file[12446] <= 8'h17;
            reg_file[12447] <= 8'h00;
            reg_file[12448] <= 8'hB3;
            reg_file[12449] <= 8'h88;
            reg_file[12450] <= 8'hE8;
            reg_file[12451] <= 8'h00;
            reg_file[12452] <= 8'h13;
            reg_file[12453] <= 8'h04;
            reg_file[12454] <= 8'h10;
            reg_file[12455] <= 8'h00;
            reg_file[12456] <= 8'h6F;
            reg_file[12457] <= 8'hF0;
            reg_file[12458] <= 8'h9F;
            reg_file[12459] <= 8'hDF;
            reg_file[12460] <= 8'h13;
            reg_file[12461] <= 8'h04;
            reg_file[12462] <= 8'h10;
            reg_file[12463] <= 8'h00;
            reg_file[12464] <= 8'hE3;
            reg_file[12465] <= 8'h88;
            reg_file[12466] <= 8'h04;
            reg_file[12467] <= 8'hDE;
            reg_file[12468] <= 8'h13;
            reg_file[12469] <= 8'h37;
            reg_file[12470] <= 8'h87;
            reg_file[12471] <= 8'hFF;
            reg_file[12472] <= 8'h13;
            reg_file[12473] <= 8'h47;
            reg_file[12474] <= 8'h17;
            reg_file[12475] <= 8'h00;
            reg_file[12476] <= 8'hB3;
            reg_file[12477] <= 8'h88;
            reg_file[12478] <= 8'hE8;
            reg_file[12479] <= 8'h00;
            reg_file[12480] <= 8'h13;
            reg_file[12481] <= 8'h84;
            reg_file[12482] <= 8'h04;
            reg_file[12483] <= 8'h00;
            reg_file[12484] <= 8'h6F;
            reg_file[12485] <= 8'hF0;
            reg_file[12486] <= 8'hDF;
            reg_file[12487] <= 8'hDD;
            reg_file[12488] <= 8'h93;
            reg_file[12489] <= 8'h07;
            reg_file[12490] <= 8'h00;
            reg_file[12491] <= 8'h00;
            reg_file[12492] <= 8'h13;
            reg_file[12493] <= 8'h08;
            reg_file[12494] <= 8'hF0;
            reg_file[12495] <= 8'h7F;
            reg_file[12496] <= 8'h6F;
            reg_file[12497] <= 8'hF0;
            reg_file[12498] <= 8'h8F;
            reg_file[12499] <= 8'hE9;
            reg_file[12500] <= 8'h93;
            reg_file[12501] <= 8'h07;
            reg_file[12502] <= 8'h07;
            reg_file[12503] <= 8'h00;
            reg_file[12504] <= 8'h13;
            reg_file[12505] <= 8'h05;
            reg_file[12506] <= 8'h06;
            reg_file[12507] <= 8'h00;
            reg_file[12508] <= 8'h13;
            reg_file[12509] <= 8'h08;
            reg_file[12510] <= 8'hF0;
            reg_file[12511] <= 8'h7F;
            reg_file[12512] <= 8'h6F;
            reg_file[12513] <= 8'hF0;
            reg_file[12514] <= 8'h5F;
            reg_file[12515] <= 8'hA6;
            reg_file[12516] <= 8'h93;
            reg_file[12517] <= 8'h07;
            reg_file[12518] <= 8'hF0;
            reg_file[12519] <= 8'hFF;
            reg_file[12520] <= 8'h13;
            reg_file[12521] <= 8'h05;
            reg_file[12522] <= 8'hF0;
            reg_file[12523] <= 8'hFF;
            reg_file[12524] <= 8'h13;
            reg_file[12525] <= 8'h08;
            reg_file[12526] <= 8'hE0;
            reg_file[12527] <= 8'h7F;
            reg_file[12528] <= 8'h93;
            reg_file[12529] <= 8'h08;
            reg_file[12530] <= 8'h00;
            reg_file[12531] <= 8'h00;
            reg_file[12532] <= 8'h6F;
            reg_file[12533] <= 8'hF0;
            reg_file[12534] <= 8'h1F;
            reg_file[12535] <= 8'hA9;
            reg_file[12536] <= 8'h93;
            reg_file[12537] <= 8'h07;
            reg_file[12538] <= 8'h00;
            reg_file[12539] <= 8'h00;
            reg_file[12540] <= 8'h13;
            reg_file[12541] <= 8'h05;
            reg_file[12542] <= 8'h00;
            reg_file[12543] <= 8'h00;
            reg_file[12544] <= 8'h6F;
            reg_file[12545] <= 8'hF0;
            reg_file[12546] <= 8'h1F;
            reg_file[12547] <= 8'h98;
            reg_file[12548] <= 8'h93;
            reg_file[12549] <= 8'h07;
            reg_file[12550] <= 8'h00;
            reg_file[12551] <= 8'h00;
            reg_file[12552] <= 8'h13;
            reg_file[12553] <= 8'h05;
            reg_file[12554] <= 8'h00;
            reg_file[12555] <= 8'h00;
            reg_file[12556] <= 8'h6F;
            reg_file[12557] <= 8'hF0;
            reg_file[12558] <= 8'h1F;
            reg_file[12559] <= 8'hFC;
            reg_file[12560] <= 8'h93;
            reg_file[12561] <= 8'h07;
            reg_file[12562] <= 8'h07;
            reg_file[12563] <= 8'h00;
            reg_file[12564] <= 8'h13;
            reg_file[12565] <= 8'h05;
            reg_file[12566] <= 8'h06;
            reg_file[12567] <= 8'h00;
            reg_file[12568] <= 8'h93;
            reg_file[12569] <= 8'h08;
            reg_file[12570] <= 8'h00;
            reg_file[12571] <= 8'h00;
            reg_file[12572] <= 8'h6F;
            reg_file[12573] <= 8'hF0;
            reg_file[12574] <= 8'h1F;
            reg_file[12575] <= 8'h8D;
            reg_file[12576] <= 8'h93;
            reg_file[12577] <= 8'h07;
            reg_file[12578] <= 8'h00;
            reg_file[12579] <= 8'h00;
            reg_file[12580] <= 8'h93;
            reg_file[12581] <= 8'h84;
            reg_file[12582] <= 8'h06;
            reg_file[12583] <= 8'h00;
            reg_file[12584] <= 8'h6F;
            reg_file[12585] <= 8'hF0;
            reg_file[12586] <= 8'h9F;
            reg_file[12587] <= 8'h95;
            reg_file[12588] <= 8'h93;
            reg_file[12589] <= 8'h07;
            reg_file[12590] <= 8'h07;
            reg_file[12591] <= 8'h00;
            reg_file[12592] <= 8'h13;
            reg_file[12593] <= 8'h05;
            reg_file[12594] <= 8'h06;
            reg_file[12595] <= 8'h00;
            reg_file[12596] <= 8'h93;
            reg_file[12597] <= 8'h84;
            reg_file[12598] <= 8'h06;
            reg_file[12599] <= 8'h00;
            reg_file[12600] <= 8'h6F;
            reg_file[12601] <= 8'hF0;
            reg_file[12602] <= 8'h1F;
            reg_file[12603] <= 8'hFE;
            reg_file[12604] <= 8'h93;
            reg_file[12605] <= 8'h07;
            reg_file[12606] <= 8'h00;
            reg_file[12607] <= 8'h00;
            reg_file[12608] <= 8'h13;
            reg_file[12609] <= 8'h08;
            reg_file[12610] <= 8'hF0;
            reg_file[12611] <= 8'h7F;
            reg_file[12612] <= 8'h93;
            reg_file[12613] <= 8'h84;
            reg_file[12614] <= 8'h06;
            reg_file[12615] <= 8'h00;
            reg_file[12616] <= 8'h6F;
            reg_file[12617] <= 8'hF0;
            reg_file[12618] <= 8'h0F;
            reg_file[12619] <= 8'hE2;
            reg_file[12620] <= 8'h93;
            reg_file[12621] <= 8'h07;
            reg_file[12622] <= 8'h07;
            reg_file[12623] <= 8'h00;
            reg_file[12624] <= 8'h13;
            reg_file[12625] <= 8'h05;
            reg_file[12626] <= 8'h06;
            reg_file[12627] <= 8'h00;
            reg_file[12628] <= 8'h13;
            reg_file[12629] <= 8'h08;
            reg_file[12630] <= 8'hF0;
            reg_file[12631] <= 8'h7F;
            reg_file[12632] <= 8'h93;
            reg_file[12633] <= 8'h84;
            reg_file[12634] <= 8'h06;
            reg_file[12635] <= 8'h00;
            reg_file[12636] <= 8'h6F;
            reg_file[12637] <= 8'hF0;
            reg_file[12638] <= 8'h9F;
            reg_file[12639] <= 8'h9E;
            reg_file[12640] <= 8'h13;
            reg_file[12641] <= 8'h05;
            reg_file[12642] <= 8'h00;
            reg_file[12643] <= 8'h00;
            reg_file[12644] <= 8'h93;
            reg_file[12645] <= 8'h04;
            reg_file[12646] <= 8'h00;
            reg_file[12647] <= 8'h00;
            reg_file[12648] <= 8'hB7;
            reg_file[12649] <= 8'h07;
            reg_file[12650] <= 8'h40;
            reg_file[12651] <= 8'h00;
            reg_file[12652] <= 8'h13;
            reg_file[12653] <= 8'h08;
            reg_file[12654] <= 8'hF0;
            reg_file[12655] <= 8'h7F;
            reg_file[12656] <= 8'h13;
            reg_file[12657] <= 8'h04;
            reg_file[12658] <= 8'h00;
            reg_file[12659] <= 8'h01;
            reg_file[12660] <= 8'h6F;
            reg_file[12661] <= 8'hF0;
            reg_file[12662] <= 8'hDF;
            reg_file[12663] <= 8'h90;
            reg_file[12664] <= 8'h93;
            reg_file[12665] <= 8'h07;
            reg_file[12666] <= 8'h00;
            reg_file[12667] <= 8'h00;
            reg_file[12668] <= 8'h13;
            reg_file[12669] <= 8'h05;
            reg_file[12670] <= 8'h00;
            reg_file[12671] <= 8'h00;
            reg_file[12672] <= 8'h13;
            reg_file[12673] <= 8'h08;
            reg_file[12674] <= 8'h00;
            reg_file[12675] <= 8'h00;
            reg_file[12676] <= 8'h6F;
            reg_file[12677] <= 8'hF0;
            reg_file[12678] <= 8'h4F;
            reg_file[12679] <= 8'hDE;
            reg_file[12680] <= 8'h63;
            reg_file[12681] <= 8'h98;
            reg_file[12682] <= 8'h04;
            reg_file[12683] <= 8'h00;
            reg_file[12684] <= 8'h13;
            reg_file[12685] <= 8'h07;
            reg_file[12686] <= 8'h85;
            reg_file[12687] <= 8'h00;
            reg_file[12688] <= 8'h6F;
            reg_file[12689] <= 8'hF0;
            reg_file[12690] <= 8'h1F;
            reg_file[12691] <= 8'hA2;
            reg_file[12692] <= 8'hE3;
            reg_file[12693] <= 8'h9C;
            reg_file[12694] <= 8'h04;
            reg_file[12695] <= 8'hFE;
            reg_file[12696] <= 8'hE3;
            reg_file[12697] <= 8'h94;
            reg_file[12698] <= 8'h08;
            reg_file[12699] <= 8'h86;
            reg_file[12700] <= 8'h6F;
            reg_file[12701] <= 8'hF0;
            reg_file[12702] <= 8'h5F;
            reg_file[12703] <= 8'h8E;
            reg_file[12704] <= 8'h13;
            reg_file[12705] <= 8'h05;
            reg_file[12706] <= 8'h00;
            reg_file[12707] <= 8'h00;
            reg_file[12708] <= 8'h63;
            reg_file[12709] <= 8'h84;
            reg_file[12710] <= 8'h09;
            reg_file[12711] <= 8'h02;
            reg_file[12712] <= 8'h93;
            reg_file[12713] <= 8'h07;
            reg_file[12714] <= 8'h30;
            reg_file[12715] <= 8'h00;
            reg_file[12716] <= 8'h63;
            reg_file[12717] <= 8'h9A;
            reg_file[12718] <= 8'hF9;
            reg_file[12719] <= 8'h00;
            reg_file[12720] <= 8'h63;
            reg_file[12721] <= 8'h8E;
            reg_file[12722] <= 8'h04;
            reg_file[12723] <= 8'h00;
            reg_file[12724] <= 8'h13;
            reg_file[12725] <= 8'h05;
            reg_file[12726] <= 8'hF0;
            reg_file[12727] <= 8'hFF;
            reg_file[12728] <= 8'h13;
            reg_file[12729] <= 8'h08;
            reg_file[12730] <= 8'hE0;
            reg_file[12731] <= 8'h7F;
            reg_file[12732] <= 8'h6F;
            reg_file[12733] <= 8'h00;
            reg_file[12734] <= 8'h00;
            reg_file[12735] <= 8'h01;
            reg_file[12736] <= 8'h93;
            reg_file[12737] <= 8'h07;
            reg_file[12738] <= 8'h20;
            reg_file[12739] <= 8'h00;
            reg_file[12740] <= 8'hE3;
            reg_file[12741] <= 8'h98;
            reg_file[12742] <= 8'hF9;
            reg_file[12743] <= 8'hFE;
            reg_file[12744] <= 8'hE3;
            reg_file[12745] <= 8'h86;
            reg_file[12746] <= 8'h04;
            reg_file[12747] <= 8'hFE;
            reg_file[12748] <= 8'h13;
            reg_file[12749] <= 8'h64;
            reg_file[12750] <= 8'h54;
            reg_file[12751] <= 8'h00;
            reg_file[12752] <= 8'h93;
            reg_file[12753] <= 8'h07;
            reg_file[12754] <= 8'h05;
            reg_file[12755] <= 8'h00;
            reg_file[12756] <= 8'h6F;
            reg_file[12757] <= 8'hF0;
            reg_file[12758] <= 8'hDF;
            reg_file[12759] <= 8'h8C;
            reg_file[12760] <= 8'hE3;
            reg_file[12761] <= 8'h8E;
            reg_file[12762] <= 8'h88;
            reg_file[12763] <= 8'hD6;
            reg_file[12764] <= 8'h13;
            reg_file[12765] <= 8'h04;
            reg_file[12766] <= 8'h00;
            reg_file[12767] <= 8'h00;
            reg_file[12768] <= 8'h6F;
            reg_file[12769] <= 8'hF0;
            reg_file[12770] <= 8'h1F;
            reg_file[12771] <= 8'hD6;
            reg_file[12772] <= 8'hE3;
            reg_file[12773] <= 8'h8E;
            reg_file[12774] <= 8'h88;
            reg_file[12775] <= 8'h86;
            reg_file[12776] <= 8'h13;
            reg_file[12777] <= 8'h04;
            reg_file[12778] <= 8'h00;
            reg_file[12779] <= 8'h00;
            reg_file[12780] <= 8'h6F;
            reg_file[12781] <= 8'hF0;
            reg_file[12782] <= 8'h1F;
            reg_file[12783] <= 8'h86;
            reg_file[12784] <= 8'hB7;
            reg_file[12785] <= 8'h07;
            reg_file[12786] <= 8'h01;
            reg_file[12787] <= 8'h00;
            reg_file[12788] <= 8'h63;
            reg_file[12789] <= 8'h7A;
            reg_file[12790] <= 8'hF5;
            reg_file[12791] <= 8'h02;
            reg_file[12792] <= 8'h93;
            reg_file[12793] <= 8'h07;
            reg_file[12794] <= 8'hF0;
            reg_file[12795] <= 8'h0F;
            reg_file[12796] <= 8'hB3;
            reg_file[12797] <= 8'hB7;
            reg_file[12798] <= 8'hA7;
            reg_file[12799] <= 8'h00;
            reg_file[12800] <= 8'h93;
            reg_file[12801] <= 8'h97;
            reg_file[12802] <= 8'h37;
            reg_file[12803] <= 8'h00;
            reg_file[12804] <= 8'h37;
            reg_file[12805] <= 8'h37;
            reg_file[12806] <= 8'h00;
            reg_file[12807] <= 8'h80;
            reg_file[12808] <= 8'h93;
            reg_file[12809] <= 8'h06;
            reg_file[12810] <= 8'h00;
            reg_file[12811] <= 8'h02;
            reg_file[12812] <= 8'hB3;
            reg_file[12813] <= 8'h86;
            reg_file[12814] <= 8'hF6;
            reg_file[12815] <= 8'h40;
            reg_file[12816] <= 8'h33;
            reg_file[12817] <= 8'h55;
            reg_file[12818] <= 8'hF5;
            reg_file[12819] <= 8'h00;
            reg_file[12820] <= 8'h93;
            reg_file[12821] <= 8'h07;
            reg_file[12822] <= 8'h47;
            reg_file[12823] <= 8'h6B;
            reg_file[12824] <= 8'h33;
            reg_file[12825] <= 8'h85;
            reg_file[12826] <= 8'hA7;
            reg_file[12827] <= 8'h00;
            reg_file[12828] <= 8'h03;
            reg_file[12829] <= 8'h45;
            reg_file[12830] <= 8'h05;
            reg_file[12831] <= 8'h00;
            reg_file[12832] <= 8'h33;
            reg_file[12833] <= 8'h85;
            reg_file[12834] <= 8'hA6;
            reg_file[12835] <= 8'h40;
            reg_file[12836] <= 8'h67;
            reg_file[12837] <= 8'h80;
            reg_file[12838] <= 8'h00;
            reg_file[12839] <= 8'h00;
            reg_file[12840] <= 8'h37;
            reg_file[12841] <= 8'h07;
            reg_file[12842] <= 8'h00;
            reg_file[12843] <= 8'h01;
            reg_file[12844] <= 8'h93;
            reg_file[12845] <= 8'h07;
            reg_file[12846] <= 8'h00;
            reg_file[12847] <= 8'h01;
            reg_file[12848] <= 8'hE3;
            reg_file[12849] <= 8'h6A;
            reg_file[12850] <= 8'hE5;
            reg_file[12851] <= 8'hFC;
            reg_file[12852] <= 8'h93;
            reg_file[12853] <= 8'h07;
            reg_file[12854] <= 8'h80;
            reg_file[12855] <= 8'h01;
            reg_file[12856] <= 8'h6F;
            reg_file[12857] <= 8'hF0;
            reg_file[12858] <= 8'hDF;
            reg_file[12859] <= 8'hFC;
            reg_file[12860] <= 8'h93;
            reg_file[12861] <= 8'h05;
            reg_file[12862] <= 8'h05;
            reg_file[12863] <= 8'h00;
            reg_file[12864] <= 8'h93;
            reg_file[12865] <= 8'h06;
            reg_file[12866] <= 8'h00;
            reg_file[12867] <= 8'h00;
            reg_file[12868] <= 8'h13;
            reg_file[12869] <= 8'h06;
            reg_file[12870] <= 8'h00;
            reg_file[12871] <= 8'h00;
            reg_file[12872] <= 8'h13;
            reg_file[12873] <= 8'h05;
            reg_file[12874] <= 8'h00;
            reg_file[12875] <= 8'h00;
            reg_file[12876] <= 8'h6F;
            reg_file[12877] <= 8'h00;
            reg_file[12878] <= 8'h00;
            reg_file[12879] <= 8'h23;
            reg_file[12880] <= 8'h13;
            reg_file[12881] <= 8'h01;
            reg_file[12882] <= 8'h01;
            reg_file[12883] <= 8'hFF;
            reg_file[12884] <= 8'h93;
            reg_file[12885] <= 8'h05;
            reg_file[12886] <= 8'h00;
            reg_file[12887] <= 8'h00;
            reg_file[12888] <= 8'h23;
            reg_file[12889] <= 8'h24;
            reg_file[12890] <= 8'h81;
            reg_file[12891] <= 8'h00;
            reg_file[12892] <= 8'h23;
            reg_file[12893] <= 8'h26;
            reg_file[12894] <= 8'h11;
            reg_file[12895] <= 8'h00;
            reg_file[12896] <= 8'h13;
            reg_file[12897] <= 8'h04;
            reg_file[12898] <= 8'h05;
            reg_file[12899] <= 8'h00;
            reg_file[12900] <= 8'hEF;
            reg_file[12901] <= 8'h00;
            reg_file[12902] <= 8'h40;
            reg_file[12903] <= 8'h2B;
            reg_file[12904] <= 8'hB7;
            reg_file[12905] <= 8'h57;
            reg_file[12906] <= 8'h00;
            reg_file[12907] <= 8'h80;
            reg_file[12908] <= 8'h03;
            reg_file[12909] <= 8'hA5;
            reg_file[12910] <= 8'h07;
            reg_file[12911] <= 8'hCF;
            reg_file[12912] <= 8'h83;
            reg_file[12913] <= 8'h27;
            reg_file[12914] <= 8'hC5;
            reg_file[12915] <= 8'h03;
            reg_file[12916] <= 8'h63;
            reg_file[12917] <= 8'h84;
            reg_file[12918] <= 8'h07;
            reg_file[12919] <= 8'h00;
            reg_file[12920] <= 8'hE7;
            reg_file[12921] <= 8'h80;
            reg_file[12922] <= 8'h07;
            reg_file[12923] <= 8'h00;
            reg_file[12924] <= 8'h13;
            reg_file[12925] <= 8'h05;
            reg_file[12926] <= 8'h04;
            reg_file[12927] <= 8'h00;
            reg_file[12928] <= 8'hEF;
            reg_file[12929] <= 8'hC0;
            reg_file[12930] <= 8'hDF;
            reg_file[12931] <= 8'hF3;
            reg_file[12932] <= 8'hB3;
            reg_file[12933] <= 8'hC7;
            reg_file[12934] <= 8'hA5;
            reg_file[12935] <= 8'h00;
            reg_file[12936] <= 8'h93;
            reg_file[12937] <= 8'hF7;
            reg_file[12938] <= 8'h37;
            reg_file[12939] <= 8'h00;
            reg_file[12940] <= 8'hB3;
            reg_file[12941] <= 8'h08;
            reg_file[12942] <= 8'hC5;
            reg_file[12943] <= 8'h00;
            reg_file[12944] <= 8'h63;
            reg_file[12945] <= 8'h92;
            reg_file[12946] <= 8'h07;
            reg_file[12947] <= 8'h06;
            reg_file[12948] <= 8'h93;
            reg_file[12949] <= 8'h07;
            reg_file[12950] <= 8'h30;
            reg_file[12951] <= 8'h00;
            reg_file[12952] <= 8'h63;
            reg_file[12953] <= 8'hFE;
            reg_file[12954] <= 8'hC7;
            reg_file[12955] <= 8'h04;
            reg_file[12956] <= 8'h93;
            reg_file[12957] <= 8'h77;
            reg_file[12958] <= 8'h35;
            reg_file[12959] <= 8'h00;
            reg_file[12960] <= 8'h13;
            reg_file[12961] <= 8'h07;
            reg_file[12962] <= 8'h05;
            reg_file[12963] <= 8'h00;
            reg_file[12964] <= 8'h63;
            reg_file[12965] <= 8'h98;
            reg_file[12966] <= 8'h07;
            reg_file[12967] <= 8'h06;
            reg_file[12968] <= 8'h13;
            reg_file[12969] <= 8'hF6;
            reg_file[12970] <= 8'hC8;
            reg_file[12971] <= 8'hFF;
            reg_file[12972] <= 8'h93;
            reg_file[12973] <= 8'h07;
            reg_file[12974] <= 8'h06;
            reg_file[12975] <= 8'hFE;
            reg_file[12976] <= 8'h63;
            reg_file[12977] <= 8'h6C;
            reg_file[12978] <= 8'hF7;
            reg_file[12979] <= 8'h08;
            reg_file[12980] <= 8'h63;
            reg_file[12981] <= 8'h7C;
            reg_file[12982] <= 8'hC7;
            reg_file[12983] <= 8'h02;
            reg_file[12984] <= 8'h93;
            reg_file[12985] <= 8'h86;
            reg_file[12986] <= 8'h05;
            reg_file[12987] <= 8'h00;
            reg_file[12988] <= 8'h93;
            reg_file[12989] <= 8'h07;
            reg_file[12990] <= 8'h07;
            reg_file[12991] <= 8'h00;
            reg_file[12992] <= 8'h03;
            reg_file[12993] <= 8'hA8;
            reg_file[12994] <= 8'h06;
            reg_file[12995] <= 8'h00;
            reg_file[12996] <= 8'h93;
            reg_file[12997] <= 8'h87;
            reg_file[12998] <= 8'h47;
            reg_file[12999] <= 8'h00;
            reg_file[13000] <= 8'h93;
            reg_file[13001] <= 8'h86;
            reg_file[13002] <= 8'h46;
            reg_file[13003] <= 8'h00;
            reg_file[13004] <= 8'h23;
            reg_file[13005] <= 8'hAE;
            reg_file[13006] <= 8'h07;
            reg_file[13007] <= 8'hFF;
            reg_file[13008] <= 8'hE3;
            reg_file[13009] <= 8'hE8;
            reg_file[13010] <= 8'hC7;
            reg_file[13011] <= 8'hFE;
            reg_file[13012] <= 8'h93;
            reg_file[13013] <= 8'h07;
            reg_file[13014] <= 8'hF6;
            reg_file[13015] <= 8'hFF;
            reg_file[13016] <= 8'hB3;
            reg_file[13017] <= 8'h87;
            reg_file[13018] <= 8'hE7;
            reg_file[13019] <= 8'h40;
            reg_file[13020] <= 8'h93;
            reg_file[13021] <= 8'hF7;
            reg_file[13022] <= 8'hC7;
            reg_file[13023] <= 8'hFF;
            reg_file[13024] <= 8'h93;
            reg_file[13025] <= 8'h87;
            reg_file[13026] <= 8'h47;
            reg_file[13027] <= 8'h00;
            reg_file[13028] <= 8'h33;
            reg_file[13029] <= 8'h07;
            reg_file[13030] <= 8'hF7;
            reg_file[13031] <= 8'h00;
            reg_file[13032] <= 8'hB3;
            reg_file[13033] <= 8'h85;
            reg_file[13034] <= 8'hF5;
            reg_file[13035] <= 8'h00;
            reg_file[13036] <= 8'h63;
            reg_file[13037] <= 8'h68;
            reg_file[13038] <= 8'h17;
            reg_file[13039] <= 8'h01;
            reg_file[13040] <= 8'h67;
            reg_file[13041] <= 8'h80;
            reg_file[13042] <= 8'h00;
            reg_file[13043] <= 8'h00;
            reg_file[13044] <= 8'h13;
            reg_file[13045] <= 8'h07;
            reg_file[13046] <= 8'h05;
            reg_file[13047] <= 8'h00;
            reg_file[13048] <= 8'hE3;
            reg_file[13049] <= 8'h7C;
            reg_file[13050] <= 8'h15;
            reg_file[13051] <= 8'hFF;
            reg_file[13052] <= 8'h83;
            reg_file[13053] <= 8'hC7;
            reg_file[13054] <= 8'h05;
            reg_file[13055] <= 8'h00;
            reg_file[13056] <= 8'h13;
            reg_file[13057] <= 8'h07;
            reg_file[13058] <= 8'h17;
            reg_file[13059] <= 8'h00;
            reg_file[13060] <= 8'h93;
            reg_file[13061] <= 8'h85;
            reg_file[13062] <= 8'h15;
            reg_file[13063] <= 8'h00;
            reg_file[13064] <= 8'hA3;
            reg_file[13065] <= 8'h0F;
            reg_file[13066] <= 8'hF7;
            reg_file[13067] <= 8'hFE;
            reg_file[13068] <= 8'hE3;
            reg_file[13069] <= 8'h68;
            reg_file[13070] <= 8'h17;
            reg_file[13071] <= 8'hFF;
            reg_file[13072] <= 8'h67;
            reg_file[13073] <= 8'h80;
            reg_file[13074] <= 8'h00;
            reg_file[13075] <= 8'h00;
            reg_file[13076] <= 8'h83;
            reg_file[13077] <= 8'hC6;
            reg_file[13078] <= 8'h05;
            reg_file[13079] <= 8'h00;
            reg_file[13080] <= 8'h13;
            reg_file[13081] <= 8'h07;
            reg_file[13082] <= 8'h17;
            reg_file[13083] <= 8'h00;
            reg_file[13084] <= 8'h93;
            reg_file[13085] <= 8'h77;
            reg_file[13086] <= 8'h37;
            reg_file[13087] <= 8'h00;
            reg_file[13088] <= 8'hA3;
            reg_file[13089] <= 8'h0F;
            reg_file[13090] <= 8'hD7;
            reg_file[13091] <= 8'hFE;
            reg_file[13092] <= 8'h93;
            reg_file[13093] <= 8'h85;
            reg_file[13094] <= 8'h15;
            reg_file[13095] <= 8'h00;
            reg_file[13096] <= 8'hE3;
            reg_file[13097] <= 8'h80;
            reg_file[13098] <= 8'h07;
            reg_file[13099] <= 8'hF8;
            reg_file[13100] <= 8'h83;
            reg_file[13101] <= 8'hC6;
            reg_file[13102] <= 8'h05;
            reg_file[13103] <= 8'h00;
            reg_file[13104] <= 8'h13;
            reg_file[13105] <= 8'h07;
            reg_file[13106] <= 8'h17;
            reg_file[13107] <= 8'h00;
            reg_file[13108] <= 8'h93;
            reg_file[13109] <= 8'h77;
            reg_file[13110] <= 8'h37;
            reg_file[13111] <= 8'h00;
            reg_file[13112] <= 8'hA3;
            reg_file[13113] <= 8'h0F;
            reg_file[13114] <= 8'hD7;
            reg_file[13115] <= 8'hFE;
            reg_file[13116] <= 8'h93;
            reg_file[13117] <= 8'h85;
            reg_file[13118] <= 8'h15;
            reg_file[13119] <= 8'h00;
            reg_file[13120] <= 8'hE3;
            reg_file[13121] <= 8'h9A;
            reg_file[13122] <= 8'h07;
            reg_file[13123] <= 8'hFC;
            reg_file[13124] <= 8'h6F;
            reg_file[13125] <= 8'hF0;
            reg_file[13126] <= 8'h5F;
            reg_file[13127] <= 8'hF6;
            reg_file[13128] <= 8'h83;
            reg_file[13129] <= 8'hA6;
            reg_file[13130] <= 8'h45;
            reg_file[13131] <= 8'h00;
            reg_file[13132] <= 8'h83;
            reg_file[13133] <= 8'hA2;
            reg_file[13134] <= 8'h05;
            reg_file[13135] <= 8'h00;
            reg_file[13136] <= 8'h83;
            reg_file[13137] <= 8'hAF;
            reg_file[13138] <= 8'h85;
            reg_file[13139] <= 8'h00;
            reg_file[13140] <= 8'h03;
            reg_file[13141] <= 8'hAF;
            reg_file[13142] <= 8'hC5;
            reg_file[13143] <= 8'h00;
            reg_file[13144] <= 8'h83;
            reg_file[13145] <= 8'hAE;
            reg_file[13146] <= 8'h05;
            reg_file[13147] <= 8'h01;
            reg_file[13148] <= 8'h03;
            reg_file[13149] <= 8'hAE;
            reg_file[13150] <= 8'h45;
            reg_file[13151] <= 8'h01;
            reg_file[13152] <= 8'h03;
            reg_file[13153] <= 8'hA3;
            reg_file[13154] <= 8'h85;
            reg_file[13155] <= 8'h01;
            reg_file[13156] <= 8'h03;
            reg_file[13157] <= 8'hA8;
            reg_file[13158] <= 8'hC5;
            reg_file[13159] <= 8'h01;
            reg_file[13160] <= 8'h23;
            reg_file[13161] <= 8'h22;
            reg_file[13162] <= 8'hD7;
            reg_file[13163] <= 8'h00;
            reg_file[13164] <= 8'h83;
            reg_file[13165] <= 8'hA6;
            reg_file[13166] <= 8'h05;
            reg_file[13167] <= 8'h02;
            reg_file[13168] <= 8'h23;
            reg_file[13169] <= 8'h20;
            reg_file[13170] <= 8'h57;
            reg_file[13171] <= 8'h00;
            reg_file[13172] <= 8'h23;
            reg_file[13173] <= 8'h24;
            reg_file[13174] <= 8'hF7;
            reg_file[13175] <= 8'h01;
            reg_file[13176] <= 8'h23;
            reg_file[13177] <= 8'h26;
            reg_file[13178] <= 8'hE7;
            reg_file[13179] <= 8'h01;
            reg_file[13180] <= 8'h23;
            reg_file[13181] <= 8'h28;
            reg_file[13182] <= 8'hD7;
            reg_file[13183] <= 8'h01;
            reg_file[13184] <= 8'h23;
            reg_file[13185] <= 8'h2A;
            reg_file[13186] <= 8'hC7;
            reg_file[13187] <= 8'h01;
            reg_file[13188] <= 8'h23;
            reg_file[13189] <= 8'h2C;
            reg_file[13190] <= 8'h67;
            reg_file[13191] <= 8'h00;
            reg_file[13192] <= 8'h23;
            reg_file[13193] <= 8'h2E;
            reg_file[13194] <= 8'h07;
            reg_file[13195] <= 8'h01;
            reg_file[13196] <= 8'h23;
            reg_file[13197] <= 8'h20;
            reg_file[13198] <= 8'hD7;
            reg_file[13199] <= 8'h02;
            reg_file[13200] <= 8'h13;
            reg_file[13201] <= 8'h07;
            reg_file[13202] <= 8'h47;
            reg_file[13203] <= 8'h02;
            reg_file[13204] <= 8'h93;
            reg_file[13205] <= 8'h85;
            reg_file[13206] <= 8'h45;
            reg_file[13207] <= 8'h02;
            reg_file[13208] <= 8'hE3;
            reg_file[13209] <= 8'h68;
            reg_file[13210] <= 8'hF7;
            reg_file[13211] <= 8'hFA;
            reg_file[13212] <= 8'h6F;
            reg_file[13213] <= 8'hF0;
            reg_file[13214] <= 8'h9F;
            reg_file[13215] <= 8'hF1;
            reg_file[13216] <= 8'h13;
            reg_file[13217] <= 8'h03;
            reg_file[13218] <= 8'hF0;
            reg_file[13219] <= 8'h00;
            reg_file[13220] <= 8'h13;
            reg_file[13221] <= 8'h07;
            reg_file[13222] <= 8'h05;
            reg_file[13223] <= 8'h00;
            reg_file[13224] <= 8'h63;
            reg_file[13225] <= 8'h7E;
            reg_file[13226] <= 8'hC3;
            reg_file[13227] <= 8'h02;
            reg_file[13228] <= 8'h93;
            reg_file[13229] <= 8'h77;
            reg_file[13230] <= 8'hF7;
            reg_file[13231] <= 8'h00;
            reg_file[13232] <= 8'h63;
            reg_file[13233] <= 8'h90;
            reg_file[13234] <= 8'h07;
            reg_file[13235] <= 8'h0A;
            reg_file[13236] <= 8'h63;
            reg_file[13237] <= 8'h92;
            reg_file[13238] <= 8'h05;
            reg_file[13239] <= 8'h08;
            reg_file[13240] <= 8'h93;
            reg_file[13241] <= 8'h76;
            reg_file[13242] <= 8'h06;
            reg_file[13243] <= 8'hFF;
            reg_file[13244] <= 8'h13;
            reg_file[13245] <= 8'h76;
            reg_file[13246] <= 8'hF6;
            reg_file[13247] <= 8'h00;
            reg_file[13248] <= 8'hB3;
            reg_file[13249] <= 8'h86;
            reg_file[13250] <= 8'hE6;
            reg_file[13251] <= 8'h00;
            reg_file[13252] <= 8'h23;
            reg_file[13253] <= 8'h20;
            reg_file[13254] <= 8'hB7;
            reg_file[13255] <= 8'h00;
            reg_file[13256] <= 8'h23;
            reg_file[13257] <= 8'h22;
            reg_file[13258] <= 8'hB7;
            reg_file[13259] <= 8'h00;
            reg_file[13260] <= 8'h23;
            reg_file[13261] <= 8'h24;
            reg_file[13262] <= 8'hB7;
            reg_file[13263] <= 8'h00;
            reg_file[13264] <= 8'h23;
            reg_file[13265] <= 8'h26;
            reg_file[13266] <= 8'hB7;
            reg_file[13267] <= 8'h00;
            reg_file[13268] <= 8'h13;
            reg_file[13269] <= 8'h07;
            reg_file[13270] <= 8'h07;
            reg_file[13271] <= 8'h01;
            reg_file[13272] <= 8'hE3;
            reg_file[13273] <= 8'h66;
            reg_file[13274] <= 8'hD7;
            reg_file[13275] <= 8'hFE;
            reg_file[13276] <= 8'h63;
            reg_file[13277] <= 8'h14;
            reg_file[13278] <= 8'h06;
            reg_file[13279] <= 8'h00;
            reg_file[13280] <= 8'h67;
            reg_file[13281] <= 8'h80;
            reg_file[13282] <= 8'h00;
            reg_file[13283] <= 8'h00;
            reg_file[13284] <= 8'hB3;
            reg_file[13285] <= 8'h06;
            reg_file[13286] <= 8'hC3;
            reg_file[13287] <= 8'h40;
            reg_file[13288] <= 8'h93;
            reg_file[13289] <= 8'h96;
            reg_file[13290] <= 8'h26;
            reg_file[13291] <= 8'h00;
            reg_file[13292] <= 8'h97;
            reg_file[13293] <= 8'h02;
            reg_file[13294] <= 8'h00;
            reg_file[13295] <= 8'h00;
            reg_file[13296] <= 8'hB3;
            reg_file[13297] <= 8'h86;
            reg_file[13298] <= 8'h56;
            reg_file[13299] <= 8'h00;
            reg_file[13300] <= 8'h67;
            reg_file[13301] <= 8'h80;
            reg_file[13302] <= 8'hC6;
            reg_file[13303] <= 8'h00;
            reg_file[13304] <= 8'h23;
            reg_file[13305] <= 8'h07;
            reg_file[13306] <= 8'hB7;
            reg_file[13307] <= 8'h00;
            reg_file[13308] <= 8'hA3;
            reg_file[13309] <= 8'h06;
            reg_file[13310] <= 8'hB7;
            reg_file[13311] <= 8'h00;
            reg_file[13312] <= 8'h23;
            reg_file[13313] <= 8'h06;
            reg_file[13314] <= 8'hB7;
            reg_file[13315] <= 8'h00;
            reg_file[13316] <= 8'hA3;
            reg_file[13317] <= 8'h05;
            reg_file[13318] <= 8'hB7;
            reg_file[13319] <= 8'h00;
            reg_file[13320] <= 8'h23;
            reg_file[13321] <= 8'h05;
            reg_file[13322] <= 8'hB7;
            reg_file[13323] <= 8'h00;
            reg_file[13324] <= 8'hA3;
            reg_file[13325] <= 8'h04;
            reg_file[13326] <= 8'hB7;
            reg_file[13327] <= 8'h00;
            reg_file[13328] <= 8'h23;
            reg_file[13329] <= 8'h04;
            reg_file[13330] <= 8'hB7;
            reg_file[13331] <= 8'h00;
            reg_file[13332] <= 8'hA3;
            reg_file[13333] <= 8'h03;
            reg_file[13334] <= 8'hB7;
            reg_file[13335] <= 8'h00;
            reg_file[13336] <= 8'h23;
            reg_file[13337] <= 8'h03;
            reg_file[13338] <= 8'hB7;
            reg_file[13339] <= 8'h00;
            reg_file[13340] <= 8'hA3;
            reg_file[13341] <= 8'h02;
            reg_file[13342] <= 8'hB7;
            reg_file[13343] <= 8'h00;
            reg_file[13344] <= 8'h23;
            reg_file[13345] <= 8'h02;
            reg_file[13346] <= 8'hB7;
            reg_file[13347] <= 8'h00;
            reg_file[13348] <= 8'hA3;
            reg_file[13349] <= 8'h01;
            reg_file[13350] <= 8'hB7;
            reg_file[13351] <= 8'h00;
            reg_file[13352] <= 8'h23;
            reg_file[13353] <= 8'h01;
            reg_file[13354] <= 8'hB7;
            reg_file[13355] <= 8'h00;
            reg_file[13356] <= 8'hA3;
            reg_file[13357] <= 8'h00;
            reg_file[13358] <= 8'hB7;
            reg_file[13359] <= 8'h00;
            reg_file[13360] <= 8'h23;
            reg_file[13361] <= 8'h00;
            reg_file[13362] <= 8'hB7;
            reg_file[13363] <= 8'h00;
            reg_file[13364] <= 8'h67;
            reg_file[13365] <= 8'h80;
            reg_file[13366] <= 8'h00;
            reg_file[13367] <= 8'h00;
            reg_file[13368] <= 8'h93;
            reg_file[13369] <= 8'hF5;
            reg_file[13370] <= 8'hF5;
            reg_file[13371] <= 8'h0F;
            reg_file[13372] <= 8'h93;
            reg_file[13373] <= 8'h96;
            reg_file[13374] <= 8'h85;
            reg_file[13375] <= 8'h00;
            reg_file[13376] <= 8'hB3;
            reg_file[13377] <= 8'hE5;
            reg_file[13378] <= 8'hD5;
            reg_file[13379] <= 8'h00;
            reg_file[13380] <= 8'h93;
            reg_file[13381] <= 8'h96;
            reg_file[13382] <= 8'h05;
            reg_file[13383] <= 8'h01;
            reg_file[13384] <= 8'hB3;
            reg_file[13385] <= 8'hE5;
            reg_file[13386] <= 8'hD5;
            reg_file[13387] <= 8'h00;
            reg_file[13388] <= 8'h6F;
            reg_file[13389] <= 8'hF0;
            reg_file[13390] <= 8'hDF;
            reg_file[13391] <= 8'hF6;
            reg_file[13392] <= 8'h93;
            reg_file[13393] <= 8'h96;
            reg_file[13394] <= 8'h27;
            reg_file[13395] <= 8'h00;
            reg_file[13396] <= 8'h97;
            reg_file[13397] <= 8'h02;
            reg_file[13398] <= 8'h00;
            reg_file[13399] <= 8'h00;
            reg_file[13400] <= 8'hB3;
            reg_file[13401] <= 8'h86;
            reg_file[13402] <= 8'h56;
            reg_file[13403] <= 8'h00;
            reg_file[13404] <= 8'h93;
            reg_file[13405] <= 8'h82;
            reg_file[13406] <= 8'h00;
            reg_file[13407] <= 8'h00;
            reg_file[13408] <= 8'hE7;
            reg_file[13409] <= 8'h80;
            reg_file[13410] <= 8'h06;
            reg_file[13411] <= 8'hFA;
            reg_file[13412] <= 8'h93;
            reg_file[13413] <= 8'h80;
            reg_file[13414] <= 8'h02;
            reg_file[13415] <= 8'h00;
            reg_file[13416] <= 8'h93;
            reg_file[13417] <= 8'h87;
            reg_file[13418] <= 8'h07;
            reg_file[13419] <= 8'hFF;
            reg_file[13420] <= 8'h33;
            reg_file[13421] <= 8'h07;
            reg_file[13422] <= 8'hF7;
            reg_file[13423] <= 8'h40;
            reg_file[13424] <= 8'h33;
            reg_file[13425] <= 8'h06;
            reg_file[13426] <= 8'hF6;
            reg_file[13427] <= 8'h00;
            reg_file[13428] <= 8'hE3;
            reg_file[13429] <= 8'h78;
            reg_file[13430] <= 8'hC3;
            reg_file[13431] <= 8'hF6;
            reg_file[13432] <= 8'h6F;
            reg_file[13433] <= 8'hF0;
            reg_file[13434] <= 8'hDF;
            reg_file[13435] <= 8'hF3;
            reg_file[13436] <= 8'hB7;
            reg_file[13437] <= 8'h57;
            reg_file[13438] <= 8'h00;
            reg_file[13439] <= 8'h80;
            reg_file[13440] <= 8'h03;
            reg_file[13441] <= 8'hA7;
            reg_file[13442] <= 8'h07;
            reg_file[13443] <= 8'hCF;
            reg_file[13444] <= 8'h83;
            reg_file[13445] <= 8'h27;
            reg_file[13446] <= 8'h87;
            reg_file[13447] <= 8'h14;
            reg_file[13448] <= 8'h63;
            reg_file[13449] <= 8'h8C;
            reg_file[13450] <= 8'h07;
            reg_file[13451] <= 8'h04;
            reg_file[13452] <= 8'h03;
            reg_file[13453] <= 8'hA7;
            reg_file[13454] <= 8'h47;
            reg_file[13455] <= 8'h00;
            reg_file[13456] <= 8'h13;
            reg_file[13457] <= 8'h08;
            reg_file[13458] <= 8'hF0;
            reg_file[13459] <= 8'h01;
            reg_file[13460] <= 8'h63;
            reg_file[13461] <= 8'h4E;
            reg_file[13462] <= 8'hE8;
            reg_file[13463] <= 8'h06;
            reg_file[13464] <= 8'h13;
            reg_file[13465] <= 8'h18;
            reg_file[13466] <= 8'h27;
            reg_file[13467] <= 8'h00;
            reg_file[13468] <= 8'h63;
            reg_file[13469] <= 8'h06;
            reg_file[13470] <= 8'h05;
            reg_file[13471] <= 8'h02;
            reg_file[13472] <= 8'h33;
            reg_file[13473] <= 8'h83;
            reg_file[13474] <= 8'h07;
            reg_file[13475] <= 8'h01;
            reg_file[13476] <= 8'h23;
            reg_file[13477] <= 8'h24;
            reg_file[13478] <= 8'hC3;
            reg_file[13479] <= 8'h08;
            reg_file[13480] <= 8'h83;
            reg_file[13481] <= 8'hA8;
            reg_file[13482] <= 8'h87;
            reg_file[13483] <= 8'h18;
            reg_file[13484] <= 8'h13;
            reg_file[13485] <= 8'h06;
            reg_file[13486] <= 8'h10;
            reg_file[13487] <= 8'h00;
            reg_file[13488] <= 8'h33;
            reg_file[13489] <= 8'h16;
            reg_file[13490] <= 8'hE6;
            reg_file[13491] <= 8'h00;
            reg_file[13492] <= 8'hB3;
            reg_file[13493] <= 8'hE8;
            reg_file[13494] <= 8'hC8;
            reg_file[13495] <= 8'h00;
            reg_file[13496] <= 8'h23;
            reg_file[13497] <= 8'hA4;
            reg_file[13498] <= 8'h17;
            reg_file[13499] <= 8'h19;
            reg_file[13500] <= 8'h23;
            reg_file[13501] <= 8'h24;
            reg_file[13502] <= 8'hD3;
            reg_file[13503] <= 8'h10;
            reg_file[13504] <= 8'h93;
            reg_file[13505] <= 8'h06;
            reg_file[13506] <= 8'h20;
            reg_file[13507] <= 8'h00;
            reg_file[13508] <= 8'h63;
            reg_file[13509] <= 8'h04;
            reg_file[13510] <= 8'hD5;
            reg_file[13511] <= 8'h02;
            reg_file[13512] <= 8'h13;
            reg_file[13513] <= 8'h07;
            reg_file[13514] <= 8'h17;
            reg_file[13515] <= 8'h00;
            reg_file[13516] <= 8'h23;
            reg_file[13517] <= 8'hA2;
            reg_file[13518] <= 8'hE7;
            reg_file[13519] <= 8'h00;
            reg_file[13520] <= 8'hB3;
            reg_file[13521] <= 8'h87;
            reg_file[13522] <= 8'h07;
            reg_file[13523] <= 8'h01;
            reg_file[13524] <= 8'h23;
            reg_file[13525] <= 8'hA4;
            reg_file[13526] <= 8'hB7;
            reg_file[13527] <= 8'h00;
            reg_file[13528] <= 8'h13;
            reg_file[13529] <= 8'h05;
            reg_file[13530] <= 8'h00;
            reg_file[13531] <= 8'h00;
            reg_file[13532] <= 8'h67;
            reg_file[13533] <= 8'h80;
            reg_file[13534] <= 8'h00;
            reg_file[13535] <= 8'h00;
            reg_file[13536] <= 8'h93;
            reg_file[13537] <= 8'h07;
            reg_file[13538] <= 8'hC7;
            reg_file[13539] <= 8'h14;
            reg_file[13540] <= 8'h23;
            reg_file[13541] <= 8'h24;
            reg_file[13542] <= 8'hF7;
            reg_file[13543] <= 8'h14;
            reg_file[13544] <= 8'h6F;
            reg_file[13545] <= 8'hF0;
            reg_file[13546] <= 8'h5F;
            reg_file[13547] <= 8'hFA;
            reg_file[13548] <= 8'h83;
            reg_file[13549] <= 8'hA6;
            reg_file[13550] <= 8'hC7;
            reg_file[13551] <= 8'h18;
            reg_file[13552] <= 8'h13;
            reg_file[13553] <= 8'h07;
            reg_file[13554] <= 8'h17;
            reg_file[13555] <= 8'h00;
            reg_file[13556] <= 8'h23;
            reg_file[13557] <= 8'hA2;
            reg_file[13558] <= 8'hE7;
            reg_file[13559] <= 8'h00;
            reg_file[13560] <= 8'h33;
            reg_file[13561] <= 8'hE6;
            reg_file[13562] <= 8'hC6;
            reg_file[13563] <= 8'h00;
            reg_file[13564] <= 8'h23;
            reg_file[13565] <= 8'hA6;
            reg_file[13566] <= 8'hC7;
            reg_file[13567] <= 8'h18;
            reg_file[13568] <= 8'hB3;
            reg_file[13569] <= 8'h87;
            reg_file[13570] <= 8'h07;
            reg_file[13571] <= 8'h01;
            reg_file[13572] <= 8'h23;
            reg_file[13573] <= 8'hA4;
            reg_file[13574] <= 8'hB7;
            reg_file[13575] <= 8'h00;
            reg_file[13576] <= 8'h13;
            reg_file[13577] <= 8'h05;
            reg_file[13578] <= 8'h00;
            reg_file[13579] <= 8'h00;
            reg_file[13580] <= 8'h67;
            reg_file[13581] <= 8'h80;
            reg_file[13582] <= 8'h00;
            reg_file[13583] <= 8'h00;
            reg_file[13584] <= 8'h13;
            reg_file[13585] <= 8'h05;
            reg_file[13586] <= 8'hF0;
            reg_file[13587] <= 8'hFF;
            reg_file[13588] <= 8'h67;
            reg_file[13589] <= 8'h80;
            reg_file[13590] <= 8'h00;
            reg_file[13591] <= 8'h00;
            reg_file[13592] <= 8'h13;
            reg_file[13593] <= 8'h01;
            reg_file[13594] <= 8'h01;
            reg_file[13595] <= 8'hFD;
            reg_file[13596] <= 8'hB7;
            reg_file[13597] <= 8'h57;
            reg_file[13598] <= 8'h00;
            reg_file[13599] <= 8'h80;
            reg_file[13600] <= 8'h23;
            reg_file[13601] <= 8'h2C;
            reg_file[13602] <= 8'h41;
            reg_file[13603] <= 8'h01;
            reg_file[13604] <= 8'h03;
            reg_file[13605] <= 8'hAA;
            reg_file[13606] <= 8'h07;
            reg_file[13607] <= 8'hCF;
            reg_file[13608] <= 8'h23;
            reg_file[13609] <= 8'h20;
            reg_file[13610] <= 8'h21;
            reg_file[13611] <= 8'h03;
            reg_file[13612] <= 8'h23;
            reg_file[13613] <= 8'h26;
            reg_file[13614] <= 8'h11;
            reg_file[13615] <= 8'h02;
            reg_file[13616] <= 8'h03;
            reg_file[13617] <= 8'h29;
            reg_file[13618] <= 8'h8A;
            reg_file[13619] <= 8'h14;
            reg_file[13620] <= 8'h23;
            reg_file[13621] <= 8'h24;
            reg_file[13622] <= 8'h81;
            reg_file[13623] <= 8'h02;
            reg_file[13624] <= 8'h23;
            reg_file[13625] <= 8'h22;
            reg_file[13626] <= 8'h91;
            reg_file[13627] <= 8'h02;
            reg_file[13628] <= 8'h23;
            reg_file[13629] <= 8'h2E;
            reg_file[13630] <= 8'h31;
            reg_file[13631] <= 8'h01;
            reg_file[13632] <= 8'h23;
            reg_file[13633] <= 8'h2A;
            reg_file[13634] <= 8'h51;
            reg_file[13635] <= 8'h01;
            reg_file[13636] <= 8'h23;
            reg_file[13637] <= 8'h28;
            reg_file[13638] <= 8'h61;
            reg_file[13639] <= 8'h01;
            reg_file[13640] <= 8'h23;
            reg_file[13641] <= 8'h26;
            reg_file[13642] <= 8'h71;
            reg_file[13643] <= 8'h01;
            reg_file[13644] <= 8'h23;
            reg_file[13645] <= 8'h24;
            reg_file[13646] <= 8'h81;
            reg_file[13647] <= 8'h01;
            reg_file[13648] <= 8'h63;
            reg_file[13649] <= 8'h00;
            reg_file[13650] <= 8'h09;
            reg_file[13651] <= 8'h04;
            reg_file[13652] <= 8'h13;
            reg_file[13653] <= 8'h0B;
            reg_file[13654] <= 8'h05;
            reg_file[13655] <= 8'h00;
            reg_file[13656] <= 8'h93;
            reg_file[13657] <= 8'h8B;
            reg_file[13658] <= 8'h05;
            reg_file[13659] <= 8'h00;
            reg_file[13660] <= 8'h93;
            reg_file[13661] <= 8'h0A;
            reg_file[13662] <= 8'h10;
            reg_file[13663] <= 8'h00;
            reg_file[13664] <= 8'h93;
            reg_file[13665] <= 8'h09;
            reg_file[13666] <= 8'hF0;
            reg_file[13667] <= 8'hFF;
            reg_file[13668] <= 8'h83;
            reg_file[13669] <= 8'h24;
            reg_file[13670] <= 8'h49;
            reg_file[13671] <= 8'h00;
            reg_file[13672] <= 8'h13;
            reg_file[13673] <= 8'h84;
            reg_file[13674] <= 8'hF4;
            reg_file[13675] <= 8'hFF;
            reg_file[13676] <= 8'h63;
            reg_file[13677] <= 8'h42;
            reg_file[13678] <= 8'h04;
            reg_file[13679] <= 8'h02;
            reg_file[13680] <= 8'h93;
            reg_file[13681] <= 8'h94;
            reg_file[13682] <= 8'h24;
            reg_file[13683] <= 8'h00;
            reg_file[13684] <= 8'hB3;
            reg_file[13685] <= 8'h04;
            reg_file[13686] <= 8'h99;
            reg_file[13687] <= 8'h00;
            reg_file[13688] <= 8'h63;
            reg_file[13689] <= 8'h84;
            reg_file[13690] <= 8'h0B;
            reg_file[13691] <= 8'h04;
            reg_file[13692] <= 8'h83;
            reg_file[13693] <= 8'hA7;
            reg_file[13694] <= 8'h44;
            reg_file[13695] <= 8'h10;
            reg_file[13696] <= 8'h63;
            reg_file[13697] <= 8'h80;
            reg_file[13698] <= 8'h77;
            reg_file[13699] <= 8'h05;
            reg_file[13700] <= 8'h13;
            reg_file[13701] <= 8'h04;
            reg_file[13702] <= 8'hF4;
            reg_file[13703] <= 8'hFF;
            reg_file[13704] <= 8'h93;
            reg_file[13705] <= 8'h84;
            reg_file[13706] <= 8'hC4;
            reg_file[13707] <= 8'hFF;
            reg_file[13708] <= 8'hE3;
            reg_file[13709] <= 8'h16;
            reg_file[13710] <= 8'h34;
            reg_file[13711] <= 8'hFF;
            reg_file[13712] <= 8'h83;
            reg_file[13713] <= 8'h20;
            reg_file[13714] <= 8'hC1;
            reg_file[13715] <= 8'h02;
            reg_file[13716] <= 8'h03;
            reg_file[13717] <= 8'h24;
            reg_file[13718] <= 8'h81;
            reg_file[13719] <= 8'h02;
            reg_file[13720] <= 8'h83;
            reg_file[13721] <= 8'h24;
            reg_file[13722] <= 8'h41;
            reg_file[13723] <= 8'h02;
            reg_file[13724] <= 8'h03;
            reg_file[13725] <= 8'h29;
            reg_file[13726] <= 8'h01;
            reg_file[13727] <= 8'h02;
            reg_file[13728] <= 8'h83;
            reg_file[13729] <= 8'h29;
            reg_file[13730] <= 8'hC1;
            reg_file[13731] <= 8'h01;
            reg_file[13732] <= 8'h03;
            reg_file[13733] <= 8'h2A;
            reg_file[13734] <= 8'h81;
            reg_file[13735] <= 8'h01;
            reg_file[13736] <= 8'h83;
            reg_file[13737] <= 8'h2A;
            reg_file[13738] <= 8'h41;
            reg_file[13739] <= 8'h01;
            reg_file[13740] <= 8'h03;
            reg_file[13741] <= 8'h2B;
            reg_file[13742] <= 8'h01;
            reg_file[13743] <= 8'h01;
            reg_file[13744] <= 8'h83;
            reg_file[13745] <= 8'h2B;
            reg_file[13746] <= 8'hC1;
            reg_file[13747] <= 8'h00;
            reg_file[13748] <= 8'h03;
            reg_file[13749] <= 8'h2C;
            reg_file[13750] <= 8'h81;
            reg_file[13751] <= 8'h00;
            reg_file[13752] <= 8'h13;
            reg_file[13753] <= 8'h01;
            reg_file[13754] <= 8'h01;
            reg_file[13755] <= 8'h03;
            reg_file[13756] <= 8'h67;
            reg_file[13757] <= 8'h80;
            reg_file[13758] <= 8'h00;
            reg_file[13759] <= 8'h00;
            reg_file[13760] <= 8'h83;
            reg_file[13761] <= 8'h27;
            reg_file[13762] <= 8'h49;
            reg_file[13763] <= 8'h00;
            reg_file[13764] <= 8'h83;
            reg_file[13765] <= 8'hA6;
            reg_file[13766] <= 8'h44;
            reg_file[13767] <= 8'h00;
            reg_file[13768] <= 8'h93;
            reg_file[13769] <= 8'h87;
            reg_file[13770] <= 8'hF7;
            reg_file[13771] <= 8'hFF;
            reg_file[13772] <= 8'h63;
            reg_file[13773] <= 8'h8E;
            reg_file[13774] <= 8'h87;
            reg_file[13775] <= 8'h04;
            reg_file[13776] <= 8'h23;
            reg_file[13777] <= 8'hA2;
            reg_file[13778] <= 8'h04;
            reg_file[13779] <= 8'h00;
            reg_file[13780] <= 8'hE3;
            reg_file[13781] <= 8'h88;
            reg_file[13782] <= 8'h06;
            reg_file[13783] <= 8'hFA;
            reg_file[13784] <= 8'h83;
            reg_file[13785] <= 8'h27;
            reg_file[13786] <= 8'h89;
            reg_file[13787] <= 8'h18;
            reg_file[13788] <= 8'h33;
            reg_file[13789] <= 8'h97;
            reg_file[13790] <= 8'h8A;
            reg_file[13791] <= 8'h00;
            reg_file[13792] <= 8'h03;
            reg_file[13793] <= 8'h2C;
            reg_file[13794] <= 8'h49;
            reg_file[13795] <= 8'h00;
            reg_file[13796] <= 8'hB3;
            reg_file[13797] <= 8'h77;
            reg_file[13798] <= 8'hF7;
            reg_file[13799] <= 8'h00;
            reg_file[13800] <= 8'h63;
            reg_file[13801] <= 8'h92;
            reg_file[13802] <= 8'h07;
            reg_file[13803] <= 8'h02;
            reg_file[13804] <= 8'hE7;
            reg_file[13805] <= 8'h80;
            reg_file[13806] <= 8'h06;
            reg_file[13807] <= 8'h00;
            reg_file[13808] <= 8'h03;
            reg_file[13809] <= 8'h27;
            reg_file[13810] <= 8'h49;
            reg_file[13811] <= 8'h00;
            reg_file[13812] <= 8'h83;
            reg_file[13813] <= 8'h27;
            reg_file[13814] <= 8'h8A;
            reg_file[13815] <= 8'h14;
            reg_file[13816] <= 8'h63;
            reg_file[13817] <= 8'h14;
            reg_file[13818] <= 8'h87;
            reg_file[13819] <= 8'h01;
            reg_file[13820] <= 8'hE3;
            reg_file[13821] <= 8'h04;
            reg_file[13822] <= 8'hF9;
            reg_file[13823] <= 8'hF8;
            reg_file[13824] <= 8'hE3;
            reg_file[13825] <= 8'h88;
            reg_file[13826] <= 8'h07;
            reg_file[13827] <= 8'hF8;
            reg_file[13828] <= 8'h13;
            reg_file[13829] <= 8'h89;
            reg_file[13830] <= 8'h07;
            reg_file[13831] <= 8'h00;
            reg_file[13832] <= 8'h6F;
            reg_file[13833] <= 8'hF0;
            reg_file[13834] <= 8'hDF;
            reg_file[13835] <= 8'hF5;
            reg_file[13836] <= 8'h83;
            reg_file[13837] <= 8'h27;
            reg_file[13838] <= 8'hC9;
            reg_file[13839] <= 8'h18;
            reg_file[13840] <= 8'h83;
            reg_file[13841] <= 8'hA5;
            reg_file[13842] <= 8'h44;
            reg_file[13843] <= 8'h08;
            reg_file[13844] <= 8'h33;
            reg_file[13845] <= 8'h77;
            reg_file[13846] <= 8'hF7;
            reg_file[13847] <= 8'h00;
            reg_file[13848] <= 8'h63;
            reg_file[13849] <= 8'h1C;
            reg_file[13850] <= 8'h07;
            reg_file[13851] <= 8'h00;
            reg_file[13852] <= 8'h13;
            reg_file[13853] <= 8'h05;
            reg_file[13854] <= 8'h0B;
            reg_file[13855] <= 8'h00;
            reg_file[13856] <= 8'hE7;
            reg_file[13857] <= 8'h80;
            reg_file[13858] <= 8'h06;
            reg_file[13859] <= 8'h00;
            reg_file[13860] <= 8'h6F;
            reg_file[13861] <= 8'hF0;
            reg_file[13862] <= 8'hDF;
            reg_file[13863] <= 8'hFC;
            reg_file[13864] <= 8'h23;
            reg_file[13865] <= 8'h22;
            reg_file[13866] <= 8'h89;
            reg_file[13867] <= 8'h00;
            reg_file[13868] <= 8'h6F;
            reg_file[13869] <= 8'hF0;
            reg_file[13870] <= 8'h9F;
            reg_file[13871] <= 8'hFA;
            reg_file[13872] <= 8'h13;
            reg_file[13873] <= 8'h85;
            reg_file[13874] <= 8'h05;
            reg_file[13875] <= 8'h00;
            reg_file[13876] <= 8'hE7;
            reg_file[13877] <= 8'h80;
            reg_file[13878] <= 8'h06;
            reg_file[13879] <= 8'h00;
            reg_file[13880] <= 8'h6F;
            reg_file[13881] <= 8'hF0;
            reg_file[13882] <= 8'h9F;
            reg_file[13883] <= 8'hFB;
            reg_file[13884] <= 8'hAC;
            reg_file[13885] <= 8'h1B;
            reg_file[13886] <= 8'h00;
            reg_file[13887] <= 8'h80;
            reg_file[13888] <= 8'hA0;
            reg_file[13889] <= 8'h1E;
            reg_file[13890] <= 8'h00;
            reg_file[13891] <= 8'h80;
            reg_file[13892] <= 8'hA4;
            reg_file[13893] <= 8'h1B;
            reg_file[13894] <= 8'h00;
            reg_file[13895] <= 8'h80;
            reg_file[13896] <= 8'hA0;
            reg_file[13897] <= 8'h1E;
            reg_file[13898] <= 8'h00;
            reg_file[13899] <= 8'h80;
            reg_file[13900] <= 8'h88;
            reg_file[13901] <= 8'h1E;
            reg_file[13902] <= 8'h00;
            reg_file[13903] <= 8'h80;
            reg_file[13904] <= 8'hA0;
            reg_file[13905] <= 8'h1E;
            reg_file[13906] <= 8'h00;
            reg_file[13907] <= 8'h80;
            reg_file[13908] <= 8'hA4;
            reg_file[13909] <= 8'h1B;
            reg_file[13910] <= 8'h00;
            reg_file[13911] <= 8'h80;
            reg_file[13912] <= 8'hB0;
            reg_file[13913] <= 8'h1B;
            reg_file[13914] <= 8'h00;
            reg_file[13915] <= 8'h80;
            reg_file[13916] <= 8'hB0;
            reg_file[13917] <= 8'h1B;
            reg_file[13918] <= 8'h00;
            reg_file[13919] <= 8'h80;
            reg_file[13920] <= 8'h88;
            reg_file[13921] <= 8'h1E;
            reg_file[13922] <= 8'h00;
            reg_file[13923] <= 8'h80;
            reg_file[13924] <= 8'hA4;
            reg_file[13925] <= 8'h1B;
            reg_file[13926] <= 8'h00;
            reg_file[13927] <= 8'h80;
            reg_file[13928] <= 8'h78;
            reg_file[13929] <= 8'h1B;
            reg_file[13930] <= 8'h00;
            reg_file[13931] <= 8'h80;
            reg_file[13932] <= 8'h78;
            reg_file[13933] <= 8'h1B;
            reg_file[13934] <= 8'h00;
            reg_file[13935] <= 8'h80;
            reg_file[13936] <= 8'h78;
            reg_file[13937] <= 8'h1B;
            reg_file[13938] <= 8'h00;
            reg_file[13939] <= 8'h80;
            reg_file[13940] <= 8'hC0;
            reg_file[13941] <= 8'h1B;
            reg_file[13942] <= 8'h00;
            reg_file[13943] <= 8'h80;
            reg_file[13944] <= 8'hC8;
            reg_file[13945] <= 8'h23;
            reg_file[13946] <= 8'h00;
            reg_file[13947] <= 8'h80;
            reg_file[13948] <= 8'hC8;
            reg_file[13949] <= 8'h23;
            reg_file[13950] <= 8'h00;
            reg_file[13951] <= 8'h80;
            reg_file[13952] <= 8'hEC;
            reg_file[13953] <= 8'h23;
            reg_file[13954] <= 8'h00;
            reg_file[13955] <= 8'h80;
            reg_file[13956] <= 8'hBC;
            reg_file[13957] <= 8'h23;
            reg_file[13958] <= 8'h00;
            reg_file[13959] <= 8'h80;
            reg_file[13960] <= 8'hBC;
            reg_file[13961] <= 8'h23;
            reg_file[13962] <= 8'h00;
            reg_file[13963] <= 8'h80;
            reg_file[13964] <= 8'h3C;
            reg_file[13965] <= 8'h21;
            reg_file[13966] <= 8'h00;
            reg_file[13967] <= 8'h80;
            reg_file[13968] <= 8'hEC;
            reg_file[13969] <= 8'h23;
            reg_file[13970] <= 8'h00;
            reg_file[13971] <= 8'h80;
            reg_file[13972] <= 8'hBC;
            reg_file[13973] <= 8'h23;
            reg_file[13974] <= 8'h00;
            reg_file[13975] <= 8'h80;
            reg_file[13976] <= 8'h3C;
            reg_file[13977] <= 8'h21;
            reg_file[13978] <= 8'h00;
            reg_file[13979] <= 8'h80;
            reg_file[13980] <= 8'hBC;
            reg_file[13981] <= 8'h23;
            reg_file[13982] <= 8'h00;
            reg_file[13983] <= 8'h80;
            reg_file[13984] <= 8'hEC;
            reg_file[13985] <= 8'h23;
            reg_file[13986] <= 8'h00;
            reg_file[13987] <= 8'h80;
            reg_file[13988] <= 8'hB8;
            reg_file[13989] <= 8'h23;
            reg_file[13990] <= 8'h00;
            reg_file[13991] <= 8'h80;
            reg_file[13992] <= 8'hB8;
            reg_file[13993] <= 8'h23;
            reg_file[13994] <= 8'h00;
            reg_file[13995] <= 8'h80;
            reg_file[13996] <= 8'hB8;
            reg_file[13997] <= 8'h23;
            reg_file[13998] <= 8'h00;
            reg_file[13999] <= 8'h80;
            reg_file[14000] <= 8'h60;
            reg_file[14001] <= 8'h26;
            reg_file[14002] <= 8'h00;
            reg_file[14003] <= 8'h80;
            reg_file[14004] <= 8'h00;
            reg_file[14005] <= 8'h01;
            reg_file[14006] <= 8'h02;
            reg_file[14007] <= 8'h02;
            reg_file[14008] <= 8'h03;
            reg_file[14009] <= 8'h03;
            reg_file[14010] <= 8'h03;
            reg_file[14011] <= 8'h03;
            reg_file[14012] <= 8'h04;
            reg_file[14013] <= 8'h04;
            reg_file[14014] <= 8'h04;
            reg_file[14015] <= 8'h04;
            reg_file[14016] <= 8'h04;
            reg_file[14017] <= 8'h04;
            reg_file[14018] <= 8'h04;
            reg_file[14019] <= 8'h04;
            reg_file[14020] <= 8'h05;
            reg_file[14021] <= 8'h05;
            reg_file[14022] <= 8'h05;
            reg_file[14023] <= 8'h05;
            reg_file[14024] <= 8'h05;
            reg_file[14025] <= 8'h05;
            reg_file[14026] <= 8'h05;
            reg_file[14027] <= 8'h05;
            reg_file[14028] <= 8'h05;
            reg_file[14029] <= 8'h05;
            reg_file[14030] <= 8'h05;
            reg_file[14031] <= 8'h05;
            reg_file[14032] <= 8'h05;
            reg_file[14033] <= 8'h05;
            reg_file[14034] <= 8'h05;
            reg_file[14035] <= 8'h05;
            reg_file[14036] <= 8'h06;
            reg_file[14037] <= 8'h06;
            reg_file[14038] <= 8'h06;
            reg_file[14039] <= 8'h06;
            reg_file[14040] <= 8'h06;
            reg_file[14041] <= 8'h06;
            reg_file[14042] <= 8'h06;
            reg_file[14043] <= 8'h06;
            reg_file[14044] <= 8'h06;
            reg_file[14045] <= 8'h06;
            reg_file[14046] <= 8'h06;
            reg_file[14047] <= 8'h06;
            reg_file[14048] <= 8'h06;
            reg_file[14049] <= 8'h06;
            reg_file[14050] <= 8'h06;
            reg_file[14051] <= 8'h06;
            reg_file[14052] <= 8'h06;
            reg_file[14053] <= 8'h06;
            reg_file[14054] <= 8'h06;
            reg_file[14055] <= 8'h06;
            reg_file[14056] <= 8'h06;
            reg_file[14057] <= 8'h06;
            reg_file[14058] <= 8'h06;
            reg_file[14059] <= 8'h06;
            reg_file[14060] <= 8'h06;
            reg_file[14061] <= 8'h06;
            reg_file[14062] <= 8'h06;
            reg_file[14063] <= 8'h06;
            reg_file[14064] <= 8'h06;
            reg_file[14065] <= 8'h06;
            reg_file[14066] <= 8'h06;
            reg_file[14067] <= 8'h06;
            reg_file[14068] <= 8'h07;
            reg_file[14069] <= 8'h07;
            reg_file[14070] <= 8'h07;
            reg_file[14071] <= 8'h07;
            reg_file[14072] <= 8'h07;
            reg_file[14073] <= 8'h07;
            reg_file[14074] <= 8'h07;
            reg_file[14075] <= 8'h07;
            reg_file[14076] <= 8'h07;
            reg_file[14077] <= 8'h07;
            reg_file[14078] <= 8'h07;
            reg_file[14079] <= 8'h07;
            reg_file[14080] <= 8'h07;
            reg_file[14081] <= 8'h07;
            reg_file[14082] <= 8'h07;
            reg_file[14083] <= 8'h07;
            reg_file[14084] <= 8'h07;
            reg_file[14085] <= 8'h07;
            reg_file[14086] <= 8'h07;
            reg_file[14087] <= 8'h07;
            reg_file[14088] <= 8'h07;
            reg_file[14089] <= 8'h07;
            reg_file[14090] <= 8'h07;
            reg_file[14091] <= 8'h07;
            reg_file[14092] <= 8'h07;
            reg_file[14093] <= 8'h07;
            reg_file[14094] <= 8'h07;
            reg_file[14095] <= 8'h07;
            reg_file[14096] <= 8'h07;
            reg_file[14097] <= 8'h07;
            reg_file[14098] <= 8'h07;
            reg_file[14099] <= 8'h07;
            reg_file[14100] <= 8'h07;
            reg_file[14101] <= 8'h07;
            reg_file[14102] <= 8'h07;
            reg_file[14103] <= 8'h07;
            reg_file[14104] <= 8'h07;
            reg_file[14105] <= 8'h07;
            reg_file[14106] <= 8'h07;
            reg_file[14107] <= 8'h07;
            reg_file[14108] <= 8'h07;
            reg_file[14109] <= 8'h07;
            reg_file[14110] <= 8'h07;
            reg_file[14111] <= 8'h07;
            reg_file[14112] <= 8'h07;
            reg_file[14113] <= 8'h07;
            reg_file[14114] <= 8'h07;
            reg_file[14115] <= 8'h07;
            reg_file[14116] <= 8'h07;
            reg_file[14117] <= 8'h07;
            reg_file[14118] <= 8'h07;
            reg_file[14119] <= 8'h07;
            reg_file[14120] <= 8'h07;
            reg_file[14121] <= 8'h07;
            reg_file[14122] <= 8'h07;
            reg_file[14123] <= 8'h07;
            reg_file[14124] <= 8'h07;
            reg_file[14125] <= 8'h07;
            reg_file[14126] <= 8'h07;
            reg_file[14127] <= 8'h07;
            reg_file[14128] <= 8'h07;
            reg_file[14129] <= 8'h07;
            reg_file[14130] <= 8'h07;
            reg_file[14131] <= 8'h07;
            reg_file[14132] <= 8'h08;
            reg_file[14133] <= 8'h08;
            reg_file[14134] <= 8'h08;
            reg_file[14135] <= 8'h08;
            reg_file[14136] <= 8'h08;
            reg_file[14137] <= 8'h08;
            reg_file[14138] <= 8'h08;
            reg_file[14139] <= 8'h08;
            reg_file[14140] <= 8'h08;
            reg_file[14141] <= 8'h08;
            reg_file[14142] <= 8'h08;
            reg_file[14143] <= 8'h08;
            reg_file[14144] <= 8'h08;
            reg_file[14145] <= 8'h08;
            reg_file[14146] <= 8'h08;
            reg_file[14147] <= 8'h08;
            reg_file[14148] <= 8'h08;
            reg_file[14149] <= 8'h08;
            reg_file[14150] <= 8'h08;
            reg_file[14151] <= 8'h08;
            reg_file[14152] <= 8'h08;
            reg_file[14153] <= 8'h08;
            reg_file[14154] <= 8'h08;
            reg_file[14155] <= 8'h08;
            reg_file[14156] <= 8'h08;
            reg_file[14157] <= 8'h08;
            reg_file[14158] <= 8'h08;
            reg_file[14159] <= 8'h08;
            reg_file[14160] <= 8'h08;
            reg_file[14161] <= 8'h08;
            reg_file[14162] <= 8'h08;
            reg_file[14163] <= 8'h08;
            reg_file[14164] <= 8'h08;
            reg_file[14165] <= 8'h08;
            reg_file[14166] <= 8'h08;
            reg_file[14167] <= 8'h08;
            reg_file[14168] <= 8'h08;
            reg_file[14169] <= 8'h08;
            reg_file[14170] <= 8'h08;
            reg_file[14171] <= 8'h08;
            reg_file[14172] <= 8'h08;
            reg_file[14173] <= 8'h08;
            reg_file[14174] <= 8'h08;
            reg_file[14175] <= 8'h08;
            reg_file[14176] <= 8'h08;
            reg_file[14177] <= 8'h08;
            reg_file[14178] <= 8'h08;
            reg_file[14179] <= 8'h08;
            reg_file[14180] <= 8'h08;
            reg_file[14181] <= 8'h08;
            reg_file[14182] <= 8'h08;
            reg_file[14183] <= 8'h08;
            reg_file[14184] <= 8'h08;
            reg_file[14185] <= 8'h08;
            reg_file[14186] <= 8'h08;
            reg_file[14187] <= 8'h08;
            reg_file[14188] <= 8'h08;
            reg_file[14189] <= 8'h08;
            reg_file[14190] <= 8'h08;
            reg_file[14191] <= 8'h08;
            reg_file[14192] <= 8'h08;
            reg_file[14193] <= 8'h08;
            reg_file[14194] <= 8'h08;
            reg_file[14195] <= 8'h08;
            reg_file[14196] <= 8'h08;
            reg_file[14197] <= 8'h08;
            reg_file[14198] <= 8'h08;
            reg_file[14199] <= 8'h08;
            reg_file[14200] <= 8'h08;
            reg_file[14201] <= 8'h08;
            reg_file[14202] <= 8'h08;
            reg_file[14203] <= 8'h08;
            reg_file[14204] <= 8'h08;
            reg_file[14205] <= 8'h08;
            reg_file[14206] <= 8'h08;
            reg_file[14207] <= 8'h08;
            reg_file[14208] <= 8'h08;
            reg_file[14209] <= 8'h08;
            reg_file[14210] <= 8'h08;
            reg_file[14211] <= 8'h08;
            reg_file[14212] <= 8'h08;
            reg_file[14213] <= 8'h08;
            reg_file[14214] <= 8'h08;
            reg_file[14215] <= 8'h08;
            reg_file[14216] <= 8'h08;
            reg_file[14217] <= 8'h08;
            reg_file[14218] <= 8'h08;
            reg_file[14219] <= 8'h08;
            reg_file[14220] <= 8'h08;
            reg_file[14221] <= 8'h08;
            reg_file[14222] <= 8'h08;
            reg_file[14223] <= 8'h08;
            reg_file[14224] <= 8'h08;
            reg_file[14225] <= 8'h08;
            reg_file[14226] <= 8'h08;
            reg_file[14227] <= 8'h08;
            reg_file[14228] <= 8'h08;
            reg_file[14229] <= 8'h08;
            reg_file[14230] <= 8'h08;
            reg_file[14231] <= 8'h08;
            reg_file[14232] <= 8'h08;
            reg_file[14233] <= 8'h08;
            reg_file[14234] <= 8'h08;
            reg_file[14235] <= 8'h08;
            reg_file[14236] <= 8'h08;
            reg_file[14237] <= 8'h08;
            reg_file[14238] <= 8'h08;
            reg_file[14239] <= 8'h08;
            reg_file[14240] <= 8'h08;
            reg_file[14241] <= 8'h08;
            reg_file[14242] <= 8'h08;
            reg_file[14243] <= 8'h08;
            reg_file[14244] <= 8'h08;
            reg_file[14245] <= 8'h08;
            reg_file[14246] <= 8'h08;
            reg_file[14247] <= 8'h08;
            reg_file[14248] <= 8'h08;
            reg_file[14249] <= 8'h08;
            reg_file[14250] <= 8'h08;
            reg_file[14251] <= 8'h08;
            reg_file[14252] <= 8'h08;
            reg_file[14253] <= 8'h08;
            reg_file[14254] <= 8'h08;
            reg_file[14255] <= 8'h08;
            reg_file[14256] <= 8'h08;
            reg_file[14257] <= 8'h08;
            reg_file[14258] <= 8'h08;
            reg_file[14259] <= 8'h08;
            reg_file[14260] <= 8'h10;
            reg_file[14261] <= 8'h00;
            reg_file[14262] <= 8'h00;
            reg_file[14263] <= 8'h00;
            reg_file[14264] <= 8'h00;
            reg_file[14265] <= 8'h00;
            reg_file[14266] <= 8'h00;
            reg_file[14267] <= 8'h00;
            reg_file[14268] <= 8'h03;
            reg_file[14269] <= 8'h7A;
            reg_file[14270] <= 8'h52;
            reg_file[14271] <= 8'h00;
            reg_file[14272] <= 8'h01;
            reg_file[14273] <= 8'h7C;
            reg_file[14274] <= 8'h01;
            reg_file[14275] <= 8'h01;
            reg_file[14276] <= 8'h1B;
            reg_file[14277] <= 8'h0D;
            reg_file[14278] <= 8'h02;
            reg_file[14279] <= 8'h00;
            reg_file[14280] <= 8'h10;
            reg_file[14281] <= 8'h00;
            reg_file[14282] <= 8'h00;
            reg_file[14283] <= 8'h00;
            reg_file[14284] <= 8'h18;
            reg_file[14285] <= 8'h00;
            reg_file[14286] <= 8'h00;
            reg_file[14287] <= 8'h00;
            reg_file[14288] <= 8'h80;
            reg_file[14289] <= 8'hD2;
            reg_file[14290] <= 8'hFF;
            reg_file[14291] <= 8'hFF;
            reg_file[14292] <= 8'h08;
            reg_file[14293] <= 8'h00;
            reg_file[14294] <= 8'h00;
            reg_file[14295] <= 8'h00;
            reg_file[14296] <= 8'h00;
            reg_file[14297] <= 8'h00;
            reg_file[14298] <= 8'h00;
            reg_file[14299] <= 8'h00;
            reg_file[14300] <= 8'h10;
            reg_file[14301] <= 8'h00;
            reg_file[14302] <= 8'h00;
            reg_file[14303] <= 8'h00;
            reg_file[14304] <= 8'h2C;
            reg_file[14305] <= 8'h00;
            reg_file[14306] <= 8'h00;
            reg_file[14307] <= 8'h00;
            reg_file[14308] <= 8'h74;
            reg_file[14309] <= 8'hD2;
            reg_file[14310] <= 8'hFF;
            reg_file[14311] <= 8'hFF;
            reg_file[14312] <= 8'h08;
            reg_file[14313] <= 8'h00;
            reg_file[14314] <= 8'h00;
            reg_file[14315] <= 8'h00;
            reg_file[14316] <= 8'h00;
            reg_file[14317] <= 8'h00;
            reg_file[14318] <= 8'h00;
            reg_file[14319] <= 8'h00;
            reg_file[14320] <= 8'h10;
            reg_file[14321] <= 8'h00;
            reg_file[14322] <= 8'h00;
            reg_file[14323] <= 8'h00;
            reg_file[14324] <= 8'h40;
            reg_file[14325] <= 8'h00;
            reg_file[14326] <= 8'h00;
            reg_file[14327] <= 8'h00;
            reg_file[14328] <= 8'h68;
            reg_file[14329] <= 8'hD2;
            reg_file[14330] <= 8'hFF;
            reg_file[14331] <= 8'hFF;
            reg_file[14332] <= 8'h08;
            reg_file[14333] <= 8'h00;
            reg_file[14334] <= 8'h00;
            reg_file[14335] <= 8'h00;
            reg_file[14336] <= 8'h00;
            reg_file[14337] <= 8'h00;
            reg_file[14338] <= 8'h00;
            reg_file[14339] <= 8'h00;
            reg_file[14340] <= 8'h10;
            reg_file[14341] <= 8'h00;
            reg_file[14342] <= 8'h00;
            reg_file[14343] <= 8'h00;
            reg_file[14344] <= 8'h54;
            reg_file[14345] <= 8'h00;
            reg_file[14346] <= 8'h00;
            reg_file[14347] <= 8'h00;
            reg_file[14348] <= 8'h5C;
            reg_file[14349] <= 8'hD2;
            reg_file[14350] <= 8'hFF;
            reg_file[14351] <= 8'hFF;
            reg_file[14352] <= 8'h08;
            reg_file[14353] <= 8'h00;
            reg_file[14354] <= 8'h00;
            reg_file[14355] <= 8'h00;
            reg_file[14356] <= 8'h00;
            reg_file[14357] <= 8'h00;
            reg_file[14358] <= 8'h00;
            reg_file[14359] <= 8'h00;
            reg_file[14360] <= 8'h10;
            reg_file[14361] <= 8'h00;
            reg_file[14362] <= 8'h00;
            reg_file[14363] <= 8'h00;
            reg_file[14364] <= 8'h68;
            reg_file[14365] <= 8'h00;
            reg_file[14366] <= 8'h00;
            reg_file[14367] <= 8'h00;
            reg_file[14368] <= 8'h50;
            reg_file[14369] <= 8'hD2;
            reg_file[14370] <= 8'hFF;
            reg_file[14371] <= 8'hFF;
            reg_file[14372] <= 8'h08;
            reg_file[14373] <= 8'h00;
            reg_file[14374] <= 8'h00;
            reg_file[14375] <= 8'h00;
            reg_file[14376] <= 8'h00;
            reg_file[14377] <= 8'h00;
            reg_file[14378] <= 8'h00;
            reg_file[14379] <= 8'h00;
            reg_file[14380] <= 8'h10;
            reg_file[14381] <= 8'h00;
            reg_file[14382] <= 8'h00;
            reg_file[14383] <= 8'h00;
            reg_file[14384] <= 8'h7C;
            reg_file[14385] <= 8'h00;
            reg_file[14386] <= 8'h00;
            reg_file[14387] <= 8'h00;
            reg_file[14388] <= 8'h44;
            reg_file[14389] <= 8'hD2;
            reg_file[14390] <= 8'hFF;
            reg_file[14391] <= 8'hFF;
            reg_file[14392] <= 8'h08;
            reg_file[14393] <= 8'h00;
            reg_file[14394] <= 8'h00;
            reg_file[14395] <= 8'h00;
            reg_file[14396] <= 8'h00;
            reg_file[14397] <= 8'h00;
            reg_file[14398] <= 8'h00;
            reg_file[14399] <= 8'h00;
            reg_file[14400] <= 8'h10;
            reg_file[14401] <= 8'h00;
            reg_file[14402] <= 8'h00;
            reg_file[14403] <= 8'h00;
            reg_file[14404] <= 8'h90;
            reg_file[14405] <= 8'h00;
            reg_file[14406] <= 8'h00;
            reg_file[14407] <= 8'h00;
            reg_file[14408] <= 8'h38;
            reg_file[14409] <= 8'hD2;
            reg_file[14410] <= 8'hFF;
            reg_file[14411] <= 8'hFF;
            reg_file[14412] <= 8'h08;
            reg_file[14413] <= 8'h00;
            reg_file[14414] <= 8'h00;
            reg_file[14415] <= 8'h00;
            reg_file[14416] <= 8'h00;
            reg_file[14417] <= 8'h00;
            reg_file[14418] <= 8'h00;
            reg_file[14419] <= 8'h00;
            reg_file[14420] <= 8'h10;
            reg_file[14421] <= 8'h00;
            reg_file[14422] <= 8'h00;
            reg_file[14423] <= 8'h00;
            reg_file[14424] <= 8'hA4;
            reg_file[14425] <= 8'h00;
            reg_file[14426] <= 8'h00;
            reg_file[14427] <= 8'h00;
            reg_file[14428] <= 8'h2C;
            reg_file[14429] <= 8'hD2;
            reg_file[14430] <= 8'hFF;
            reg_file[14431] <= 8'hFF;
            reg_file[14432] <= 8'h08;
            reg_file[14433] <= 8'h00;
            reg_file[14434] <= 8'h00;
            reg_file[14435] <= 8'h00;
            reg_file[14436] <= 8'h00;
            reg_file[14437] <= 8'h00;
            reg_file[14438] <= 8'h00;
            reg_file[14439] <= 8'h00;
            reg_file[14440] <= 8'h10;
            reg_file[14441] <= 8'h00;
            reg_file[14442] <= 8'h00;
            reg_file[14443] <= 8'h00;
            reg_file[14444] <= 8'hB8;
            reg_file[14445] <= 8'h00;
            reg_file[14446] <= 8'h00;
            reg_file[14447] <= 8'h00;
            reg_file[14448] <= 8'h20;
            reg_file[14449] <= 8'hD2;
            reg_file[14450] <= 8'hFF;
            reg_file[14451] <= 8'hFF;
            reg_file[14452] <= 8'h08;
            reg_file[14453] <= 8'h00;
            reg_file[14454] <= 8'h00;
            reg_file[14455] <= 8'h00;
            reg_file[14456] <= 8'h00;
            reg_file[14457] <= 8'h00;
            reg_file[14458] <= 8'h00;
            reg_file[14459] <= 8'h00;
            reg_file[14460] <= 8'h10;
            reg_file[14461] <= 8'h00;
            reg_file[14462] <= 8'h00;
            reg_file[14463] <= 8'h00;
            reg_file[14464] <= 8'hCC;
            reg_file[14465] <= 8'h00;
            reg_file[14466] <= 8'h00;
            reg_file[14467] <= 8'h00;
            reg_file[14468] <= 8'h14;
            reg_file[14469] <= 8'hD2;
            reg_file[14470] <= 8'hFF;
            reg_file[14471] <= 8'hFF;
            reg_file[14472] <= 8'h08;
            reg_file[14473] <= 8'h00;
            reg_file[14474] <= 8'h00;
            reg_file[14475] <= 8'h00;
            reg_file[14476] <= 8'h00;
            reg_file[14477] <= 8'h00;
            reg_file[14478] <= 8'h00;
            reg_file[14479] <= 8'h00;
            reg_file[14480] <= 8'h10;
            reg_file[14481] <= 8'h00;
            reg_file[14482] <= 8'h00;
            reg_file[14483] <= 8'h00;
            reg_file[14484] <= 8'hE0;
            reg_file[14485] <= 8'h00;
            reg_file[14486] <= 8'h00;
            reg_file[14487] <= 8'h00;
            reg_file[14488] <= 8'h08;
            reg_file[14489] <= 8'hD2;
            reg_file[14490] <= 8'hFF;
            reg_file[14491] <= 8'hFF;
            reg_file[14492] <= 8'h08;
            reg_file[14493] <= 8'h00;
            reg_file[14494] <= 8'h00;
            reg_file[14495] <= 8'h00;
            reg_file[14496] <= 8'h00;
            reg_file[14497] <= 8'h00;
            reg_file[14498] <= 8'h00;
            reg_file[14499] <= 8'h00;
            reg_file[14500] <= 8'h10;
            reg_file[14501] <= 8'h00;
            reg_file[14502] <= 8'h00;
            reg_file[14503] <= 8'h00;
            reg_file[14504] <= 8'hF4;
            reg_file[14505] <= 8'h00;
            reg_file[14506] <= 8'h00;
            reg_file[14507] <= 8'h00;
            reg_file[14508] <= 8'hFC;
            reg_file[14509] <= 8'hD1;
            reg_file[14510] <= 8'hFF;
            reg_file[14511] <= 8'hFF;
            reg_file[14512] <= 8'h08;
            reg_file[14513] <= 8'h00;
            reg_file[14514] <= 8'h00;
            reg_file[14515] <= 8'h00;
            reg_file[14516] <= 8'h00;
            reg_file[14517] <= 8'h00;
            reg_file[14518] <= 8'h00;
            reg_file[14519] <= 8'h00;
            reg_file[14520] <= 8'h00;
            reg_file[14521] <= 8'h00;
            reg_file[14522] <= 8'h00;
            reg_file[14523] <= 8'h00;
            reg_file[14524] <= 8'h00;
            reg_file[14525] <= 8'h00;
            reg_file[14526] <= 8'h00;
            reg_file[14527] <= 8'h00;
            reg_file[14528] <= 8'h00;
            reg_file[14529] <= 8'h00;
            reg_file[14530] <= 8'h00;
            reg_file[14531] <= 8'h00;
            reg_file[14532] <= 8'h00;
            reg_file[14533] <= 8'h00;
            reg_file[14534] <= 8'h00;
            reg_file[14535] <= 8'h00;
            reg_file[14536] <= 8'h00;
            reg_file[14537] <= 8'h00;
            reg_file[14538] <= 8'h00;
            reg_file[14539] <= 8'h00;
            reg_file[14540] <= 8'h00;
            reg_file[14541] <= 8'h00;
            reg_file[14542] <= 8'h00;
            reg_file[14543] <= 8'h00;
            reg_file[14544] <= 8'h00;
            reg_file[14545] <= 8'h00;
            reg_file[14546] <= 8'h00;
            reg_file[14547] <= 8'h00;
            reg_file[14548] <= 8'h00;
            reg_file[14549] <= 8'h00;
            reg_file[14550] <= 8'h00;
            reg_file[14551] <= 8'h00;
            reg_file[14552] <= 8'h00;
            reg_file[14553] <= 8'h00;
            reg_file[14554] <= 8'h00;
            reg_file[14555] <= 8'h00;
            reg_file[14556] <= 8'h00;
            reg_file[14557] <= 8'h00;
            reg_file[14558] <= 8'h00;
            reg_file[14559] <= 8'h00;
            reg_file[14560] <= 8'h00;
            reg_file[14561] <= 8'h00;
            reg_file[14562] <= 8'h00;
            reg_file[14563] <= 8'h00;
            reg_file[14564] <= 8'h00;
            reg_file[14565] <= 8'h00;
            reg_file[14566] <= 8'h00;
            reg_file[14567] <= 8'h00;
            reg_file[14568] <= 8'h00;
            reg_file[14569] <= 8'h00;
            reg_file[14570] <= 8'h00;
            reg_file[14571] <= 8'h00;
            reg_file[14572] <= 8'h00;
            reg_file[14573] <= 8'h00;
            reg_file[14574] <= 8'h00;
            reg_file[14575] <= 8'h00;
            reg_file[14576] <= 8'h00;
            reg_file[14577] <= 8'h00;
            reg_file[14578] <= 8'h00;
            reg_file[14579] <= 8'h00;
            reg_file[14580] <= 8'h00;
            reg_file[14581] <= 8'h00;
            reg_file[14582] <= 8'h00;
            reg_file[14583] <= 8'h00;
            reg_file[14584] <= 8'h00;
            reg_file[14585] <= 8'h00;
            reg_file[14586] <= 8'h00;
            reg_file[14587] <= 8'h00;
            reg_file[14588] <= 8'h00;
            reg_file[14589] <= 8'h00;
            reg_file[14590] <= 8'h00;
            reg_file[14591] <= 8'h00;
            reg_file[14592] <= 8'h00;
            reg_file[14593] <= 8'h00;
            reg_file[14594] <= 8'h00;
            reg_file[14595] <= 8'h00;
            reg_file[14596] <= 8'h00;
            reg_file[14597] <= 8'h00;
            reg_file[14598] <= 8'h00;
            reg_file[14599] <= 8'h00;
            reg_file[14600] <= 8'h00;
            reg_file[14601] <= 8'h00;
            reg_file[14602] <= 8'h00;
            reg_file[14603] <= 8'h00;
            reg_file[14604] <= 8'h00;
            reg_file[14605] <= 8'h00;
            reg_file[14606] <= 8'h00;
            reg_file[14607] <= 8'h00;
            reg_file[14608] <= 8'h00;
            reg_file[14609] <= 8'h00;
            reg_file[14610] <= 8'h00;
            reg_file[14611] <= 8'h00;
            reg_file[14612] <= 8'h00;
            reg_file[14613] <= 8'h00;
            reg_file[14614] <= 8'h00;
            reg_file[14615] <= 8'h00;
            reg_file[14616] <= 8'h00;
            reg_file[14617] <= 8'h00;
            reg_file[14618] <= 8'h00;
            reg_file[14619] <= 8'h00;
            reg_file[14620] <= 8'h00;
            reg_file[14621] <= 8'h00;
            reg_file[14622] <= 8'h00;
            reg_file[14623] <= 8'h00;
            reg_file[14624] <= 8'h00;
            reg_file[14625] <= 8'h00;
            reg_file[14626] <= 8'h00;
            reg_file[14627] <= 8'h00;
            reg_file[14628] <= 8'h00;
            reg_file[14629] <= 8'h00;
            reg_file[14630] <= 8'h00;
            reg_file[14631] <= 8'h00;
            reg_file[14632] <= 8'h00;
            reg_file[14633] <= 8'h00;
            reg_file[14634] <= 8'h00;
            reg_file[14635] <= 8'h00;
            reg_file[14636] <= 8'h00;
            reg_file[14637] <= 8'h00;
            reg_file[14638] <= 8'h00;
            reg_file[14639] <= 8'h00;
            reg_file[14640] <= 8'h00;
            reg_file[14641] <= 8'h00;
            reg_file[14642] <= 8'h00;
            reg_file[14643] <= 8'h00;
            reg_file[14644] <= 8'h00;
            reg_file[14645] <= 8'h00;
            reg_file[14646] <= 8'h00;
            reg_file[14647] <= 8'h00;
            reg_file[14648] <= 8'h00;
            reg_file[14649] <= 8'h00;
            reg_file[14650] <= 8'h00;
            reg_file[14651] <= 8'h00;
            reg_file[14652] <= 8'h00;
            reg_file[14653] <= 8'h00;
            reg_file[14654] <= 8'h00;
            reg_file[14655] <= 8'h00;
            reg_file[14656] <= 8'h00;
            reg_file[14657] <= 8'h00;
            reg_file[14658] <= 8'h00;
            reg_file[14659] <= 8'h00;
            reg_file[14660] <= 8'h00;
            reg_file[14661] <= 8'h00;
            reg_file[14662] <= 8'h00;
            reg_file[14663] <= 8'h00;
            reg_file[14664] <= 8'h00;
            reg_file[14665] <= 8'h00;
            reg_file[14666] <= 8'h00;
            reg_file[14667] <= 8'h00;
            reg_file[14668] <= 8'h00;
            reg_file[14669] <= 8'h00;
            reg_file[14670] <= 8'h00;
            reg_file[14671] <= 8'h00;
            reg_file[14672] <= 8'h00;
            reg_file[14673] <= 8'h00;
            reg_file[14674] <= 8'h00;
            reg_file[14675] <= 8'h00;
            reg_file[14676] <= 8'h00;
            reg_file[14677] <= 8'h00;
            reg_file[14678] <= 8'h00;
            reg_file[14679] <= 8'h00;
            reg_file[14680] <= 8'h00;
            reg_file[14681] <= 8'h00;
            reg_file[14682] <= 8'h00;
            reg_file[14683] <= 8'h00;
            reg_file[14684] <= 8'h00;
            reg_file[14685] <= 8'h00;
            reg_file[14686] <= 8'h00;
            reg_file[14687] <= 8'h00;
            reg_file[14688] <= 8'h00;
            reg_file[14689] <= 8'h00;
            reg_file[14690] <= 8'h00;
            reg_file[14691] <= 8'h00;
            reg_file[14692] <= 8'h00;
            reg_file[14693] <= 8'h00;
            reg_file[14694] <= 8'h00;
            reg_file[14695] <= 8'h00;
            reg_file[14696] <= 8'h00;
            reg_file[14697] <= 8'h00;
            reg_file[14698] <= 8'h00;
            reg_file[14699] <= 8'h00;
            reg_file[14700] <= 8'h00;
            reg_file[14701] <= 8'h00;
            reg_file[14702] <= 8'h00;
            reg_file[14703] <= 8'h00;
            reg_file[14704] <= 8'h00;
            reg_file[14705] <= 8'h00;
            reg_file[14706] <= 8'h00;
            reg_file[14707] <= 8'h00;
            reg_file[14708] <= 8'h00;
            reg_file[14709] <= 8'h00;
            reg_file[14710] <= 8'h00;
            reg_file[14711] <= 8'h00;
            reg_file[14712] <= 8'h00;
            reg_file[14713] <= 8'h00;
            reg_file[14714] <= 8'h00;
            reg_file[14715] <= 8'h00;
            reg_file[14716] <= 8'h00;
            reg_file[14717] <= 8'h00;
            reg_file[14718] <= 8'h00;
            reg_file[14719] <= 8'h00;
            reg_file[14720] <= 8'h00;
            reg_file[14721] <= 8'h00;
            reg_file[14722] <= 8'h00;
            reg_file[14723] <= 8'h00;
            reg_file[14724] <= 8'h00;
            reg_file[14725] <= 8'h00;
            reg_file[14726] <= 8'h00;
            reg_file[14727] <= 8'h00;
            reg_file[14728] <= 8'h00;
            reg_file[14729] <= 8'h00;
            reg_file[14730] <= 8'h00;
            reg_file[14731] <= 8'h00;
            reg_file[14732] <= 8'h00;
            reg_file[14733] <= 8'h00;
            reg_file[14734] <= 8'h00;
            reg_file[14735] <= 8'h00;
            reg_file[14736] <= 8'h00;
            reg_file[14737] <= 8'h00;
            reg_file[14738] <= 8'h00;
            reg_file[14739] <= 8'h00;
            reg_file[14740] <= 8'h00;
            reg_file[14741] <= 8'h00;
            reg_file[14742] <= 8'h00;
            reg_file[14743] <= 8'h00;
            reg_file[14744] <= 8'h00;
            reg_file[14745] <= 8'h00;
            reg_file[14746] <= 8'h00;
            reg_file[14747] <= 8'h00;
            reg_file[14748] <= 8'h00;
            reg_file[14749] <= 8'h00;
            reg_file[14750] <= 8'h00;
            reg_file[14751] <= 8'h00;
            reg_file[14752] <= 8'h00;
            reg_file[14753] <= 8'h00;
            reg_file[14754] <= 8'h00;
            reg_file[14755] <= 8'h00;
            reg_file[14756] <= 8'h00;
            reg_file[14757] <= 8'h00;
            reg_file[14758] <= 8'h00;
            reg_file[14759] <= 8'h00;
            reg_file[14760] <= 8'h00;
            reg_file[14761] <= 8'h00;
            reg_file[14762] <= 8'h00;
            reg_file[14763] <= 8'h00;
            reg_file[14764] <= 8'h00;
            reg_file[14765] <= 8'h00;
            reg_file[14766] <= 8'h00;
            reg_file[14767] <= 8'h00;
            reg_file[14768] <= 8'h00;
            reg_file[14769] <= 8'h00;
            reg_file[14770] <= 8'h00;
            reg_file[14771] <= 8'h00;
            reg_file[14772] <= 8'h00;
            reg_file[14773] <= 8'h00;
            reg_file[14774] <= 8'h00;
            reg_file[14775] <= 8'h00;
            reg_file[14776] <= 8'h00;
            reg_file[14777] <= 8'h00;
            reg_file[14778] <= 8'h00;
            reg_file[14779] <= 8'h00;
            reg_file[14780] <= 8'h00;
            reg_file[14781] <= 8'h00;
            reg_file[14782] <= 8'h00;
            reg_file[14783] <= 8'h00;
            reg_file[14784] <= 8'h00;
            reg_file[14785] <= 8'h00;
            reg_file[14786] <= 8'h00;
            reg_file[14787] <= 8'h00;
            reg_file[14788] <= 8'h00;
            reg_file[14789] <= 8'h00;
            reg_file[14790] <= 8'h00;
            reg_file[14791] <= 8'h00;
            reg_file[14792] <= 8'h00;
            reg_file[14793] <= 8'h00;
            reg_file[14794] <= 8'h00;
            reg_file[14795] <= 8'h00;
            reg_file[14796] <= 8'h00;
            reg_file[14797] <= 8'h00;
            reg_file[14798] <= 8'h00;
            reg_file[14799] <= 8'h00;
            reg_file[14800] <= 8'h00;
            reg_file[14801] <= 8'h00;
            reg_file[14802] <= 8'h00;
            reg_file[14803] <= 8'h00;
            reg_file[14804] <= 8'h00;
            reg_file[14805] <= 8'h00;
            reg_file[14806] <= 8'h00;
            reg_file[14807] <= 8'h00;
            reg_file[14808] <= 8'h00;
            reg_file[14809] <= 8'h00;
            reg_file[14810] <= 8'h00;
            reg_file[14811] <= 8'h00;
            reg_file[14812] <= 8'h00;
            reg_file[14813] <= 8'h00;
            reg_file[14814] <= 8'h00;
            reg_file[14815] <= 8'h00;
            reg_file[14816] <= 8'h00;
            reg_file[14817] <= 8'h00;
            reg_file[14818] <= 8'h00;
            reg_file[14819] <= 8'h00;
            reg_file[14820] <= 8'h00;
            reg_file[14821] <= 8'h00;
            reg_file[14822] <= 8'h00;
            reg_file[14823] <= 8'h00;
            reg_file[14824] <= 8'h00;
            reg_file[14825] <= 8'h00;
            reg_file[14826] <= 8'h00;
            reg_file[14827] <= 8'h00;
            reg_file[14828] <= 8'h00;
            reg_file[14829] <= 8'h00;
            reg_file[14830] <= 8'h00;
            reg_file[14831] <= 8'h00;
            reg_file[14832] <= 8'h00;
            reg_file[14833] <= 8'h00;
            reg_file[14834] <= 8'h00;
            reg_file[14835] <= 8'h00;
            reg_file[14836] <= 8'h00;
            reg_file[14837] <= 8'h00;
            reg_file[14838] <= 8'h00;
            reg_file[14839] <= 8'h00;
            reg_file[14840] <= 8'h00;
            reg_file[14841] <= 8'h00;
            reg_file[14842] <= 8'h00;
            reg_file[14843] <= 8'h00;
            reg_file[14844] <= 8'h00;
            reg_file[14845] <= 8'h00;
            reg_file[14846] <= 8'h00;
            reg_file[14847] <= 8'h00;
            reg_file[14848] <= 8'h00;
            reg_file[14849] <= 8'h00;
            reg_file[14850] <= 8'h00;
            reg_file[14851] <= 8'h00;
            reg_file[14852] <= 8'h00;
            reg_file[14853] <= 8'h00;
            reg_file[14854] <= 8'h00;
            reg_file[14855] <= 8'h00;
            reg_file[14856] <= 8'h00;
            reg_file[14857] <= 8'h00;
            reg_file[14858] <= 8'h00;
            reg_file[14859] <= 8'h00;
            reg_file[14860] <= 8'h00;
            reg_file[14861] <= 8'h00;
            reg_file[14862] <= 8'h00;
            reg_file[14863] <= 8'h00;
            reg_file[14864] <= 8'h00;
            reg_file[14865] <= 8'h00;
            reg_file[14866] <= 8'h00;
            reg_file[14867] <= 8'h00;
            reg_file[14868] <= 8'h00;
            reg_file[14869] <= 8'h00;
            reg_file[14870] <= 8'h00;
            reg_file[14871] <= 8'h00;
            reg_file[14872] <= 8'h00;
            reg_file[14873] <= 8'h00;
            reg_file[14874] <= 8'h00;
            reg_file[14875] <= 8'h00;
            reg_file[14876] <= 8'h00;
            reg_file[14877] <= 8'h00;
            reg_file[14878] <= 8'h00;
            reg_file[14879] <= 8'h00;
            reg_file[14880] <= 8'h00;
            reg_file[14881] <= 8'h00;
            reg_file[14882] <= 8'h00;
            reg_file[14883] <= 8'h00;
            reg_file[14884] <= 8'h00;
            reg_file[14885] <= 8'h00;
            reg_file[14886] <= 8'h00;
            reg_file[14887] <= 8'h00;
            reg_file[14888] <= 8'h00;
            reg_file[14889] <= 8'h00;
            reg_file[14890] <= 8'h00;
            reg_file[14891] <= 8'h00;
            reg_file[14892] <= 8'h00;
            reg_file[14893] <= 8'h00;
            reg_file[14894] <= 8'h00;
            reg_file[14895] <= 8'h00;
            reg_file[14896] <= 8'h00;
            reg_file[14897] <= 8'h00;
            reg_file[14898] <= 8'h00;
            reg_file[14899] <= 8'h00;
            reg_file[14900] <= 8'h00;
            reg_file[14901] <= 8'h00;
            reg_file[14902] <= 8'h00;
            reg_file[14903] <= 8'h00;
            reg_file[14904] <= 8'h00;
            reg_file[14905] <= 8'h00;
            reg_file[14906] <= 8'h00;
            reg_file[14907] <= 8'h00;
            reg_file[14908] <= 8'h00;
            reg_file[14909] <= 8'h00;
            reg_file[14910] <= 8'h00;
            reg_file[14911] <= 8'h00;
            reg_file[14912] <= 8'h00;
            reg_file[14913] <= 8'h00;
            reg_file[14914] <= 8'h00;
            reg_file[14915] <= 8'h00;
            reg_file[14916] <= 8'h00;
            reg_file[14917] <= 8'h00;
            reg_file[14918] <= 8'h00;
            reg_file[14919] <= 8'h00;
            reg_file[14920] <= 8'h00;
            reg_file[14921] <= 8'h00;
            reg_file[14922] <= 8'h00;
            reg_file[14923] <= 8'h00;
            reg_file[14924] <= 8'h00;
            reg_file[14925] <= 8'h00;
            reg_file[14926] <= 8'h00;
            reg_file[14927] <= 8'h00;
            reg_file[14928] <= 8'h00;
            reg_file[14929] <= 8'h00;
            reg_file[14930] <= 8'h00;
            reg_file[14931] <= 8'h00;
            reg_file[14932] <= 8'h00;
            reg_file[14933] <= 8'h00;
            reg_file[14934] <= 8'h00;
            reg_file[14935] <= 8'h00;
            reg_file[14936] <= 8'h00;
            reg_file[14937] <= 8'h00;
            reg_file[14938] <= 8'h00;
            reg_file[14939] <= 8'h00;
            reg_file[14940] <= 8'h00;
            reg_file[14941] <= 8'h00;
            reg_file[14942] <= 8'h00;
            reg_file[14943] <= 8'h00;
            reg_file[14944] <= 8'h00;
            reg_file[14945] <= 8'h00;
            reg_file[14946] <= 8'h00;
            reg_file[14947] <= 8'h00;
            reg_file[14948] <= 8'h00;
            reg_file[14949] <= 8'h00;
            reg_file[14950] <= 8'h00;
            reg_file[14951] <= 8'h00;
            reg_file[14952] <= 8'h00;
            reg_file[14953] <= 8'h00;
            reg_file[14954] <= 8'h00;
            reg_file[14955] <= 8'h00;
            reg_file[14956] <= 8'h00;
            reg_file[14957] <= 8'h00;
            reg_file[14958] <= 8'h00;
            reg_file[14959] <= 8'h00;
            reg_file[14960] <= 8'h00;
            reg_file[14961] <= 8'h00;
            reg_file[14962] <= 8'h00;
            reg_file[14963] <= 8'h00;
            reg_file[14964] <= 8'h00;
            reg_file[14965] <= 8'h00;
            reg_file[14966] <= 8'h00;
            reg_file[14967] <= 8'h00;
            reg_file[14968] <= 8'h00;
            reg_file[14969] <= 8'h00;
            reg_file[14970] <= 8'h00;
            reg_file[14971] <= 8'h00;
            reg_file[14972] <= 8'h00;
            reg_file[14973] <= 8'h00;
            reg_file[14974] <= 8'h00;
            reg_file[14975] <= 8'h00;
            reg_file[14976] <= 8'h00;
            reg_file[14977] <= 8'h00;
            reg_file[14978] <= 8'h00;
            reg_file[14979] <= 8'h00;
            reg_file[14980] <= 8'h00;
            reg_file[14981] <= 8'h00;
            reg_file[14982] <= 8'h00;
            reg_file[14983] <= 8'h00;
            reg_file[14984] <= 8'h00;
            reg_file[14985] <= 8'h00;
            reg_file[14986] <= 8'h00;
            reg_file[14987] <= 8'h00;
            reg_file[14988] <= 8'h00;
            reg_file[14989] <= 8'h00;
            reg_file[14990] <= 8'h00;
            reg_file[14991] <= 8'h00;
            reg_file[14992] <= 8'h00;
            reg_file[14993] <= 8'h00;
            reg_file[14994] <= 8'h00;
            reg_file[14995] <= 8'h00;
            reg_file[14996] <= 8'h00;
            reg_file[14997] <= 8'h00;
            reg_file[14998] <= 8'h00;
            reg_file[14999] <= 8'h00;
            reg_file[15000] <= 8'h00;
            reg_file[15001] <= 8'h00;
            reg_file[15002] <= 8'h00;
            reg_file[15003] <= 8'h00;
            reg_file[15004] <= 8'h00;
            reg_file[15005] <= 8'h00;
            reg_file[15006] <= 8'h00;
            reg_file[15007] <= 8'h00;
            reg_file[15008] <= 8'h00;
            reg_file[15009] <= 8'h00;
            reg_file[15010] <= 8'h00;
            reg_file[15011] <= 8'h00;
            reg_file[15012] <= 8'h00;
            reg_file[15013] <= 8'h00;
            reg_file[15014] <= 8'h00;
            reg_file[15015] <= 8'h00;
            reg_file[15016] <= 8'h00;
            reg_file[15017] <= 8'h00;
            reg_file[15018] <= 8'h00;
            reg_file[15019] <= 8'h00;
            reg_file[15020] <= 8'h00;
            reg_file[15021] <= 8'h00;
            reg_file[15022] <= 8'h00;
            reg_file[15023] <= 8'h00;
            reg_file[15024] <= 8'h00;
            reg_file[15025] <= 8'h00;
            reg_file[15026] <= 8'h00;
            reg_file[15027] <= 8'h00;
            reg_file[15028] <= 8'h00;
            reg_file[15029] <= 8'h00;
            reg_file[15030] <= 8'h00;
            reg_file[15031] <= 8'h00;
            reg_file[15032] <= 8'h00;
            reg_file[15033] <= 8'h00;
            reg_file[15034] <= 8'h00;
            reg_file[15035] <= 8'h00;
            reg_file[15036] <= 8'h00;
            reg_file[15037] <= 8'h00;
            reg_file[15038] <= 8'h00;
            reg_file[15039] <= 8'h00;
            reg_file[15040] <= 8'h00;
            reg_file[15041] <= 8'h00;
            reg_file[15042] <= 8'h00;
            reg_file[15043] <= 8'h00;
            reg_file[15044] <= 8'h00;
            reg_file[15045] <= 8'h00;
            reg_file[15046] <= 8'h00;
            reg_file[15047] <= 8'h00;
            reg_file[15048] <= 8'h00;
            reg_file[15049] <= 8'h00;
            reg_file[15050] <= 8'h00;
            reg_file[15051] <= 8'h00;
            reg_file[15052] <= 8'h00;
            reg_file[15053] <= 8'h00;
            reg_file[15054] <= 8'h00;
            reg_file[15055] <= 8'h00;
            reg_file[15056] <= 8'h00;
            reg_file[15057] <= 8'h00;
            reg_file[15058] <= 8'h00;
            reg_file[15059] <= 8'h00;
            reg_file[15060] <= 8'h00;
            reg_file[15061] <= 8'h00;
            reg_file[15062] <= 8'h00;
            reg_file[15063] <= 8'h00;
            reg_file[15064] <= 8'h00;
            reg_file[15065] <= 8'h00;
            reg_file[15066] <= 8'h00;
            reg_file[15067] <= 8'h00;
            reg_file[15068] <= 8'h00;
            reg_file[15069] <= 8'h00;
            reg_file[15070] <= 8'h00;
            reg_file[15071] <= 8'h00;
            reg_file[15072] <= 8'h00;
            reg_file[15073] <= 8'h00;
            reg_file[15074] <= 8'h00;
            reg_file[15075] <= 8'h00;
            reg_file[15076] <= 8'h00;
            reg_file[15077] <= 8'h00;
            reg_file[15078] <= 8'h00;
            reg_file[15079] <= 8'h00;
            reg_file[15080] <= 8'h00;
            reg_file[15081] <= 8'h00;
            reg_file[15082] <= 8'h00;
            reg_file[15083] <= 8'h00;
            reg_file[15084] <= 8'h00;
            reg_file[15085] <= 8'h00;
            reg_file[15086] <= 8'h00;
            reg_file[15087] <= 8'h00;
            reg_file[15088] <= 8'h00;
            reg_file[15089] <= 8'h00;
            reg_file[15090] <= 8'h00;
            reg_file[15091] <= 8'h00;
            reg_file[15092] <= 8'h00;
            reg_file[15093] <= 8'h00;
            reg_file[15094] <= 8'h00;
            reg_file[15095] <= 8'h00;
            reg_file[15096] <= 8'h00;
            reg_file[15097] <= 8'h00;
            reg_file[15098] <= 8'h00;
            reg_file[15099] <= 8'h00;
            reg_file[15100] <= 8'h00;
            reg_file[15101] <= 8'h00;
            reg_file[15102] <= 8'h00;
            reg_file[15103] <= 8'h00;
            reg_file[15104] <= 8'h00;
            reg_file[15105] <= 8'h00;
            reg_file[15106] <= 8'h00;
            reg_file[15107] <= 8'h00;
            reg_file[15108] <= 8'h00;
            reg_file[15109] <= 8'h00;
            reg_file[15110] <= 8'h00;
            reg_file[15111] <= 8'h00;
            reg_file[15112] <= 8'h00;
            reg_file[15113] <= 8'h00;
            reg_file[15114] <= 8'h00;
            reg_file[15115] <= 8'h00;
            reg_file[15116] <= 8'h00;
            reg_file[15117] <= 8'h00;
            reg_file[15118] <= 8'h00;
            reg_file[15119] <= 8'h00;
            reg_file[15120] <= 8'h00;
            reg_file[15121] <= 8'h00;
            reg_file[15122] <= 8'h00;
            reg_file[15123] <= 8'h00;
            reg_file[15124] <= 8'h00;
            reg_file[15125] <= 8'h00;
            reg_file[15126] <= 8'h00;
            reg_file[15127] <= 8'h00;
            reg_file[15128] <= 8'h00;
            reg_file[15129] <= 8'h00;
            reg_file[15130] <= 8'h00;
            reg_file[15131] <= 8'h00;
            reg_file[15132] <= 8'h00;
            reg_file[15133] <= 8'h00;
            reg_file[15134] <= 8'h00;
            reg_file[15135] <= 8'h00;
            reg_file[15136] <= 8'h00;
            reg_file[15137] <= 8'h00;
            reg_file[15138] <= 8'h00;
            reg_file[15139] <= 8'h00;
            reg_file[15140] <= 8'h00;
            reg_file[15141] <= 8'h00;
            reg_file[15142] <= 8'h00;
            reg_file[15143] <= 8'h00;
            reg_file[15144] <= 8'h00;
            reg_file[15145] <= 8'h00;
            reg_file[15146] <= 8'h00;
            reg_file[15147] <= 8'h00;
            reg_file[15148] <= 8'h00;
            reg_file[15149] <= 8'h00;
            reg_file[15150] <= 8'h00;
            reg_file[15151] <= 8'h00;
            reg_file[15152] <= 8'h00;
            reg_file[15153] <= 8'h00;
            reg_file[15154] <= 8'h00;
            reg_file[15155] <= 8'h00;
            reg_file[15156] <= 8'h00;
            reg_file[15157] <= 8'h00;
            reg_file[15158] <= 8'h00;
            reg_file[15159] <= 8'h00;
            reg_file[15160] <= 8'h00;
            reg_file[15161] <= 8'h00;
            reg_file[15162] <= 8'h00;
            reg_file[15163] <= 8'h00;
            reg_file[15164] <= 8'h00;
            reg_file[15165] <= 8'h00;
            reg_file[15166] <= 8'h00;
            reg_file[15167] <= 8'h00;
            reg_file[15168] <= 8'h00;
            reg_file[15169] <= 8'h00;
            reg_file[15170] <= 8'h00;
            reg_file[15171] <= 8'h00;
            reg_file[15172] <= 8'h00;
            reg_file[15173] <= 8'h00;
            reg_file[15174] <= 8'h00;
            reg_file[15175] <= 8'h00;
            reg_file[15176] <= 8'h00;
            reg_file[15177] <= 8'h00;
            reg_file[15178] <= 8'h00;
            reg_file[15179] <= 8'h00;
            reg_file[15180] <= 8'h00;
            reg_file[15181] <= 8'h00;
            reg_file[15182] <= 8'h00;
            reg_file[15183] <= 8'h00;
            reg_file[15184] <= 8'h00;
            reg_file[15185] <= 8'h00;
            reg_file[15186] <= 8'h00;
            reg_file[15187] <= 8'h00;
            reg_file[15188] <= 8'h00;
            reg_file[15189] <= 8'h00;
            reg_file[15190] <= 8'h00;
            reg_file[15191] <= 8'h00;
            reg_file[15192] <= 8'h00;
            reg_file[15193] <= 8'h00;
            reg_file[15194] <= 8'h00;
            reg_file[15195] <= 8'h00;
            reg_file[15196] <= 8'h00;
            reg_file[15197] <= 8'h00;
            reg_file[15198] <= 8'h00;
            reg_file[15199] <= 8'h00;
            reg_file[15200] <= 8'h00;
            reg_file[15201] <= 8'h00;
            reg_file[15202] <= 8'h00;
            reg_file[15203] <= 8'h00;
            reg_file[15204] <= 8'h00;
            reg_file[15205] <= 8'h00;
            reg_file[15206] <= 8'h00;
            reg_file[15207] <= 8'h00;
            reg_file[15208] <= 8'h00;
            reg_file[15209] <= 8'h00;
            reg_file[15210] <= 8'h00;
            reg_file[15211] <= 8'h00;
            reg_file[15212] <= 8'h00;
            reg_file[15213] <= 8'h00;
            reg_file[15214] <= 8'h00;
            reg_file[15215] <= 8'h00;
            reg_file[15216] <= 8'h00;
            reg_file[15217] <= 8'h00;
            reg_file[15218] <= 8'h00;
            reg_file[15219] <= 8'h00;
            reg_file[15220] <= 8'h00;
            reg_file[15221] <= 8'h00;
            reg_file[15222] <= 8'h00;
            reg_file[15223] <= 8'h00;
            reg_file[15224] <= 8'h00;
            reg_file[15225] <= 8'h00;
            reg_file[15226] <= 8'h00;
            reg_file[15227] <= 8'h00;
            reg_file[15228] <= 8'h00;
            reg_file[15229] <= 8'h00;
            reg_file[15230] <= 8'h00;
            reg_file[15231] <= 8'h00;
            reg_file[15232] <= 8'h00;
            reg_file[15233] <= 8'h00;
            reg_file[15234] <= 8'h00;
            reg_file[15235] <= 8'h00;
            reg_file[15236] <= 8'h00;
            reg_file[15237] <= 8'h00;
            reg_file[15238] <= 8'h00;
            reg_file[15239] <= 8'h00;
            reg_file[15240] <= 8'h00;
            reg_file[15241] <= 8'h00;
            reg_file[15242] <= 8'h00;
            reg_file[15243] <= 8'h00;
            reg_file[15244] <= 8'h00;
            reg_file[15245] <= 8'h00;
            reg_file[15246] <= 8'h00;
            reg_file[15247] <= 8'h00;
            reg_file[15248] <= 8'h00;
            reg_file[15249] <= 8'h00;
            reg_file[15250] <= 8'h00;
            reg_file[15251] <= 8'h00;
            reg_file[15252] <= 8'h00;
            reg_file[15253] <= 8'h00;
            reg_file[15254] <= 8'h00;
            reg_file[15255] <= 8'h00;
            reg_file[15256] <= 8'h00;
            reg_file[15257] <= 8'h00;
            reg_file[15258] <= 8'h00;
            reg_file[15259] <= 8'h00;
            reg_file[15260] <= 8'h00;
            reg_file[15261] <= 8'h00;
            reg_file[15262] <= 8'h00;
            reg_file[15263] <= 8'h00;
            reg_file[15264] <= 8'h00;
            reg_file[15265] <= 8'h00;
            reg_file[15266] <= 8'h00;
            reg_file[15267] <= 8'h00;
            reg_file[15268] <= 8'h00;
            reg_file[15269] <= 8'h00;
            reg_file[15270] <= 8'h00;
            reg_file[15271] <= 8'h00;
            reg_file[15272] <= 8'h00;
            reg_file[15273] <= 8'h00;
            reg_file[15274] <= 8'h00;
            reg_file[15275] <= 8'h00;
            reg_file[15276] <= 8'h00;
            reg_file[15277] <= 8'h00;
            reg_file[15278] <= 8'h00;
            reg_file[15279] <= 8'h00;
            reg_file[15280] <= 8'h00;
            reg_file[15281] <= 8'h00;
            reg_file[15282] <= 8'h00;
            reg_file[15283] <= 8'h00;
            reg_file[15284] <= 8'h00;
            reg_file[15285] <= 8'h00;
            reg_file[15286] <= 8'h00;
            reg_file[15287] <= 8'h00;
            reg_file[15288] <= 8'h00;
            reg_file[15289] <= 8'h00;
            reg_file[15290] <= 8'h00;
            reg_file[15291] <= 8'h00;
            reg_file[15292] <= 8'h00;
            reg_file[15293] <= 8'h00;
            reg_file[15294] <= 8'h00;
            reg_file[15295] <= 8'h00;
            reg_file[15296] <= 8'h00;
            reg_file[15297] <= 8'h00;
            reg_file[15298] <= 8'h00;
            reg_file[15299] <= 8'h00;
            reg_file[15300] <= 8'h00;
            reg_file[15301] <= 8'h00;
            reg_file[15302] <= 8'h00;
            reg_file[15303] <= 8'h00;
            reg_file[15304] <= 8'h00;
            reg_file[15305] <= 8'h00;
            reg_file[15306] <= 8'h00;
            reg_file[15307] <= 8'h00;
            reg_file[15308] <= 8'h00;
            reg_file[15309] <= 8'h00;
            reg_file[15310] <= 8'h00;
            reg_file[15311] <= 8'h00;
            reg_file[15312] <= 8'h00;
            reg_file[15313] <= 8'h00;
            reg_file[15314] <= 8'h00;
            reg_file[15315] <= 8'h00;
            reg_file[15316] <= 8'h00;
            reg_file[15317] <= 8'h00;
            reg_file[15318] <= 8'h00;
            reg_file[15319] <= 8'h00;
            reg_file[15320] <= 8'h00;
            reg_file[15321] <= 8'h00;
            reg_file[15322] <= 8'h00;
            reg_file[15323] <= 8'h00;
            reg_file[15324] <= 8'h00;
            reg_file[15325] <= 8'h00;
            reg_file[15326] <= 8'h00;
            reg_file[15327] <= 8'h00;
            reg_file[15328] <= 8'h00;
            reg_file[15329] <= 8'h00;
            reg_file[15330] <= 8'h00;
            reg_file[15331] <= 8'h00;
            reg_file[15332] <= 8'h00;
            reg_file[15333] <= 8'h00;
            reg_file[15334] <= 8'h00;
            reg_file[15335] <= 8'h00;
            reg_file[15336] <= 8'h00;
            reg_file[15337] <= 8'h00;
            reg_file[15338] <= 8'h00;
            reg_file[15339] <= 8'h00;
            reg_file[15340] <= 8'h00;
            reg_file[15341] <= 8'h00;
            reg_file[15342] <= 8'h00;
            reg_file[15343] <= 8'h00;
            reg_file[15344] <= 8'h00;
            reg_file[15345] <= 8'h00;
            reg_file[15346] <= 8'h00;
            reg_file[15347] <= 8'h00;
            reg_file[15348] <= 8'h00;
            reg_file[15349] <= 8'h00;
            reg_file[15350] <= 8'h00;
            reg_file[15351] <= 8'h00;
            reg_file[15352] <= 8'h00;
            reg_file[15353] <= 8'h00;
            reg_file[15354] <= 8'h00;
            reg_file[15355] <= 8'h00;
            reg_file[15356] <= 8'h00;
            reg_file[15357] <= 8'h00;
            reg_file[15358] <= 8'h00;
            reg_file[15359] <= 8'h00;
            reg_file[15360] <= 8'h00;
            reg_file[15361] <= 8'h00;
            reg_file[15362] <= 8'h00;
            reg_file[15363] <= 8'h00;
            reg_file[15364] <= 8'h00;
            reg_file[15365] <= 8'h00;
            reg_file[15366] <= 8'h00;
            reg_file[15367] <= 8'h00;
            reg_file[15368] <= 8'h00;
            reg_file[15369] <= 8'h00;
            reg_file[15370] <= 8'h00;
            reg_file[15371] <= 8'h00;
            reg_file[15372] <= 8'h00;
            reg_file[15373] <= 8'h00;
            reg_file[15374] <= 8'h00;
            reg_file[15375] <= 8'h00;
            reg_file[15376] <= 8'h00;
            reg_file[15377] <= 8'h00;
            reg_file[15378] <= 8'h00;
            reg_file[15379] <= 8'h00;
            reg_file[15380] <= 8'h00;
            reg_file[15381] <= 8'h00;
            reg_file[15382] <= 8'h00;
            reg_file[15383] <= 8'h00;
            reg_file[15384] <= 8'h00;
            reg_file[15385] <= 8'h00;
            reg_file[15386] <= 8'h00;
            reg_file[15387] <= 8'h00;
            reg_file[15388] <= 8'h00;
            reg_file[15389] <= 8'h00;
            reg_file[15390] <= 8'h00;
            reg_file[15391] <= 8'h00;
            reg_file[15392] <= 8'h00;
            reg_file[15393] <= 8'h00;
            reg_file[15394] <= 8'h00;
            reg_file[15395] <= 8'h00;
            reg_file[15396] <= 8'h00;
            reg_file[15397] <= 8'h00;
            reg_file[15398] <= 8'h00;
            reg_file[15399] <= 8'h00;
            reg_file[15400] <= 8'h00;
            reg_file[15401] <= 8'h00;
            reg_file[15402] <= 8'h00;
            reg_file[15403] <= 8'h00;
            reg_file[15404] <= 8'h00;
            reg_file[15405] <= 8'h00;
            reg_file[15406] <= 8'h00;
            reg_file[15407] <= 8'h00;
            reg_file[15408] <= 8'h00;
            reg_file[15409] <= 8'h00;
            reg_file[15410] <= 8'h00;
            reg_file[15411] <= 8'h00;
            reg_file[15412] <= 8'h00;
            reg_file[15413] <= 8'h00;
            reg_file[15414] <= 8'h00;
            reg_file[15415] <= 8'h00;
            reg_file[15416] <= 8'h00;
            reg_file[15417] <= 8'h00;
            reg_file[15418] <= 8'h00;
            reg_file[15419] <= 8'h00;
            reg_file[15420] <= 8'h00;
            reg_file[15421] <= 8'h00;
            reg_file[15422] <= 8'h00;
            reg_file[15423] <= 8'h00;
            reg_file[15424] <= 8'h00;
            reg_file[15425] <= 8'h00;
            reg_file[15426] <= 8'h00;
            reg_file[15427] <= 8'h00;
            reg_file[15428] <= 8'h00;
            reg_file[15429] <= 8'h00;
            reg_file[15430] <= 8'h00;
            reg_file[15431] <= 8'h00;
            reg_file[15432] <= 8'h00;
            reg_file[15433] <= 8'h00;
            reg_file[15434] <= 8'h00;
            reg_file[15435] <= 8'h00;
            reg_file[15436] <= 8'h00;
            reg_file[15437] <= 8'h00;
            reg_file[15438] <= 8'h00;
            reg_file[15439] <= 8'h00;
            reg_file[15440] <= 8'h00;
            reg_file[15441] <= 8'h00;
            reg_file[15442] <= 8'h00;
            reg_file[15443] <= 8'h00;
            reg_file[15444] <= 8'h00;
            reg_file[15445] <= 8'h00;
            reg_file[15446] <= 8'h00;
            reg_file[15447] <= 8'h00;
            reg_file[15448] <= 8'h00;
            reg_file[15449] <= 8'h00;
            reg_file[15450] <= 8'h00;
            reg_file[15451] <= 8'h00;
            reg_file[15452] <= 8'h00;
            reg_file[15453] <= 8'h00;
            reg_file[15454] <= 8'h00;
            reg_file[15455] <= 8'h00;
            reg_file[15456] <= 8'h00;
            reg_file[15457] <= 8'h00;
            reg_file[15458] <= 8'h00;
            reg_file[15459] <= 8'h00;
            reg_file[15460] <= 8'h00;
            reg_file[15461] <= 8'h00;
            reg_file[15462] <= 8'h00;
            reg_file[15463] <= 8'h00;
            reg_file[15464] <= 8'h00;
            reg_file[15465] <= 8'h00;
            reg_file[15466] <= 8'h00;
            reg_file[15467] <= 8'h00;
            reg_file[15468] <= 8'h00;
            reg_file[15469] <= 8'h00;
            reg_file[15470] <= 8'h00;
            reg_file[15471] <= 8'h00;
            reg_file[15472] <= 8'h00;
            reg_file[15473] <= 8'h00;
            reg_file[15474] <= 8'h00;
            reg_file[15475] <= 8'h00;
            reg_file[15476] <= 8'h00;
            reg_file[15477] <= 8'h00;
            reg_file[15478] <= 8'h00;
            reg_file[15479] <= 8'h00;
            reg_file[15480] <= 8'h00;
            reg_file[15481] <= 8'h00;
            reg_file[15482] <= 8'h00;
            reg_file[15483] <= 8'h00;
            reg_file[15484] <= 8'h00;
            reg_file[15485] <= 8'h00;
            reg_file[15486] <= 8'h00;
            reg_file[15487] <= 8'h00;
            reg_file[15488] <= 8'h00;
            reg_file[15489] <= 8'h00;
            reg_file[15490] <= 8'h00;
            reg_file[15491] <= 8'h00;
            reg_file[15492] <= 8'h00;
            reg_file[15493] <= 8'h00;
            reg_file[15494] <= 8'h00;
            reg_file[15495] <= 8'h00;
            reg_file[15496] <= 8'h00;
            reg_file[15497] <= 8'h00;
            reg_file[15498] <= 8'h00;
            reg_file[15499] <= 8'h00;
            reg_file[15500] <= 8'h00;
            reg_file[15501] <= 8'h00;
            reg_file[15502] <= 8'h00;
            reg_file[15503] <= 8'h00;
            reg_file[15504] <= 8'h00;
            reg_file[15505] <= 8'h00;
            reg_file[15506] <= 8'h00;
            reg_file[15507] <= 8'h00;
            reg_file[15508] <= 8'h00;
            reg_file[15509] <= 8'h00;
            reg_file[15510] <= 8'h00;
            reg_file[15511] <= 8'h00;
            reg_file[15512] <= 8'h00;
            reg_file[15513] <= 8'h00;
            reg_file[15514] <= 8'h00;
            reg_file[15515] <= 8'h00;
            reg_file[15516] <= 8'h00;
            reg_file[15517] <= 8'h00;
            reg_file[15518] <= 8'h00;
            reg_file[15519] <= 8'h00;
            reg_file[15520] <= 8'h00;
            reg_file[15521] <= 8'h00;
            reg_file[15522] <= 8'h00;
            reg_file[15523] <= 8'h00;
            reg_file[15524] <= 8'h00;
            reg_file[15525] <= 8'h00;
            reg_file[15526] <= 8'h00;
            reg_file[15527] <= 8'h00;
            reg_file[15528] <= 8'h00;
            reg_file[15529] <= 8'h00;
            reg_file[15530] <= 8'h00;
            reg_file[15531] <= 8'h00;
            reg_file[15532] <= 8'h00;
            reg_file[15533] <= 8'h00;
            reg_file[15534] <= 8'h00;
            reg_file[15535] <= 8'h00;
            reg_file[15536] <= 8'h00;
            reg_file[15537] <= 8'h00;
            reg_file[15538] <= 8'h00;
            reg_file[15539] <= 8'h00;
            reg_file[15540] <= 8'h00;
            reg_file[15541] <= 8'h00;
            reg_file[15542] <= 8'h00;
            reg_file[15543] <= 8'h00;
            reg_file[15544] <= 8'h00;
            reg_file[15545] <= 8'h00;
            reg_file[15546] <= 8'h00;
            reg_file[15547] <= 8'h00;
            reg_file[15548] <= 8'h00;
            reg_file[15549] <= 8'h00;
            reg_file[15550] <= 8'h00;
            reg_file[15551] <= 8'h00;
            reg_file[15552] <= 8'h00;
            reg_file[15553] <= 8'h00;
            reg_file[15554] <= 8'h00;
            reg_file[15555] <= 8'h00;
            reg_file[15556] <= 8'h00;
            reg_file[15557] <= 8'h00;
            reg_file[15558] <= 8'h00;
            reg_file[15559] <= 8'h00;
            reg_file[15560] <= 8'h00;
            reg_file[15561] <= 8'h00;
            reg_file[15562] <= 8'h00;
            reg_file[15563] <= 8'h00;
            reg_file[15564] <= 8'h00;
            reg_file[15565] <= 8'h00;
            reg_file[15566] <= 8'h00;
            reg_file[15567] <= 8'h00;
            reg_file[15568] <= 8'h00;
            reg_file[15569] <= 8'h00;
            reg_file[15570] <= 8'h00;
            reg_file[15571] <= 8'h00;
            reg_file[15572] <= 8'h00;
            reg_file[15573] <= 8'h00;
            reg_file[15574] <= 8'h00;
            reg_file[15575] <= 8'h00;
            reg_file[15576] <= 8'h00;
            reg_file[15577] <= 8'h00;
            reg_file[15578] <= 8'h00;
            reg_file[15579] <= 8'h00;
            reg_file[15580] <= 8'h00;
            reg_file[15581] <= 8'h00;
            reg_file[15582] <= 8'h00;
            reg_file[15583] <= 8'h00;
            reg_file[15584] <= 8'h00;
            reg_file[15585] <= 8'h00;
            reg_file[15586] <= 8'h00;
            reg_file[15587] <= 8'h00;
            reg_file[15588] <= 8'h00;
            reg_file[15589] <= 8'h00;
            reg_file[15590] <= 8'h00;
            reg_file[15591] <= 8'h00;
            reg_file[15592] <= 8'h00;
            reg_file[15593] <= 8'h00;
            reg_file[15594] <= 8'h00;
            reg_file[15595] <= 8'h00;
            reg_file[15596] <= 8'h00;
            reg_file[15597] <= 8'h00;
            reg_file[15598] <= 8'h00;
            reg_file[15599] <= 8'h00;
            reg_file[15600] <= 8'h00;
            reg_file[15601] <= 8'h00;
            reg_file[15602] <= 8'h00;
            reg_file[15603] <= 8'h00;
            reg_file[15604] <= 8'h00;
            reg_file[15605] <= 8'h00;
            reg_file[15606] <= 8'h00;
            reg_file[15607] <= 8'h00;
            reg_file[15608] <= 8'h00;
            reg_file[15609] <= 8'h00;
            reg_file[15610] <= 8'h00;
            reg_file[15611] <= 8'h00;
            reg_file[15612] <= 8'h00;
            reg_file[15613] <= 8'h00;
            reg_file[15614] <= 8'h00;
            reg_file[15615] <= 8'h00;
            reg_file[15616] <= 8'h00;
            reg_file[15617] <= 8'h00;
            reg_file[15618] <= 8'h00;
            reg_file[15619] <= 8'h00;
            reg_file[15620] <= 8'h00;
            reg_file[15621] <= 8'h00;
            reg_file[15622] <= 8'h00;
            reg_file[15623] <= 8'h00;
            reg_file[15624] <= 8'h00;
            reg_file[15625] <= 8'h00;
            reg_file[15626] <= 8'h00;
            reg_file[15627] <= 8'h00;
            reg_file[15628] <= 8'h00;
            reg_file[15629] <= 8'h00;
            reg_file[15630] <= 8'h00;
            reg_file[15631] <= 8'h00;
            reg_file[15632] <= 8'h00;
            reg_file[15633] <= 8'h00;
            reg_file[15634] <= 8'h00;
            reg_file[15635] <= 8'h00;
            reg_file[15636] <= 8'h00;
            reg_file[15637] <= 8'h00;
            reg_file[15638] <= 8'h00;
            reg_file[15639] <= 8'h00;
            reg_file[15640] <= 8'h00;
            reg_file[15641] <= 8'h00;
            reg_file[15642] <= 8'h00;
            reg_file[15643] <= 8'h00;
            reg_file[15644] <= 8'h00;
            reg_file[15645] <= 8'h00;
            reg_file[15646] <= 8'h00;
            reg_file[15647] <= 8'h00;
            reg_file[15648] <= 8'h00;
            reg_file[15649] <= 8'h00;
            reg_file[15650] <= 8'h00;
            reg_file[15651] <= 8'h00;
            reg_file[15652] <= 8'h00;
            reg_file[15653] <= 8'h00;
            reg_file[15654] <= 8'h00;
            reg_file[15655] <= 8'h00;
            reg_file[15656] <= 8'h00;
            reg_file[15657] <= 8'h00;
            reg_file[15658] <= 8'h00;
            reg_file[15659] <= 8'h00;
            reg_file[15660] <= 8'h00;
            reg_file[15661] <= 8'h00;
            reg_file[15662] <= 8'h00;
            reg_file[15663] <= 8'h00;
            reg_file[15664] <= 8'h00;
            reg_file[15665] <= 8'h00;
            reg_file[15666] <= 8'h00;
            reg_file[15667] <= 8'h00;
            reg_file[15668] <= 8'h00;
            reg_file[15669] <= 8'h00;
            reg_file[15670] <= 8'h00;
            reg_file[15671] <= 8'h00;
            reg_file[15672] <= 8'h00;
            reg_file[15673] <= 8'h00;
            reg_file[15674] <= 8'h00;
            reg_file[15675] <= 8'h00;
            reg_file[15676] <= 8'h00;
            reg_file[15677] <= 8'h00;
            reg_file[15678] <= 8'h00;
            reg_file[15679] <= 8'h00;
            reg_file[15680] <= 8'h00;
            reg_file[15681] <= 8'h00;
            reg_file[15682] <= 8'h00;
            reg_file[15683] <= 8'h00;
            reg_file[15684] <= 8'h00;
            reg_file[15685] <= 8'h00;
            reg_file[15686] <= 8'h00;
            reg_file[15687] <= 8'h00;
            reg_file[15688] <= 8'h00;
            reg_file[15689] <= 8'h00;
            reg_file[15690] <= 8'h00;
            reg_file[15691] <= 8'h00;
            reg_file[15692] <= 8'h00;
            reg_file[15693] <= 8'h00;
            reg_file[15694] <= 8'h00;
            reg_file[15695] <= 8'h00;
            reg_file[15696] <= 8'h00;
            reg_file[15697] <= 8'h00;
            reg_file[15698] <= 8'h00;
            reg_file[15699] <= 8'h00;
            reg_file[15700] <= 8'h00;
            reg_file[15701] <= 8'h00;
            reg_file[15702] <= 8'h00;
            reg_file[15703] <= 8'h00;
            reg_file[15704] <= 8'h00;
            reg_file[15705] <= 8'h00;
            reg_file[15706] <= 8'h00;
            reg_file[15707] <= 8'h00;
            reg_file[15708] <= 8'h00;
            reg_file[15709] <= 8'h00;
            reg_file[15710] <= 8'h00;
            reg_file[15711] <= 8'h00;
            reg_file[15712] <= 8'h00;
            reg_file[15713] <= 8'h00;
            reg_file[15714] <= 8'h00;
            reg_file[15715] <= 8'h00;
            reg_file[15716] <= 8'h00;
            reg_file[15717] <= 8'h00;
            reg_file[15718] <= 8'h00;
            reg_file[15719] <= 8'h00;
            reg_file[15720] <= 8'h00;
            reg_file[15721] <= 8'h00;
            reg_file[15722] <= 8'h00;
            reg_file[15723] <= 8'h00;
            reg_file[15724] <= 8'h00;
            reg_file[15725] <= 8'h00;
            reg_file[15726] <= 8'h00;
            reg_file[15727] <= 8'h00;
            reg_file[15728] <= 8'h00;
            reg_file[15729] <= 8'h00;
            reg_file[15730] <= 8'h00;
            reg_file[15731] <= 8'h00;
            reg_file[15732] <= 8'h00;
            reg_file[15733] <= 8'h00;
            reg_file[15734] <= 8'h00;
            reg_file[15735] <= 8'h00;
            reg_file[15736] <= 8'h00;
            reg_file[15737] <= 8'h00;
            reg_file[15738] <= 8'h00;
            reg_file[15739] <= 8'h00;
            reg_file[15740] <= 8'h00;
            reg_file[15741] <= 8'h00;
            reg_file[15742] <= 8'h00;
            reg_file[15743] <= 8'h00;
            reg_file[15744] <= 8'h00;
            reg_file[15745] <= 8'h00;
            reg_file[15746] <= 8'h00;
            reg_file[15747] <= 8'h00;
            reg_file[15748] <= 8'h00;
            reg_file[15749] <= 8'h00;
            reg_file[15750] <= 8'h00;
            reg_file[15751] <= 8'h00;
            reg_file[15752] <= 8'h00;
            reg_file[15753] <= 8'h00;
            reg_file[15754] <= 8'h00;
            reg_file[15755] <= 8'h00;
            reg_file[15756] <= 8'h00;
            reg_file[15757] <= 8'h00;
            reg_file[15758] <= 8'h00;
            reg_file[15759] <= 8'h00;
            reg_file[15760] <= 8'h00;
            reg_file[15761] <= 8'h00;
            reg_file[15762] <= 8'h00;
            reg_file[15763] <= 8'h00;
            reg_file[15764] <= 8'h00;
            reg_file[15765] <= 8'h00;
            reg_file[15766] <= 8'h00;
            reg_file[15767] <= 8'h00;
            reg_file[15768] <= 8'h00;
            reg_file[15769] <= 8'h00;
            reg_file[15770] <= 8'h00;
            reg_file[15771] <= 8'h00;
            reg_file[15772] <= 8'h00;
            reg_file[15773] <= 8'h00;
            reg_file[15774] <= 8'h00;
            reg_file[15775] <= 8'h00;
            reg_file[15776] <= 8'h00;
            reg_file[15777] <= 8'h00;
            reg_file[15778] <= 8'h00;
            reg_file[15779] <= 8'h00;
            reg_file[15780] <= 8'h00;
            reg_file[15781] <= 8'h00;
            reg_file[15782] <= 8'h00;
            reg_file[15783] <= 8'h00;
            reg_file[15784] <= 8'h00;
            reg_file[15785] <= 8'h00;
            reg_file[15786] <= 8'h00;
            reg_file[15787] <= 8'h00;
            reg_file[15788] <= 8'h00;
            reg_file[15789] <= 8'h00;
            reg_file[15790] <= 8'h00;
            reg_file[15791] <= 8'h00;
            reg_file[15792] <= 8'h00;
            reg_file[15793] <= 8'h00;
            reg_file[15794] <= 8'h00;
            reg_file[15795] <= 8'h00;
            reg_file[15796] <= 8'h00;
            reg_file[15797] <= 8'h00;
            reg_file[15798] <= 8'h00;
            reg_file[15799] <= 8'h00;
            reg_file[15800] <= 8'h00;
            reg_file[15801] <= 8'h00;
            reg_file[15802] <= 8'h00;
            reg_file[15803] <= 8'h00;
            reg_file[15804] <= 8'h00;
            reg_file[15805] <= 8'h00;
            reg_file[15806] <= 8'h00;
            reg_file[15807] <= 8'h00;
            reg_file[15808] <= 8'h00;
            reg_file[15809] <= 8'h00;
            reg_file[15810] <= 8'h00;
            reg_file[15811] <= 8'h00;
            reg_file[15812] <= 8'h00;
            reg_file[15813] <= 8'h00;
            reg_file[15814] <= 8'h00;
            reg_file[15815] <= 8'h00;
            reg_file[15816] <= 8'h00;
            reg_file[15817] <= 8'h00;
            reg_file[15818] <= 8'h00;
            reg_file[15819] <= 8'h00;
            reg_file[15820] <= 8'h00;
            reg_file[15821] <= 8'h00;
            reg_file[15822] <= 8'h00;
            reg_file[15823] <= 8'h00;
            reg_file[15824] <= 8'h00;
            reg_file[15825] <= 8'h00;
            reg_file[15826] <= 8'h00;
            reg_file[15827] <= 8'h00;
            reg_file[15828] <= 8'h00;
            reg_file[15829] <= 8'h00;
            reg_file[15830] <= 8'h00;
            reg_file[15831] <= 8'h00;
            reg_file[15832] <= 8'h00;
            reg_file[15833] <= 8'h00;
            reg_file[15834] <= 8'h00;
            reg_file[15835] <= 8'h00;
            reg_file[15836] <= 8'h00;
            reg_file[15837] <= 8'h00;
            reg_file[15838] <= 8'h00;
            reg_file[15839] <= 8'h00;
            reg_file[15840] <= 8'h00;
            reg_file[15841] <= 8'h00;
            reg_file[15842] <= 8'h00;
            reg_file[15843] <= 8'h00;
            reg_file[15844] <= 8'h00;
            reg_file[15845] <= 8'h00;
            reg_file[15846] <= 8'h00;
            reg_file[15847] <= 8'h00;
            reg_file[15848] <= 8'h00;
            reg_file[15849] <= 8'h00;
            reg_file[15850] <= 8'h00;
            reg_file[15851] <= 8'h00;
            reg_file[15852] <= 8'h00;
            reg_file[15853] <= 8'h00;
            reg_file[15854] <= 8'h00;
            reg_file[15855] <= 8'h00;
            reg_file[15856] <= 8'h00;
            reg_file[15857] <= 8'h00;
            reg_file[15858] <= 8'h00;
            reg_file[15859] <= 8'h00;
            reg_file[15860] <= 8'h00;
            reg_file[15861] <= 8'h00;
            reg_file[15862] <= 8'h00;
            reg_file[15863] <= 8'h00;
            reg_file[15864] <= 8'h00;
            reg_file[15865] <= 8'h00;
            reg_file[15866] <= 8'h00;
            reg_file[15867] <= 8'h00;
            reg_file[15868] <= 8'h00;
            reg_file[15869] <= 8'h00;
            reg_file[15870] <= 8'h00;
            reg_file[15871] <= 8'h00;
            reg_file[15872] <= 8'h00;
            reg_file[15873] <= 8'h00;
            reg_file[15874] <= 8'h00;
            reg_file[15875] <= 8'h00;
            reg_file[15876] <= 8'h00;
            reg_file[15877] <= 8'h00;
            reg_file[15878] <= 8'h00;
            reg_file[15879] <= 8'h00;
            reg_file[15880] <= 8'h00;
            reg_file[15881] <= 8'h00;
            reg_file[15882] <= 8'h00;
            reg_file[15883] <= 8'h00;
            reg_file[15884] <= 8'h00;
            reg_file[15885] <= 8'h00;
            reg_file[15886] <= 8'h00;
            reg_file[15887] <= 8'h00;
            reg_file[15888] <= 8'h00;
            reg_file[15889] <= 8'h00;
            reg_file[15890] <= 8'h00;
            reg_file[15891] <= 8'h00;
            reg_file[15892] <= 8'h00;
            reg_file[15893] <= 8'h00;
            reg_file[15894] <= 8'h00;
            reg_file[15895] <= 8'h00;
            reg_file[15896] <= 8'h00;
            reg_file[15897] <= 8'h00;
            reg_file[15898] <= 8'h00;
            reg_file[15899] <= 8'h00;
            reg_file[15900] <= 8'h00;
            reg_file[15901] <= 8'h00;
            reg_file[15902] <= 8'h00;
            reg_file[15903] <= 8'h00;
            reg_file[15904] <= 8'h00;
            reg_file[15905] <= 8'h00;
            reg_file[15906] <= 8'h00;
            reg_file[15907] <= 8'h00;
            reg_file[15908] <= 8'h00;
            reg_file[15909] <= 8'h00;
            reg_file[15910] <= 8'h00;
            reg_file[15911] <= 8'h00;
            reg_file[15912] <= 8'h00;
            reg_file[15913] <= 8'h00;
            reg_file[15914] <= 8'h00;
            reg_file[15915] <= 8'h00;
            reg_file[15916] <= 8'h00;
            reg_file[15917] <= 8'h00;
            reg_file[15918] <= 8'h00;
            reg_file[15919] <= 8'h00;
            reg_file[15920] <= 8'h00;
            reg_file[15921] <= 8'h00;
            reg_file[15922] <= 8'h00;
            reg_file[15923] <= 8'h00;
            reg_file[15924] <= 8'h00;
            reg_file[15925] <= 8'h00;
            reg_file[15926] <= 8'h00;
            reg_file[15927] <= 8'h00;
            reg_file[15928] <= 8'h00;
            reg_file[15929] <= 8'h00;
            reg_file[15930] <= 8'h00;
            reg_file[15931] <= 8'h00;
            reg_file[15932] <= 8'h00;
            reg_file[15933] <= 8'h00;
            reg_file[15934] <= 8'h00;
            reg_file[15935] <= 8'h00;
            reg_file[15936] <= 8'h00;
            reg_file[15937] <= 8'h00;
            reg_file[15938] <= 8'h00;
            reg_file[15939] <= 8'h00;
            reg_file[15940] <= 8'h00;
            reg_file[15941] <= 8'h00;
            reg_file[15942] <= 8'h00;
            reg_file[15943] <= 8'h00;
            reg_file[15944] <= 8'h00;
            reg_file[15945] <= 8'h00;
            reg_file[15946] <= 8'h00;
            reg_file[15947] <= 8'h00;
            reg_file[15948] <= 8'h00;
            reg_file[15949] <= 8'h00;
            reg_file[15950] <= 8'h00;
            reg_file[15951] <= 8'h00;
            reg_file[15952] <= 8'h00;
            reg_file[15953] <= 8'h00;
            reg_file[15954] <= 8'h00;
            reg_file[15955] <= 8'h00;
            reg_file[15956] <= 8'h00;
            reg_file[15957] <= 8'h00;
            reg_file[15958] <= 8'h00;
            reg_file[15959] <= 8'h00;
            reg_file[15960] <= 8'h00;
            reg_file[15961] <= 8'h00;
            reg_file[15962] <= 8'h00;
            reg_file[15963] <= 8'h00;
            reg_file[15964] <= 8'h00;
            reg_file[15965] <= 8'h00;
            reg_file[15966] <= 8'h00;
            reg_file[15967] <= 8'h00;
            reg_file[15968] <= 8'h00;
            reg_file[15969] <= 8'h00;
            reg_file[15970] <= 8'h00;
            reg_file[15971] <= 8'h00;
            reg_file[15972] <= 8'h00;
            reg_file[15973] <= 8'h00;
            reg_file[15974] <= 8'h00;
            reg_file[15975] <= 8'h00;
            reg_file[15976] <= 8'h00;
            reg_file[15977] <= 8'h00;
            reg_file[15978] <= 8'h00;
            reg_file[15979] <= 8'h00;
            reg_file[15980] <= 8'h00;
            reg_file[15981] <= 8'h00;
            reg_file[15982] <= 8'h00;
            reg_file[15983] <= 8'h00;
            reg_file[15984] <= 8'h00;
            reg_file[15985] <= 8'h00;
            reg_file[15986] <= 8'h00;
            reg_file[15987] <= 8'h00;
            reg_file[15988] <= 8'h00;
            reg_file[15989] <= 8'h00;
            reg_file[15990] <= 8'h00;
            reg_file[15991] <= 8'h00;
            reg_file[15992] <= 8'h00;
            reg_file[15993] <= 8'h00;
            reg_file[15994] <= 8'h00;
            reg_file[15995] <= 8'h00;
            reg_file[15996] <= 8'h00;
            reg_file[15997] <= 8'h00;
            reg_file[15998] <= 8'h00;
            reg_file[15999] <= 8'h00;
            reg_file[16000] <= 8'h00;
            reg_file[16001] <= 8'h00;
            reg_file[16002] <= 8'h00;
            reg_file[16003] <= 8'h00;
            reg_file[16004] <= 8'h00;
            reg_file[16005] <= 8'h00;
            reg_file[16006] <= 8'h00;
            reg_file[16007] <= 8'h00;
            reg_file[16008] <= 8'h00;
            reg_file[16009] <= 8'h00;
            reg_file[16010] <= 8'h00;
            reg_file[16011] <= 8'h00;
            reg_file[16012] <= 8'h00;
            reg_file[16013] <= 8'h00;
            reg_file[16014] <= 8'h00;
            reg_file[16015] <= 8'h00;
            reg_file[16016] <= 8'h00;
            reg_file[16017] <= 8'h00;
            reg_file[16018] <= 8'h00;
            reg_file[16019] <= 8'h00;
            reg_file[16020] <= 8'h00;
            reg_file[16021] <= 8'h00;
            reg_file[16022] <= 8'h00;
            reg_file[16023] <= 8'h00;
            reg_file[16024] <= 8'h00;
            reg_file[16025] <= 8'h00;
            reg_file[16026] <= 8'h00;
            reg_file[16027] <= 8'h00;
            reg_file[16028] <= 8'h00;
            reg_file[16029] <= 8'h00;
            reg_file[16030] <= 8'h00;
            reg_file[16031] <= 8'h00;
            reg_file[16032] <= 8'h00;
            reg_file[16033] <= 8'h00;
            reg_file[16034] <= 8'h00;
            reg_file[16035] <= 8'h00;
            reg_file[16036] <= 8'h00;
            reg_file[16037] <= 8'h00;
            reg_file[16038] <= 8'h00;
            reg_file[16039] <= 8'h00;
            reg_file[16040] <= 8'h00;
            reg_file[16041] <= 8'h00;
            reg_file[16042] <= 8'h00;
            reg_file[16043] <= 8'h00;
            reg_file[16044] <= 8'h00;
            reg_file[16045] <= 8'h00;
            reg_file[16046] <= 8'h00;
            reg_file[16047] <= 8'h00;
            reg_file[16048] <= 8'h00;
            reg_file[16049] <= 8'h00;
            reg_file[16050] <= 8'h00;
            reg_file[16051] <= 8'h00;
            reg_file[16052] <= 8'h00;
            reg_file[16053] <= 8'h00;
            reg_file[16054] <= 8'h00;
            reg_file[16055] <= 8'h00;
            reg_file[16056] <= 8'h00;
            reg_file[16057] <= 8'h00;
            reg_file[16058] <= 8'h00;
            reg_file[16059] <= 8'h00;
            reg_file[16060] <= 8'h00;
            reg_file[16061] <= 8'h00;
            reg_file[16062] <= 8'h00;
            reg_file[16063] <= 8'h00;
            reg_file[16064] <= 8'h00;
            reg_file[16065] <= 8'h00;
            reg_file[16066] <= 8'h00;
            reg_file[16067] <= 8'h00;
            reg_file[16068] <= 8'h00;
            reg_file[16069] <= 8'h00;
            reg_file[16070] <= 8'h00;
            reg_file[16071] <= 8'h00;
            reg_file[16072] <= 8'h00;
            reg_file[16073] <= 8'h00;
            reg_file[16074] <= 8'h00;
            reg_file[16075] <= 8'h00;
            reg_file[16076] <= 8'h00;
            reg_file[16077] <= 8'h00;
            reg_file[16078] <= 8'h00;
            reg_file[16079] <= 8'h00;
            reg_file[16080] <= 8'h00;
            reg_file[16081] <= 8'h00;
            reg_file[16082] <= 8'h00;
            reg_file[16083] <= 8'h00;
            reg_file[16084] <= 8'h00;
            reg_file[16085] <= 8'h00;
            reg_file[16086] <= 8'h00;
            reg_file[16087] <= 8'h00;
            reg_file[16088] <= 8'h00;
            reg_file[16089] <= 8'h00;
            reg_file[16090] <= 8'h00;
            reg_file[16091] <= 8'h00;
            reg_file[16092] <= 8'h00;
            reg_file[16093] <= 8'h00;
            reg_file[16094] <= 8'h00;
            reg_file[16095] <= 8'h00;
            reg_file[16096] <= 8'h00;
            reg_file[16097] <= 8'h00;
            reg_file[16098] <= 8'h00;
            reg_file[16099] <= 8'h00;
            reg_file[16100] <= 8'h00;
            reg_file[16101] <= 8'h00;
            reg_file[16102] <= 8'h00;
            reg_file[16103] <= 8'h00;
            reg_file[16104] <= 8'h00;
            reg_file[16105] <= 8'h00;
            reg_file[16106] <= 8'h00;
            reg_file[16107] <= 8'h00;
            reg_file[16108] <= 8'h00;
            reg_file[16109] <= 8'h00;
            reg_file[16110] <= 8'h00;
            reg_file[16111] <= 8'h00;
            reg_file[16112] <= 8'h00;
            reg_file[16113] <= 8'h00;
            reg_file[16114] <= 8'h00;
            reg_file[16115] <= 8'h00;
            reg_file[16116] <= 8'h00;
            reg_file[16117] <= 8'h00;
            reg_file[16118] <= 8'h00;
            reg_file[16119] <= 8'h00;
            reg_file[16120] <= 8'h00;
            reg_file[16121] <= 8'h00;
            reg_file[16122] <= 8'h00;
            reg_file[16123] <= 8'h00;
            reg_file[16124] <= 8'h00;
            reg_file[16125] <= 8'h00;
            reg_file[16126] <= 8'h00;
            reg_file[16127] <= 8'h00;
            reg_file[16128] <= 8'h00;
            reg_file[16129] <= 8'h00;
            reg_file[16130] <= 8'h00;
            reg_file[16131] <= 8'h00;
            reg_file[16132] <= 8'h00;
            reg_file[16133] <= 8'h00;
            reg_file[16134] <= 8'h00;
            reg_file[16135] <= 8'h00;
            reg_file[16136] <= 8'h00;
            reg_file[16137] <= 8'h00;
            reg_file[16138] <= 8'h00;
            reg_file[16139] <= 8'h00;
            reg_file[16140] <= 8'h00;
            reg_file[16141] <= 8'h00;
            reg_file[16142] <= 8'h00;
            reg_file[16143] <= 8'h00;
            reg_file[16144] <= 8'h00;
            reg_file[16145] <= 8'h00;
            reg_file[16146] <= 8'h00;
            reg_file[16147] <= 8'h00;
            reg_file[16148] <= 8'h00;
            reg_file[16149] <= 8'h00;
            reg_file[16150] <= 8'h00;
            reg_file[16151] <= 8'h00;
            reg_file[16152] <= 8'h00;
            reg_file[16153] <= 8'h00;
            reg_file[16154] <= 8'h00;
            reg_file[16155] <= 8'h00;
            reg_file[16156] <= 8'h00;
            reg_file[16157] <= 8'h00;
            reg_file[16158] <= 8'h00;
            reg_file[16159] <= 8'h00;
            reg_file[16160] <= 8'h00;
            reg_file[16161] <= 8'h00;
            reg_file[16162] <= 8'h00;
            reg_file[16163] <= 8'h00;
            reg_file[16164] <= 8'h00;
            reg_file[16165] <= 8'h00;
            reg_file[16166] <= 8'h00;
            reg_file[16167] <= 8'h00;
            reg_file[16168] <= 8'h00;
            reg_file[16169] <= 8'h00;
            reg_file[16170] <= 8'h00;
            reg_file[16171] <= 8'h00;
            reg_file[16172] <= 8'h00;
            reg_file[16173] <= 8'h00;
            reg_file[16174] <= 8'h00;
            reg_file[16175] <= 8'h00;
            reg_file[16176] <= 8'h00;
            reg_file[16177] <= 8'h00;
            reg_file[16178] <= 8'h00;
            reg_file[16179] <= 8'h00;
            reg_file[16180] <= 8'h00;
            reg_file[16181] <= 8'h00;
            reg_file[16182] <= 8'h00;
            reg_file[16183] <= 8'h00;
            reg_file[16184] <= 8'h00;
            reg_file[16185] <= 8'h00;
            reg_file[16186] <= 8'h00;
            reg_file[16187] <= 8'h00;
            reg_file[16188] <= 8'h00;
            reg_file[16189] <= 8'h00;
            reg_file[16190] <= 8'h00;
            reg_file[16191] <= 8'h00;
            reg_file[16192] <= 8'h00;
            reg_file[16193] <= 8'h00;
            reg_file[16194] <= 8'h00;
            reg_file[16195] <= 8'h00;
            reg_file[16196] <= 8'h00;
            reg_file[16197] <= 8'h00;
            reg_file[16198] <= 8'h00;
            reg_file[16199] <= 8'h00;
            reg_file[16200] <= 8'h00;
            reg_file[16201] <= 8'h00;
            reg_file[16202] <= 8'h00;
            reg_file[16203] <= 8'h00;
            reg_file[16204] <= 8'h00;
            reg_file[16205] <= 8'h00;
            reg_file[16206] <= 8'h00;
            reg_file[16207] <= 8'h00;
            reg_file[16208] <= 8'h00;
            reg_file[16209] <= 8'h00;
            reg_file[16210] <= 8'h00;
            reg_file[16211] <= 8'h00;
            reg_file[16212] <= 8'h00;
            reg_file[16213] <= 8'h00;
            reg_file[16214] <= 8'h00;
            reg_file[16215] <= 8'h00;
            reg_file[16216] <= 8'h00;
            reg_file[16217] <= 8'h00;
            reg_file[16218] <= 8'h00;
            reg_file[16219] <= 8'h00;
            reg_file[16220] <= 8'h00;
            reg_file[16221] <= 8'h00;
            reg_file[16222] <= 8'h00;
            reg_file[16223] <= 8'h00;
            reg_file[16224] <= 8'h00;
            reg_file[16225] <= 8'h00;
            reg_file[16226] <= 8'h00;
            reg_file[16227] <= 8'h00;
            reg_file[16228] <= 8'h00;
            reg_file[16229] <= 8'h00;
            reg_file[16230] <= 8'h00;
            reg_file[16231] <= 8'h00;
            reg_file[16232] <= 8'h00;
            reg_file[16233] <= 8'h00;
            reg_file[16234] <= 8'h00;
            reg_file[16235] <= 8'h00;
            reg_file[16236] <= 8'h00;
            reg_file[16237] <= 8'h00;
            reg_file[16238] <= 8'h00;
            reg_file[16239] <= 8'h00;
            reg_file[16240] <= 8'h00;
            reg_file[16241] <= 8'h00;
            reg_file[16242] <= 8'h00;
            reg_file[16243] <= 8'h00;
            reg_file[16244] <= 8'h00;
            reg_file[16245] <= 8'h00;
            reg_file[16246] <= 8'h00;
            reg_file[16247] <= 8'h00;
            reg_file[16248] <= 8'h00;
            reg_file[16249] <= 8'h00;
            reg_file[16250] <= 8'h00;
            reg_file[16251] <= 8'h00;
            reg_file[16252] <= 8'h00;
            reg_file[16253] <= 8'h00;
            reg_file[16254] <= 8'h00;
            reg_file[16255] <= 8'h00;
            reg_file[16256] <= 8'h00;
            reg_file[16257] <= 8'h00;
            reg_file[16258] <= 8'h00;
            reg_file[16259] <= 8'h00;
            reg_file[16260] <= 8'h00;
            reg_file[16261] <= 8'h00;
            reg_file[16262] <= 8'h00;
            reg_file[16263] <= 8'h00;
            reg_file[16264] <= 8'h00;
            reg_file[16265] <= 8'h00;
            reg_file[16266] <= 8'h00;
            reg_file[16267] <= 8'h00;
            reg_file[16268] <= 8'h00;
            reg_file[16269] <= 8'h00;
            reg_file[16270] <= 8'h00;
            reg_file[16271] <= 8'h00;
            reg_file[16272] <= 8'h00;
            reg_file[16273] <= 8'h00;
            reg_file[16274] <= 8'h00;
            reg_file[16275] <= 8'h00;
            reg_file[16276] <= 8'h00;
            reg_file[16277] <= 8'h00;
            reg_file[16278] <= 8'h00;
            reg_file[16279] <= 8'h00;
            reg_file[16280] <= 8'h00;
            reg_file[16281] <= 8'h00;
            reg_file[16282] <= 8'h00;
            reg_file[16283] <= 8'h00;
            reg_file[16284] <= 8'h00;
            reg_file[16285] <= 8'h00;
            reg_file[16286] <= 8'h00;
            reg_file[16287] <= 8'h00;
            reg_file[16288] <= 8'h00;
            reg_file[16289] <= 8'h00;
            reg_file[16290] <= 8'h00;
            reg_file[16291] <= 8'h00;
            reg_file[16292] <= 8'h00;
            reg_file[16293] <= 8'h00;
            reg_file[16294] <= 8'h00;
            reg_file[16295] <= 8'h00;
            reg_file[16296] <= 8'h00;
            reg_file[16297] <= 8'h00;
            reg_file[16298] <= 8'h00;
            reg_file[16299] <= 8'h00;
            reg_file[16300] <= 8'h00;
            reg_file[16301] <= 8'h00;
            reg_file[16302] <= 8'h00;
            reg_file[16303] <= 8'h00;
            reg_file[16304] <= 8'h00;
            reg_file[16305] <= 8'h00;
            reg_file[16306] <= 8'h00;
            reg_file[16307] <= 8'h00;
            reg_file[16308] <= 8'h00;
            reg_file[16309] <= 8'h00;
            reg_file[16310] <= 8'h00;
            reg_file[16311] <= 8'h00;
            reg_file[16312] <= 8'h00;
            reg_file[16313] <= 8'h00;
            reg_file[16314] <= 8'h00;
            reg_file[16315] <= 8'h00;
            reg_file[16316] <= 8'h00;
            reg_file[16317] <= 8'h00;
            reg_file[16318] <= 8'h00;
            reg_file[16319] <= 8'h00;
            reg_file[16320] <= 8'h00;
            reg_file[16321] <= 8'h00;
            reg_file[16322] <= 8'h00;
            reg_file[16323] <= 8'h00;
            reg_file[16324] <= 8'h00;
            reg_file[16325] <= 8'h00;
            reg_file[16326] <= 8'h00;
            reg_file[16327] <= 8'h00;
            reg_file[16328] <= 8'h00;
            reg_file[16329] <= 8'h00;
            reg_file[16330] <= 8'h00;
            reg_file[16331] <= 8'h00;
            reg_file[16332] <= 8'h00;
            reg_file[16333] <= 8'h00;
            reg_file[16334] <= 8'h00;
            reg_file[16335] <= 8'h00;
            reg_file[16336] <= 8'h00;
            reg_file[16337] <= 8'h00;
            reg_file[16338] <= 8'h00;
            reg_file[16339] <= 8'h00;
            reg_file[16340] <= 8'h00;
            reg_file[16341] <= 8'h00;
            reg_file[16342] <= 8'h00;
            reg_file[16343] <= 8'h00;
            reg_file[16344] <= 8'h00;
            reg_file[16345] <= 8'h00;
            reg_file[16346] <= 8'h00;
            reg_file[16347] <= 8'h00;
            reg_file[16348] <= 8'h00;
            reg_file[16349] <= 8'h00;
            reg_file[16350] <= 8'h00;
            reg_file[16351] <= 8'h00;
            reg_file[16352] <= 8'h00;
            reg_file[16353] <= 8'h00;
            reg_file[16354] <= 8'h00;
            reg_file[16355] <= 8'h00;
            reg_file[16356] <= 8'h00;
            reg_file[16357] <= 8'h00;
            reg_file[16358] <= 8'h00;
            reg_file[16359] <= 8'h00;
            reg_file[16360] <= 8'h00;
            reg_file[16361] <= 8'h00;
            reg_file[16362] <= 8'h00;
            reg_file[16363] <= 8'h00;
            reg_file[16364] <= 8'h00;
            reg_file[16365] <= 8'h00;
            reg_file[16366] <= 8'h00;
            reg_file[16367] <= 8'h00;
            reg_file[16368] <= 8'h00;
            reg_file[16369] <= 8'h00;
            reg_file[16370] <= 8'h00;
            reg_file[16371] <= 8'h00;
            reg_file[16372] <= 8'h00;
            reg_file[16373] <= 8'h00;
            reg_file[16374] <= 8'h00;
            reg_file[16375] <= 8'h00;
            reg_file[16376] <= 8'h00;
            reg_file[16377] <= 8'h00;
            reg_file[16378] <= 8'h00;
            reg_file[16379] <= 8'h00;
            reg_file[16380] <= 8'h00;
            reg_file[16381] <= 8'h00;
            reg_file[16382] <= 8'h00;
            reg_file[16383] <= 8'h00;
            reg_file[16384] <= 8'h00;
            reg_file[16385] <= 8'h00;
            reg_file[16386] <= 8'h00;
            reg_file[16387] <= 8'h00;
            reg_file[16388] <= 8'h00;
            reg_file[16389] <= 8'h00;
            reg_file[16390] <= 8'h00;
            reg_file[16391] <= 8'h00;
            reg_file[16392] <= 8'h00;
            reg_file[16393] <= 8'h00;
            reg_file[16394] <= 8'h00;
            reg_file[16395] <= 8'h00;
            reg_file[16396] <= 8'h00;
            reg_file[16397] <= 8'h00;
            reg_file[16398] <= 8'h00;
            reg_file[16399] <= 8'h00;
            reg_file[16400] <= 8'h00;
            reg_file[16401] <= 8'h00;
            reg_file[16402] <= 8'h00;
            reg_file[16403] <= 8'h00;
            reg_file[16404] <= 8'h00;
            reg_file[16405] <= 8'h00;
            reg_file[16406] <= 8'h00;
            reg_file[16407] <= 8'h00;
            reg_file[16408] <= 8'h00;
            reg_file[16409] <= 8'h00;
            reg_file[16410] <= 8'h00;
            reg_file[16411] <= 8'h00;
            reg_file[16412] <= 8'h00;
            reg_file[16413] <= 8'h00;
            reg_file[16414] <= 8'h00;
            reg_file[16415] <= 8'h00;
            reg_file[16416] <= 8'h00;
            reg_file[16417] <= 8'h00;
            reg_file[16418] <= 8'h00;
            reg_file[16419] <= 8'h00;
            reg_file[16420] <= 8'h00;
            reg_file[16421] <= 8'h00;
            reg_file[16422] <= 8'h00;
            reg_file[16423] <= 8'h00;
            reg_file[16424] <= 8'h00;
            reg_file[16425] <= 8'h00;
            reg_file[16426] <= 8'h00;
            reg_file[16427] <= 8'h00;
            reg_file[16428] <= 8'h00;
            reg_file[16429] <= 8'h00;
            reg_file[16430] <= 8'h00;
            reg_file[16431] <= 8'h00;
            reg_file[16432] <= 8'h00;
            reg_file[16433] <= 8'h00;
            reg_file[16434] <= 8'h00;
            reg_file[16435] <= 8'h00;
            reg_file[16436] <= 8'h00;
            reg_file[16437] <= 8'h00;
            reg_file[16438] <= 8'h00;
            reg_file[16439] <= 8'h00;
            reg_file[16440] <= 8'h00;
            reg_file[16441] <= 8'h00;
            reg_file[16442] <= 8'h00;
            reg_file[16443] <= 8'h00;
            reg_file[16444] <= 8'h00;
            reg_file[16445] <= 8'h00;
            reg_file[16446] <= 8'h00;
            reg_file[16447] <= 8'h00;
            reg_file[16448] <= 8'h00;
            reg_file[16449] <= 8'h00;
            reg_file[16450] <= 8'h00;
            reg_file[16451] <= 8'h00;
            reg_file[16452] <= 8'h00;
            reg_file[16453] <= 8'h00;
            reg_file[16454] <= 8'h00;
            reg_file[16455] <= 8'h00;
            reg_file[16456] <= 8'h00;
            reg_file[16457] <= 8'h00;
            reg_file[16458] <= 8'h00;
            reg_file[16459] <= 8'h00;
            reg_file[16460] <= 8'h00;
            reg_file[16461] <= 8'h00;
            reg_file[16462] <= 8'h00;
            reg_file[16463] <= 8'h00;
            reg_file[16464] <= 8'h00;
            reg_file[16465] <= 8'h00;
            reg_file[16466] <= 8'h00;
            reg_file[16467] <= 8'h00;
            reg_file[16468] <= 8'h00;
            reg_file[16469] <= 8'h00;
            reg_file[16470] <= 8'h00;
            reg_file[16471] <= 8'h00;
            reg_file[16472] <= 8'h00;
            reg_file[16473] <= 8'h00;
            reg_file[16474] <= 8'h00;
            reg_file[16475] <= 8'h00;
            reg_file[16476] <= 8'h00;
            reg_file[16477] <= 8'h00;
            reg_file[16478] <= 8'h00;
            reg_file[16479] <= 8'h00;
            reg_file[16480] <= 8'h00;
            reg_file[16481] <= 8'h00;
            reg_file[16482] <= 8'h00;
            reg_file[16483] <= 8'h00;
            reg_file[16484] <= 8'h00;
            reg_file[16485] <= 8'h00;
            reg_file[16486] <= 8'h00;
            reg_file[16487] <= 8'h00;
            reg_file[16488] <= 8'h00;
            reg_file[16489] <= 8'h00;
            reg_file[16490] <= 8'h00;
            reg_file[16491] <= 8'h00;
            reg_file[16492] <= 8'h00;
            reg_file[16493] <= 8'h00;
            reg_file[16494] <= 8'h00;
            reg_file[16495] <= 8'h00;
            reg_file[16496] <= 8'h00;
            reg_file[16497] <= 8'h00;
            reg_file[16498] <= 8'h00;
            reg_file[16499] <= 8'h00;
            reg_file[16500] <= 8'h00;
            reg_file[16501] <= 8'h00;
            reg_file[16502] <= 8'h00;
            reg_file[16503] <= 8'h00;
            reg_file[16504] <= 8'h00;
            reg_file[16505] <= 8'h00;
            reg_file[16506] <= 8'h00;
            reg_file[16507] <= 8'h00;
            reg_file[16508] <= 8'h00;
            reg_file[16509] <= 8'h00;
            reg_file[16510] <= 8'h00;
            reg_file[16511] <= 8'h00;
            reg_file[16512] <= 8'h00;
            reg_file[16513] <= 8'h00;
            reg_file[16514] <= 8'h00;
            reg_file[16515] <= 8'h00;
            reg_file[16516] <= 8'h00;
            reg_file[16517] <= 8'h00;
            reg_file[16518] <= 8'h00;
            reg_file[16519] <= 8'h00;
            reg_file[16520] <= 8'h00;
            reg_file[16521] <= 8'h00;
            reg_file[16522] <= 8'h00;
            reg_file[16523] <= 8'h00;
            reg_file[16524] <= 8'h00;
            reg_file[16525] <= 8'h00;
            reg_file[16526] <= 8'h00;
            reg_file[16527] <= 8'h00;
            reg_file[16528] <= 8'h00;
            reg_file[16529] <= 8'h00;
            reg_file[16530] <= 8'h00;
            reg_file[16531] <= 8'h00;
            reg_file[16532] <= 8'h00;
            reg_file[16533] <= 8'h00;
            reg_file[16534] <= 8'h00;
            reg_file[16535] <= 8'h00;
            reg_file[16536] <= 8'h00;
            reg_file[16537] <= 8'h00;
            reg_file[16538] <= 8'h00;
            reg_file[16539] <= 8'h00;
            reg_file[16540] <= 8'h00;
            reg_file[16541] <= 8'h00;
            reg_file[16542] <= 8'h00;
            reg_file[16543] <= 8'h00;
            reg_file[16544] <= 8'h00;
            reg_file[16545] <= 8'h00;
            reg_file[16546] <= 8'h00;
            reg_file[16547] <= 8'h00;
            reg_file[16548] <= 8'h00;
            reg_file[16549] <= 8'h00;
            reg_file[16550] <= 8'h00;
            reg_file[16551] <= 8'h00;
            reg_file[16552] <= 8'h00;
            reg_file[16553] <= 8'h00;
            reg_file[16554] <= 8'h00;
            reg_file[16555] <= 8'h00;
            reg_file[16556] <= 8'h00;
            reg_file[16557] <= 8'h00;
            reg_file[16558] <= 8'h00;
            reg_file[16559] <= 8'h00;
            reg_file[16560] <= 8'h00;
            reg_file[16561] <= 8'h00;
            reg_file[16562] <= 8'h00;
            reg_file[16563] <= 8'h00;
            reg_file[16564] <= 8'h00;
            reg_file[16565] <= 8'h00;
            reg_file[16566] <= 8'h00;
            reg_file[16567] <= 8'h00;
            reg_file[16568] <= 8'h00;
            reg_file[16569] <= 8'h00;
            reg_file[16570] <= 8'h00;
            reg_file[16571] <= 8'h00;
            reg_file[16572] <= 8'h00;
            reg_file[16573] <= 8'h00;
            reg_file[16574] <= 8'h00;
            reg_file[16575] <= 8'h00;
            reg_file[16576] <= 8'h00;
            reg_file[16577] <= 8'h00;
            reg_file[16578] <= 8'h00;
            reg_file[16579] <= 8'h00;
            reg_file[16580] <= 8'h00;
            reg_file[16581] <= 8'h00;
            reg_file[16582] <= 8'h00;
            reg_file[16583] <= 8'h00;
            reg_file[16584] <= 8'h00;
            reg_file[16585] <= 8'h00;
            reg_file[16586] <= 8'h00;
            reg_file[16587] <= 8'h00;
            reg_file[16588] <= 8'h00;
            reg_file[16589] <= 8'h00;
            reg_file[16590] <= 8'h00;
            reg_file[16591] <= 8'h00;
            reg_file[16592] <= 8'h00;
            reg_file[16593] <= 8'h00;
            reg_file[16594] <= 8'h00;
            reg_file[16595] <= 8'h00;
            reg_file[16596] <= 8'h00;
            reg_file[16597] <= 8'h00;
            reg_file[16598] <= 8'h00;
            reg_file[16599] <= 8'h00;
            reg_file[16600] <= 8'h00;
            reg_file[16601] <= 8'h00;
            reg_file[16602] <= 8'h00;
            reg_file[16603] <= 8'h00;
            reg_file[16604] <= 8'h00;
            reg_file[16605] <= 8'h00;
            reg_file[16606] <= 8'h00;
            reg_file[16607] <= 8'h00;
            reg_file[16608] <= 8'h00;
            reg_file[16609] <= 8'h00;
            reg_file[16610] <= 8'h00;
            reg_file[16611] <= 8'h00;
            reg_file[16612] <= 8'h00;
            reg_file[16613] <= 8'h00;
            reg_file[16614] <= 8'h00;
            reg_file[16615] <= 8'h00;
            reg_file[16616] <= 8'h00;
            reg_file[16617] <= 8'h00;
            reg_file[16618] <= 8'h00;
            reg_file[16619] <= 8'h00;
            reg_file[16620] <= 8'h00;
            reg_file[16621] <= 8'h00;
            reg_file[16622] <= 8'h00;
            reg_file[16623] <= 8'h00;
            reg_file[16624] <= 8'h00;
            reg_file[16625] <= 8'h00;
            reg_file[16626] <= 8'h00;
            reg_file[16627] <= 8'h00;
            reg_file[16628] <= 8'h00;
            reg_file[16629] <= 8'h00;
            reg_file[16630] <= 8'h00;
            reg_file[16631] <= 8'h00;
            reg_file[16632] <= 8'h00;
            reg_file[16633] <= 8'h00;
            reg_file[16634] <= 8'h00;
            reg_file[16635] <= 8'h00;
            reg_file[16636] <= 8'h00;
            reg_file[16637] <= 8'h00;
            reg_file[16638] <= 8'h00;
            reg_file[16639] <= 8'h00;
            reg_file[16640] <= 8'h00;
            reg_file[16641] <= 8'h00;
            reg_file[16642] <= 8'h00;
            reg_file[16643] <= 8'h00;
            reg_file[16644] <= 8'h00;
            reg_file[16645] <= 8'h00;
            reg_file[16646] <= 8'h00;
            reg_file[16647] <= 8'h00;
            reg_file[16648] <= 8'h00;
            reg_file[16649] <= 8'h00;
            reg_file[16650] <= 8'h00;
            reg_file[16651] <= 8'h00;
            reg_file[16652] <= 8'h00;
            reg_file[16653] <= 8'h00;
            reg_file[16654] <= 8'h00;
            reg_file[16655] <= 8'h00;
            reg_file[16656] <= 8'h00;
            reg_file[16657] <= 8'h00;
            reg_file[16658] <= 8'h00;
            reg_file[16659] <= 8'h00;
            reg_file[16660] <= 8'h00;
            reg_file[16661] <= 8'h00;
            reg_file[16662] <= 8'h00;
            reg_file[16663] <= 8'h00;
            reg_file[16664] <= 8'h00;
            reg_file[16665] <= 8'h00;
            reg_file[16666] <= 8'h00;
            reg_file[16667] <= 8'h00;
            reg_file[16668] <= 8'h00;
            reg_file[16669] <= 8'h00;
            reg_file[16670] <= 8'h00;
            reg_file[16671] <= 8'h00;
            reg_file[16672] <= 8'h00;
            reg_file[16673] <= 8'h00;
            reg_file[16674] <= 8'h00;
            reg_file[16675] <= 8'h00;
            reg_file[16676] <= 8'h00;
            reg_file[16677] <= 8'h00;
            reg_file[16678] <= 8'h00;
            reg_file[16679] <= 8'h00;
            reg_file[16680] <= 8'h00;
            reg_file[16681] <= 8'h00;
            reg_file[16682] <= 8'h00;
            reg_file[16683] <= 8'h00;
            reg_file[16684] <= 8'h00;
            reg_file[16685] <= 8'h00;
            reg_file[16686] <= 8'h00;
            reg_file[16687] <= 8'h00;
            reg_file[16688] <= 8'h00;
            reg_file[16689] <= 8'h00;
            reg_file[16690] <= 8'h00;
            reg_file[16691] <= 8'h00;
            reg_file[16692] <= 8'h00;
            reg_file[16693] <= 8'h00;
            reg_file[16694] <= 8'h00;
            reg_file[16695] <= 8'h00;
            reg_file[16696] <= 8'h00;
            reg_file[16697] <= 8'h00;
            reg_file[16698] <= 8'h00;
            reg_file[16699] <= 8'h00;
            reg_file[16700] <= 8'h00;
            reg_file[16701] <= 8'h00;
            reg_file[16702] <= 8'h00;
            reg_file[16703] <= 8'h00;
            reg_file[16704] <= 8'h00;
            reg_file[16705] <= 8'h00;
            reg_file[16706] <= 8'h00;
            reg_file[16707] <= 8'h00;
            reg_file[16708] <= 8'h00;
            reg_file[16709] <= 8'h00;
            reg_file[16710] <= 8'h00;
            reg_file[16711] <= 8'h00;
            reg_file[16712] <= 8'h00;
            reg_file[16713] <= 8'h00;
            reg_file[16714] <= 8'h00;
            reg_file[16715] <= 8'h00;
            reg_file[16716] <= 8'h00;
            reg_file[16717] <= 8'h00;
            reg_file[16718] <= 8'h00;
            reg_file[16719] <= 8'h00;
            reg_file[16720] <= 8'h00;
            reg_file[16721] <= 8'h00;
            reg_file[16722] <= 8'h00;
            reg_file[16723] <= 8'h00;
            reg_file[16724] <= 8'h00;
            reg_file[16725] <= 8'h00;
            reg_file[16726] <= 8'h00;
            reg_file[16727] <= 8'h00;
            reg_file[16728] <= 8'h00;
            reg_file[16729] <= 8'h00;
            reg_file[16730] <= 8'h00;
            reg_file[16731] <= 8'h00;
            reg_file[16732] <= 8'h00;
            reg_file[16733] <= 8'h00;
            reg_file[16734] <= 8'h00;
            reg_file[16735] <= 8'h00;
            reg_file[16736] <= 8'h00;
            reg_file[16737] <= 8'h00;
            reg_file[16738] <= 8'h00;
            reg_file[16739] <= 8'h00;
            reg_file[16740] <= 8'h00;
            reg_file[16741] <= 8'h00;
            reg_file[16742] <= 8'h00;
            reg_file[16743] <= 8'h00;
            reg_file[16744] <= 8'h00;
            reg_file[16745] <= 8'h00;
            reg_file[16746] <= 8'h00;
            reg_file[16747] <= 8'h00;
            reg_file[16748] <= 8'h00;
            reg_file[16749] <= 8'h00;
            reg_file[16750] <= 8'h00;
            reg_file[16751] <= 8'h00;
            reg_file[16752] <= 8'h00;
            reg_file[16753] <= 8'h00;
            reg_file[16754] <= 8'h00;
            reg_file[16755] <= 8'h00;
            reg_file[16756] <= 8'h00;
            reg_file[16757] <= 8'h00;
            reg_file[16758] <= 8'h00;
            reg_file[16759] <= 8'h00;
            reg_file[16760] <= 8'h00;
            reg_file[16761] <= 8'h00;
            reg_file[16762] <= 8'h00;
            reg_file[16763] <= 8'h00;
            reg_file[16764] <= 8'h00;
            reg_file[16765] <= 8'h00;
            reg_file[16766] <= 8'h00;
            reg_file[16767] <= 8'h00;
            reg_file[16768] <= 8'h00;
            reg_file[16769] <= 8'h00;
            reg_file[16770] <= 8'h00;
            reg_file[16771] <= 8'h00;
            reg_file[16772] <= 8'h00;
            reg_file[16773] <= 8'h00;
            reg_file[16774] <= 8'h00;
            reg_file[16775] <= 8'h00;
            reg_file[16776] <= 8'h00;
            reg_file[16777] <= 8'h00;
            reg_file[16778] <= 8'h00;
            reg_file[16779] <= 8'h00;
            reg_file[16780] <= 8'h00;
            reg_file[16781] <= 8'h00;
            reg_file[16782] <= 8'h00;
            reg_file[16783] <= 8'h00;
            reg_file[16784] <= 8'h00;
            reg_file[16785] <= 8'h00;
            reg_file[16786] <= 8'h00;
            reg_file[16787] <= 8'h00;
            reg_file[16788] <= 8'h00;
            reg_file[16789] <= 8'h00;
            reg_file[16790] <= 8'h00;
            reg_file[16791] <= 8'h00;
            reg_file[16792] <= 8'h00;
            reg_file[16793] <= 8'h00;
            reg_file[16794] <= 8'h00;
            reg_file[16795] <= 8'h00;
            reg_file[16796] <= 8'h00;
            reg_file[16797] <= 8'h00;
            reg_file[16798] <= 8'h00;
            reg_file[16799] <= 8'h00;
            reg_file[16800] <= 8'h00;
            reg_file[16801] <= 8'h00;
            reg_file[16802] <= 8'h00;
            reg_file[16803] <= 8'h00;
            reg_file[16804] <= 8'h00;
            reg_file[16805] <= 8'h00;
            reg_file[16806] <= 8'h00;
            reg_file[16807] <= 8'h00;
            reg_file[16808] <= 8'h00;
            reg_file[16809] <= 8'h00;
            reg_file[16810] <= 8'h00;
            reg_file[16811] <= 8'h00;
            reg_file[16812] <= 8'h00;
            reg_file[16813] <= 8'h00;
            reg_file[16814] <= 8'h00;
            reg_file[16815] <= 8'h00;
            reg_file[16816] <= 8'h00;
            reg_file[16817] <= 8'h00;
            reg_file[16818] <= 8'h00;
            reg_file[16819] <= 8'h00;
            reg_file[16820] <= 8'h00;
            reg_file[16821] <= 8'h00;
            reg_file[16822] <= 8'h00;
            reg_file[16823] <= 8'h00;
            reg_file[16824] <= 8'h00;
            reg_file[16825] <= 8'h00;
            reg_file[16826] <= 8'h00;
            reg_file[16827] <= 8'h00;
            reg_file[16828] <= 8'h00;
            reg_file[16829] <= 8'h00;
            reg_file[16830] <= 8'h00;
            reg_file[16831] <= 8'h00;
            reg_file[16832] <= 8'h00;
            reg_file[16833] <= 8'h00;
            reg_file[16834] <= 8'h00;
            reg_file[16835] <= 8'h00;
            reg_file[16836] <= 8'h00;
            reg_file[16837] <= 8'h00;
            reg_file[16838] <= 8'h00;
            reg_file[16839] <= 8'h00;
            reg_file[16840] <= 8'h00;
            reg_file[16841] <= 8'h00;
            reg_file[16842] <= 8'h00;
            reg_file[16843] <= 8'h00;
            reg_file[16844] <= 8'h00;
            reg_file[16845] <= 8'h00;
            reg_file[16846] <= 8'h00;
            reg_file[16847] <= 8'h00;
            reg_file[16848] <= 8'h00;
            reg_file[16849] <= 8'h00;
            reg_file[16850] <= 8'h00;
            reg_file[16851] <= 8'h00;
            reg_file[16852] <= 8'h00;
            reg_file[16853] <= 8'h00;
            reg_file[16854] <= 8'h00;
            reg_file[16855] <= 8'h00;
            reg_file[16856] <= 8'h00;
            reg_file[16857] <= 8'h00;
            reg_file[16858] <= 8'h00;
            reg_file[16859] <= 8'h00;
            reg_file[16860] <= 8'h00;
            reg_file[16861] <= 8'h00;
            reg_file[16862] <= 8'h00;
            reg_file[16863] <= 8'h00;
            reg_file[16864] <= 8'h00;
            reg_file[16865] <= 8'h00;
            reg_file[16866] <= 8'h00;
            reg_file[16867] <= 8'h00;
            reg_file[16868] <= 8'h00;
            reg_file[16869] <= 8'h00;
            reg_file[16870] <= 8'h00;
            reg_file[16871] <= 8'h00;
            reg_file[16872] <= 8'h00;
            reg_file[16873] <= 8'h00;
            reg_file[16874] <= 8'h00;
            reg_file[16875] <= 8'h00;
            reg_file[16876] <= 8'h00;
            reg_file[16877] <= 8'h00;
            reg_file[16878] <= 8'h00;
            reg_file[16879] <= 8'h00;
            reg_file[16880] <= 8'h00;
            reg_file[16881] <= 8'h00;
            reg_file[16882] <= 8'h00;
            reg_file[16883] <= 8'h00;
            reg_file[16884] <= 8'h00;
            reg_file[16885] <= 8'h00;
            reg_file[16886] <= 8'h00;
            reg_file[16887] <= 8'h00;
            reg_file[16888] <= 8'h00;
            reg_file[16889] <= 8'h00;
            reg_file[16890] <= 8'h00;
            reg_file[16891] <= 8'h00;
            reg_file[16892] <= 8'h00;
            reg_file[16893] <= 8'h00;
            reg_file[16894] <= 8'h00;
            reg_file[16895] <= 8'h00;
            reg_file[16896] <= 8'h00;
            reg_file[16897] <= 8'h00;
            reg_file[16898] <= 8'h00;
            reg_file[16899] <= 8'h00;
            reg_file[16900] <= 8'h00;
            reg_file[16901] <= 8'h00;
            reg_file[16902] <= 8'h00;
            reg_file[16903] <= 8'h00;
            reg_file[16904] <= 8'h00;
            reg_file[16905] <= 8'h00;
            reg_file[16906] <= 8'h00;
            reg_file[16907] <= 8'h00;
            reg_file[16908] <= 8'h00;
            reg_file[16909] <= 8'h00;
            reg_file[16910] <= 8'h00;
            reg_file[16911] <= 8'h00;
            reg_file[16912] <= 8'h00;
            reg_file[16913] <= 8'h00;
            reg_file[16914] <= 8'h00;
            reg_file[16915] <= 8'h00;
            reg_file[16916] <= 8'h00;
            reg_file[16917] <= 8'h00;
            reg_file[16918] <= 8'h00;
            reg_file[16919] <= 8'h00;
            reg_file[16920] <= 8'h00;
            reg_file[16921] <= 8'h00;
            reg_file[16922] <= 8'h00;
            reg_file[16923] <= 8'h00;
            reg_file[16924] <= 8'h00;
            reg_file[16925] <= 8'h00;
            reg_file[16926] <= 8'h00;
            reg_file[16927] <= 8'h00;
            reg_file[16928] <= 8'h00;
            reg_file[16929] <= 8'h00;
            reg_file[16930] <= 8'h00;
            reg_file[16931] <= 8'h00;
            reg_file[16932] <= 8'h00;
            reg_file[16933] <= 8'h00;
            reg_file[16934] <= 8'h00;
            reg_file[16935] <= 8'h00;
            reg_file[16936] <= 8'h00;
            reg_file[16937] <= 8'h00;
            reg_file[16938] <= 8'h00;
            reg_file[16939] <= 8'h00;
            reg_file[16940] <= 8'h00;
            reg_file[16941] <= 8'h00;
            reg_file[16942] <= 8'h00;
            reg_file[16943] <= 8'h00;
            reg_file[16944] <= 8'h00;
            reg_file[16945] <= 8'h00;
            reg_file[16946] <= 8'h00;
            reg_file[16947] <= 8'h00;
            reg_file[16948] <= 8'h00;
            reg_file[16949] <= 8'h00;
            reg_file[16950] <= 8'h00;
            reg_file[16951] <= 8'h00;
            reg_file[16952] <= 8'h00;
            reg_file[16953] <= 8'h00;
            reg_file[16954] <= 8'h00;
            reg_file[16955] <= 8'h00;
            reg_file[16956] <= 8'h00;
            reg_file[16957] <= 8'h00;
            reg_file[16958] <= 8'h00;
            reg_file[16959] <= 8'h00;
            reg_file[16960] <= 8'h00;
            reg_file[16961] <= 8'h00;
            reg_file[16962] <= 8'h00;
            reg_file[16963] <= 8'h00;
            reg_file[16964] <= 8'h00;
            reg_file[16965] <= 8'h00;
            reg_file[16966] <= 8'h00;
            reg_file[16967] <= 8'h00;
            reg_file[16968] <= 8'h00;
            reg_file[16969] <= 8'h00;
            reg_file[16970] <= 8'h00;
            reg_file[16971] <= 8'h00;
            reg_file[16972] <= 8'h00;
            reg_file[16973] <= 8'h00;
            reg_file[16974] <= 8'h00;
            reg_file[16975] <= 8'h00;
            reg_file[16976] <= 8'h00;
            reg_file[16977] <= 8'h00;
            reg_file[16978] <= 8'h00;
            reg_file[16979] <= 8'h00;
            reg_file[16980] <= 8'h00;
            reg_file[16981] <= 8'h00;
            reg_file[16982] <= 8'h00;
            reg_file[16983] <= 8'h00;
            reg_file[16984] <= 8'h00;
            reg_file[16985] <= 8'h00;
            reg_file[16986] <= 8'h00;
            reg_file[16987] <= 8'h00;
            reg_file[16988] <= 8'h00;
            reg_file[16989] <= 8'h00;
            reg_file[16990] <= 8'h00;
            reg_file[16991] <= 8'h00;
            reg_file[16992] <= 8'h00;
            reg_file[16993] <= 8'h00;
            reg_file[16994] <= 8'h00;
            reg_file[16995] <= 8'h00;
            reg_file[16996] <= 8'h00;
            reg_file[16997] <= 8'h00;
            reg_file[16998] <= 8'h00;
            reg_file[16999] <= 8'h00;
            reg_file[17000] <= 8'h00;
            reg_file[17001] <= 8'h00;
            reg_file[17002] <= 8'h00;
            reg_file[17003] <= 8'h00;
            reg_file[17004] <= 8'h00;
            reg_file[17005] <= 8'h00;
            reg_file[17006] <= 8'h00;
            reg_file[17007] <= 8'h00;
            reg_file[17008] <= 8'h00;
            reg_file[17009] <= 8'h00;
            reg_file[17010] <= 8'h00;
            reg_file[17011] <= 8'h00;
            reg_file[17012] <= 8'h00;
            reg_file[17013] <= 8'h00;
            reg_file[17014] <= 8'h00;
            reg_file[17015] <= 8'h00;
            reg_file[17016] <= 8'h00;
            reg_file[17017] <= 8'h00;
            reg_file[17018] <= 8'h00;
            reg_file[17019] <= 8'h00;
            reg_file[17020] <= 8'h00;
            reg_file[17021] <= 8'h00;
            reg_file[17022] <= 8'h00;
            reg_file[17023] <= 8'h00;
            reg_file[17024] <= 8'h00;
            reg_file[17025] <= 8'h00;
            reg_file[17026] <= 8'h00;
            reg_file[17027] <= 8'h00;
            reg_file[17028] <= 8'h00;
            reg_file[17029] <= 8'h00;
            reg_file[17030] <= 8'h00;
            reg_file[17031] <= 8'h00;
            reg_file[17032] <= 8'h00;
            reg_file[17033] <= 8'h00;
            reg_file[17034] <= 8'h00;
            reg_file[17035] <= 8'h00;
            reg_file[17036] <= 8'h00;
            reg_file[17037] <= 8'h00;
            reg_file[17038] <= 8'h00;
            reg_file[17039] <= 8'h00;
            reg_file[17040] <= 8'h00;
            reg_file[17041] <= 8'h00;
            reg_file[17042] <= 8'h00;
            reg_file[17043] <= 8'h00;
            reg_file[17044] <= 8'h00;
            reg_file[17045] <= 8'h00;
            reg_file[17046] <= 8'h00;
            reg_file[17047] <= 8'h00;
            reg_file[17048] <= 8'h00;
            reg_file[17049] <= 8'h00;
            reg_file[17050] <= 8'h00;
            reg_file[17051] <= 8'h00;
            reg_file[17052] <= 8'h00;
            reg_file[17053] <= 8'h00;
            reg_file[17054] <= 8'h00;
            reg_file[17055] <= 8'h00;
            reg_file[17056] <= 8'h00;
            reg_file[17057] <= 8'h00;
            reg_file[17058] <= 8'h00;
            reg_file[17059] <= 8'h00;
            reg_file[17060] <= 8'h00;
            reg_file[17061] <= 8'h00;
            reg_file[17062] <= 8'h00;
            reg_file[17063] <= 8'h00;
            reg_file[17064] <= 8'h00;
            reg_file[17065] <= 8'h00;
            reg_file[17066] <= 8'h00;
            reg_file[17067] <= 8'h00;
            reg_file[17068] <= 8'h00;
            reg_file[17069] <= 8'h00;
            reg_file[17070] <= 8'h00;
            reg_file[17071] <= 8'h00;
            reg_file[17072] <= 8'h00;
            reg_file[17073] <= 8'h00;
            reg_file[17074] <= 8'h00;
            reg_file[17075] <= 8'h00;
            reg_file[17076] <= 8'h00;
            reg_file[17077] <= 8'h00;
            reg_file[17078] <= 8'h00;
            reg_file[17079] <= 8'h00;
            reg_file[17080] <= 8'h00;
            reg_file[17081] <= 8'h00;
            reg_file[17082] <= 8'h00;
            reg_file[17083] <= 8'h00;
            reg_file[17084] <= 8'h00;
            reg_file[17085] <= 8'h00;
            reg_file[17086] <= 8'h00;
            reg_file[17087] <= 8'h00;
            reg_file[17088] <= 8'h00;
            reg_file[17089] <= 8'h00;
            reg_file[17090] <= 8'h00;
            reg_file[17091] <= 8'h00;
            reg_file[17092] <= 8'h00;
            reg_file[17093] <= 8'h00;
            reg_file[17094] <= 8'h00;
            reg_file[17095] <= 8'h00;
            reg_file[17096] <= 8'h00;
            reg_file[17097] <= 8'h00;
            reg_file[17098] <= 8'h00;
            reg_file[17099] <= 8'h00;
            reg_file[17100] <= 8'h00;
            reg_file[17101] <= 8'h00;
            reg_file[17102] <= 8'h00;
            reg_file[17103] <= 8'h00;
            reg_file[17104] <= 8'h00;
            reg_file[17105] <= 8'h00;
            reg_file[17106] <= 8'h00;
            reg_file[17107] <= 8'h00;
            reg_file[17108] <= 8'h00;
            reg_file[17109] <= 8'h00;
            reg_file[17110] <= 8'h00;
            reg_file[17111] <= 8'h00;
            reg_file[17112] <= 8'h00;
            reg_file[17113] <= 8'h00;
            reg_file[17114] <= 8'h00;
            reg_file[17115] <= 8'h00;
            reg_file[17116] <= 8'h00;
            reg_file[17117] <= 8'h00;
            reg_file[17118] <= 8'h00;
            reg_file[17119] <= 8'h00;
            reg_file[17120] <= 8'h00;
            reg_file[17121] <= 8'h00;
            reg_file[17122] <= 8'h00;
            reg_file[17123] <= 8'h00;
            reg_file[17124] <= 8'h00;
            reg_file[17125] <= 8'h00;
            reg_file[17126] <= 8'h00;
            reg_file[17127] <= 8'h00;
            reg_file[17128] <= 8'h00;
            reg_file[17129] <= 8'h00;
            reg_file[17130] <= 8'h00;
            reg_file[17131] <= 8'h00;
            reg_file[17132] <= 8'h00;
            reg_file[17133] <= 8'h00;
            reg_file[17134] <= 8'h00;
            reg_file[17135] <= 8'h00;
            reg_file[17136] <= 8'h00;
            reg_file[17137] <= 8'h00;
            reg_file[17138] <= 8'h00;
            reg_file[17139] <= 8'h00;
            reg_file[17140] <= 8'h00;
            reg_file[17141] <= 8'h00;
            reg_file[17142] <= 8'h00;
            reg_file[17143] <= 8'h00;
            reg_file[17144] <= 8'h00;
            reg_file[17145] <= 8'h00;
            reg_file[17146] <= 8'h00;
            reg_file[17147] <= 8'h00;
            reg_file[17148] <= 8'h00;
            reg_file[17149] <= 8'h00;
            reg_file[17150] <= 8'h00;
            reg_file[17151] <= 8'h00;
            reg_file[17152] <= 8'h00;
            reg_file[17153] <= 8'h00;
            reg_file[17154] <= 8'h00;
            reg_file[17155] <= 8'h00;
            reg_file[17156] <= 8'h00;
            reg_file[17157] <= 8'h00;
            reg_file[17158] <= 8'h00;
            reg_file[17159] <= 8'h00;
            reg_file[17160] <= 8'h00;
            reg_file[17161] <= 8'h00;
            reg_file[17162] <= 8'h00;
            reg_file[17163] <= 8'h00;
            reg_file[17164] <= 8'h00;
            reg_file[17165] <= 8'h00;
            reg_file[17166] <= 8'h00;
            reg_file[17167] <= 8'h00;
            reg_file[17168] <= 8'h00;
            reg_file[17169] <= 8'h00;
            reg_file[17170] <= 8'h00;
            reg_file[17171] <= 8'h00;
            reg_file[17172] <= 8'h00;
            reg_file[17173] <= 8'h00;
            reg_file[17174] <= 8'h00;
            reg_file[17175] <= 8'h00;
            reg_file[17176] <= 8'h00;
            reg_file[17177] <= 8'h00;
            reg_file[17178] <= 8'h00;
            reg_file[17179] <= 8'h00;
            reg_file[17180] <= 8'h00;
            reg_file[17181] <= 8'h00;
            reg_file[17182] <= 8'h00;
            reg_file[17183] <= 8'h00;
            reg_file[17184] <= 8'h00;
            reg_file[17185] <= 8'h00;
            reg_file[17186] <= 8'h00;
            reg_file[17187] <= 8'h00;
            reg_file[17188] <= 8'h00;
            reg_file[17189] <= 8'h00;
            reg_file[17190] <= 8'h00;
            reg_file[17191] <= 8'h00;
            reg_file[17192] <= 8'h00;
            reg_file[17193] <= 8'h00;
            reg_file[17194] <= 8'h00;
            reg_file[17195] <= 8'h00;
            reg_file[17196] <= 8'h00;
            reg_file[17197] <= 8'h00;
            reg_file[17198] <= 8'h00;
            reg_file[17199] <= 8'h00;
            reg_file[17200] <= 8'h00;
            reg_file[17201] <= 8'h00;
            reg_file[17202] <= 8'h00;
            reg_file[17203] <= 8'h00;
            reg_file[17204] <= 8'h00;
            reg_file[17205] <= 8'h00;
            reg_file[17206] <= 8'h00;
            reg_file[17207] <= 8'h00;
            reg_file[17208] <= 8'h00;
            reg_file[17209] <= 8'h00;
            reg_file[17210] <= 8'h00;
            reg_file[17211] <= 8'h00;
            reg_file[17212] <= 8'h00;
            reg_file[17213] <= 8'h00;
            reg_file[17214] <= 8'h00;
            reg_file[17215] <= 8'h00;
            reg_file[17216] <= 8'h00;
            reg_file[17217] <= 8'h00;
            reg_file[17218] <= 8'h00;
            reg_file[17219] <= 8'h00;
            reg_file[17220] <= 8'h00;
            reg_file[17221] <= 8'h00;
            reg_file[17222] <= 8'h00;
            reg_file[17223] <= 8'h00;
            reg_file[17224] <= 8'h00;
            reg_file[17225] <= 8'h00;
            reg_file[17226] <= 8'h00;
            reg_file[17227] <= 8'h00;
            reg_file[17228] <= 8'h00;
            reg_file[17229] <= 8'h00;
            reg_file[17230] <= 8'h00;
            reg_file[17231] <= 8'h00;
            reg_file[17232] <= 8'h00;
            reg_file[17233] <= 8'h00;
            reg_file[17234] <= 8'h00;
            reg_file[17235] <= 8'h00;
            reg_file[17236] <= 8'h00;
            reg_file[17237] <= 8'h00;
            reg_file[17238] <= 8'h00;
            reg_file[17239] <= 8'h00;
            reg_file[17240] <= 8'h00;
            reg_file[17241] <= 8'h00;
            reg_file[17242] <= 8'h00;
            reg_file[17243] <= 8'h00;
            reg_file[17244] <= 8'h00;
            reg_file[17245] <= 8'h00;
            reg_file[17246] <= 8'h00;
            reg_file[17247] <= 8'h00;
            reg_file[17248] <= 8'h00;
            reg_file[17249] <= 8'h00;
            reg_file[17250] <= 8'h00;
            reg_file[17251] <= 8'h00;
            reg_file[17252] <= 8'h00;
            reg_file[17253] <= 8'h00;
            reg_file[17254] <= 8'h00;
            reg_file[17255] <= 8'h00;
            reg_file[17256] <= 8'h00;
            reg_file[17257] <= 8'h00;
            reg_file[17258] <= 8'h00;
            reg_file[17259] <= 8'h00;
            reg_file[17260] <= 8'h00;
            reg_file[17261] <= 8'h00;
            reg_file[17262] <= 8'h00;
            reg_file[17263] <= 8'h00;
            reg_file[17264] <= 8'h00;
            reg_file[17265] <= 8'h00;
            reg_file[17266] <= 8'h00;
            reg_file[17267] <= 8'h00;
            reg_file[17268] <= 8'h00;
            reg_file[17269] <= 8'h00;
            reg_file[17270] <= 8'h00;
            reg_file[17271] <= 8'h00;
            reg_file[17272] <= 8'h00;
            reg_file[17273] <= 8'h00;
            reg_file[17274] <= 8'h00;
            reg_file[17275] <= 8'h00;
            reg_file[17276] <= 8'h00;
            reg_file[17277] <= 8'h00;
            reg_file[17278] <= 8'h00;
            reg_file[17279] <= 8'h00;
            reg_file[17280] <= 8'h00;
            reg_file[17281] <= 8'h00;
            reg_file[17282] <= 8'h00;
            reg_file[17283] <= 8'h00;
            reg_file[17284] <= 8'h00;
            reg_file[17285] <= 8'h00;
            reg_file[17286] <= 8'h00;
            reg_file[17287] <= 8'h00;
            reg_file[17288] <= 8'h00;
            reg_file[17289] <= 8'h00;
            reg_file[17290] <= 8'h00;
            reg_file[17291] <= 8'h00;
            reg_file[17292] <= 8'h00;
            reg_file[17293] <= 8'h00;
            reg_file[17294] <= 8'h00;
            reg_file[17295] <= 8'h00;
            reg_file[17296] <= 8'h00;
            reg_file[17297] <= 8'h00;
            reg_file[17298] <= 8'h00;
            reg_file[17299] <= 8'h00;
            reg_file[17300] <= 8'h00;
            reg_file[17301] <= 8'h00;
            reg_file[17302] <= 8'h00;
            reg_file[17303] <= 8'h00;
            reg_file[17304] <= 8'h00;
            reg_file[17305] <= 8'h00;
            reg_file[17306] <= 8'h00;
            reg_file[17307] <= 8'h00;
            reg_file[17308] <= 8'h00;
            reg_file[17309] <= 8'h00;
            reg_file[17310] <= 8'h00;
            reg_file[17311] <= 8'h00;
            reg_file[17312] <= 8'h00;
            reg_file[17313] <= 8'h00;
            reg_file[17314] <= 8'h00;
            reg_file[17315] <= 8'h00;
            reg_file[17316] <= 8'h00;
            reg_file[17317] <= 8'h00;
            reg_file[17318] <= 8'h00;
            reg_file[17319] <= 8'h00;
            reg_file[17320] <= 8'h00;
            reg_file[17321] <= 8'h00;
            reg_file[17322] <= 8'h00;
            reg_file[17323] <= 8'h00;
            reg_file[17324] <= 8'h00;
            reg_file[17325] <= 8'h00;
            reg_file[17326] <= 8'h00;
            reg_file[17327] <= 8'h00;
            reg_file[17328] <= 8'h00;
            reg_file[17329] <= 8'h00;
            reg_file[17330] <= 8'h00;
            reg_file[17331] <= 8'h00;
            reg_file[17332] <= 8'h00;
            reg_file[17333] <= 8'h00;
            reg_file[17334] <= 8'h00;
            reg_file[17335] <= 8'h00;
            reg_file[17336] <= 8'h00;
            reg_file[17337] <= 8'h00;
            reg_file[17338] <= 8'h00;
            reg_file[17339] <= 8'h00;
            reg_file[17340] <= 8'h00;
            reg_file[17341] <= 8'h00;
            reg_file[17342] <= 8'h00;
            reg_file[17343] <= 8'h00;
            reg_file[17344] <= 8'h00;
            reg_file[17345] <= 8'h00;
            reg_file[17346] <= 8'h00;
            reg_file[17347] <= 8'h00;
            reg_file[17348] <= 8'h00;
            reg_file[17349] <= 8'h00;
            reg_file[17350] <= 8'h00;
            reg_file[17351] <= 8'h00;
            reg_file[17352] <= 8'h00;
            reg_file[17353] <= 8'h00;
            reg_file[17354] <= 8'h00;
            reg_file[17355] <= 8'h00;
            reg_file[17356] <= 8'h00;
            reg_file[17357] <= 8'h00;
            reg_file[17358] <= 8'h00;
            reg_file[17359] <= 8'h00;
            reg_file[17360] <= 8'h00;
            reg_file[17361] <= 8'h00;
            reg_file[17362] <= 8'h00;
            reg_file[17363] <= 8'h00;
            reg_file[17364] <= 8'h00;
            reg_file[17365] <= 8'h00;
            reg_file[17366] <= 8'h00;
            reg_file[17367] <= 8'h00;
            reg_file[17368] <= 8'h00;
            reg_file[17369] <= 8'h00;
            reg_file[17370] <= 8'h00;
            reg_file[17371] <= 8'h00;
            reg_file[17372] <= 8'h00;
            reg_file[17373] <= 8'h00;
            reg_file[17374] <= 8'h00;
            reg_file[17375] <= 8'h00;
            reg_file[17376] <= 8'h00;
            reg_file[17377] <= 8'h00;
            reg_file[17378] <= 8'h00;
            reg_file[17379] <= 8'h00;
            reg_file[17380] <= 8'h00;
            reg_file[17381] <= 8'h00;
            reg_file[17382] <= 8'h00;
            reg_file[17383] <= 8'h00;
            reg_file[17384] <= 8'h00;
            reg_file[17385] <= 8'h00;
            reg_file[17386] <= 8'h00;
            reg_file[17387] <= 8'h00;
            reg_file[17388] <= 8'h00;
            reg_file[17389] <= 8'h00;
            reg_file[17390] <= 8'h00;
            reg_file[17391] <= 8'h00;
            reg_file[17392] <= 8'h00;
            reg_file[17393] <= 8'h00;
            reg_file[17394] <= 8'h00;
            reg_file[17395] <= 8'h00;
            reg_file[17396] <= 8'h00;
            reg_file[17397] <= 8'h00;
            reg_file[17398] <= 8'h00;
            reg_file[17399] <= 8'h00;
            reg_file[17400] <= 8'h00;
            reg_file[17401] <= 8'h00;
            reg_file[17402] <= 8'h00;
            reg_file[17403] <= 8'h00;
            reg_file[17404] <= 8'h00;
            reg_file[17405] <= 8'h00;
            reg_file[17406] <= 8'h00;
            reg_file[17407] <= 8'h00;
            reg_file[17408] <= 8'h00;
            reg_file[17409] <= 8'h00;
            reg_file[17410] <= 8'h00;
            reg_file[17411] <= 8'h00;
            reg_file[17412] <= 8'h00;
            reg_file[17413] <= 8'h00;
            reg_file[17414] <= 8'h00;
            reg_file[17415] <= 8'h00;
            reg_file[17416] <= 8'h00;
            reg_file[17417] <= 8'h00;
            reg_file[17418] <= 8'h00;
            reg_file[17419] <= 8'h00;
            reg_file[17420] <= 8'h00;
            reg_file[17421] <= 8'h00;
            reg_file[17422] <= 8'h00;
            reg_file[17423] <= 8'h00;
            reg_file[17424] <= 8'h00;
            reg_file[17425] <= 8'h00;
            reg_file[17426] <= 8'h00;
            reg_file[17427] <= 8'h00;
            reg_file[17428] <= 8'h00;
            reg_file[17429] <= 8'h00;
            reg_file[17430] <= 8'h00;
            reg_file[17431] <= 8'h00;
            reg_file[17432] <= 8'h00;
            reg_file[17433] <= 8'h00;
            reg_file[17434] <= 8'h00;
            reg_file[17435] <= 8'h00;
            reg_file[17436] <= 8'h00;
            reg_file[17437] <= 8'h00;
            reg_file[17438] <= 8'h00;
            reg_file[17439] <= 8'h00;
            reg_file[17440] <= 8'h00;
            reg_file[17441] <= 8'h00;
            reg_file[17442] <= 8'h00;
            reg_file[17443] <= 8'h00;
            reg_file[17444] <= 8'h00;
            reg_file[17445] <= 8'h00;
            reg_file[17446] <= 8'h00;
            reg_file[17447] <= 8'h00;
            reg_file[17448] <= 8'h00;
            reg_file[17449] <= 8'h00;
            reg_file[17450] <= 8'h00;
            reg_file[17451] <= 8'h00;
            reg_file[17452] <= 8'h00;
            reg_file[17453] <= 8'h00;
            reg_file[17454] <= 8'h00;
            reg_file[17455] <= 8'h00;
            reg_file[17456] <= 8'h00;
            reg_file[17457] <= 8'h00;
            reg_file[17458] <= 8'h00;
            reg_file[17459] <= 8'h00;
            reg_file[17460] <= 8'h00;
            reg_file[17461] <= 8'h00;
            reg_file[17462] <= 8'h00;
            reg_file[17463] <= 8'h00;
            reg_file[17464] <= 8'h00;
            reg_file[17465] <= 8'h00;
            reg_file[17466] <= 8'h00;
            reg_file[17467] <= 8'h00;
            reg_file[17468] <= 8'h00;
            reg_file[17469] <= 8'h00;
            reg_file[17470] <= 8'h00;
            reg_file[17471] <= 8'h00;
            reg_file[17472] <= 8'h00;
            reg_file[17473] <= 8'h00;
            reg_file[17474] <= 8'h00;
            reg_file[17475] <= 8'h00;
            reg_file[17476] <= 8'h00;
            reg_file[17477] <= 8'h00;
            reg_file[17478] <= 8'h00;
            reg_file[17479] <= 8'h00;
            reg_file[17480] <= 8'h00;
            reg_file[17481] <= 8'h00;
            reg_file[17482] <= 8'h00;
            reg_file[17483] <= 8'h00;
            reg_file[17484] <= 8'h00;
            reg_file[17485] <= 8'h00;
            reg_file[17486] <= 8'h00;
            reg_file[17487] <= 8'h00;
            reg_file[17488] <= 8'h00;
            reg_file[17489] <= 8'h00;
            reg_file[17490] <= 8'h00;
            reg_file[17491] <= 8'h00;
            reg_file[17492] <= 8'h00;
            reg_file[17493] <= 8'h00;
            reg_file[17494] <= 8'h00;
            reg_file[17495] <= 8'h00;
            reg_file[17496] <= 8'h00;
            reg_file[17497] <= 8'h00;
            reg_file[17498] <= 8'h00;
            reg_file[17499] <= 8'h00;
            reg_file[17500] <= 8'h00;
            reg_file[17501] <= 8'h00;
            reg_file[17502] <= 8'h00;
            reg_file[17503] <= 8'h00;
            reg_file[17504] <= 8'h00;
            reg_file[17505] <= 8'h00;
            reg_file[17506] <= 8'h00;
            reg_file[17507] <= 8'h00;
            reg_file[17508] <= 8'h00;
            reg_file[17509] <= 8'h00;
            reg_file[17510] <= 8'h00;
            reg_file[17511] <= 8'h00;
            reg_file[17512] <= 8'h00;
            reg_file[17513] <= 8'h00;
            reg_file[17514] <= 8'h00;
            reg_file[17515] <= 8'h00;
            reg_file[17516] <= 8'h00;
            reg_file[17517] <= 8'h00;
            reg_file[17518] <= 8'h00;
            reg_file[17519] <= 8'h00;
            reg_file[17520] <= 8'h00;
            reg_file[17521] <= 8'h00;
            reg_file[17522] <= 8'h00;
            reg_file[17523] <= 8'h00;
            reg_file[17524] <= 8'h00;
            reg_file[17525] <= 8'h00;
            reg_file[17526] <= 8'h00;
            reg_file[17527] <= 8'h00;
            reg_file[17528] <= 8'h00;
            reg_file[17529] <= 8'h00;
            reg_file[17530] <= 8'h00;
            reg_file[17531] <= 8'h00;
            reg_file[17532] <= 8'h00;
            reg_file[17533] <= 8'h00;
            reg_file[17534] <= 8'h00;
            reg_file[17535] <= 8'h00;
            reg_file[17536] <= 8'h00;
            reg_file[17537] <= 8'h00;
            reg_file[17538] <= 8'h00;
            reg_file[17539] <= 8'h00;
            reg_file[17540] <= 8'h00;
            reg_file[17541] <= 8'h00;
            reg_file[17542] <= 8'h00;
            reg_file[17543] <= 8'h00;
            reg_file[17544] <= 8'h00;
            reg_file[17545] <= 8'h00;
            reg_file[17546] <= 8'h00;
            reg_file[17547] <= 8'h00;
            reg_file[17548] <= 8'h00;
            reg_file[17549] <= 8'h00;
            reg_file[17550] <= 8'h00;
            reg_file[17551] <= 8'h00;
            reg_file[17552] <= 8'h00;
            reg_file[17553] <= 8'h00;
            reg_file[17554] <= 8'h00;
            reg_file[17555] <= 8'h00;
            reg_file[17556] <= 8'h00;
            reg_file[17557] <= 8'h00;
            reg_file[17558] <= 8'h00;
            reg_file[17559] <= 8'h00;
            reg_file[17560] <= 8'h00;
            reg_file[17561] <= 8'h00;
            reg_file[17562] <= 8'h00;
            reg_file[17563] <= 8'h00;
            reg_file[17564] <= 8'h00;
            reg_file[17565] <= 8'h00;
            reg_file[17566] <= 8'h00;
            reg_file[17567] <= 8'h00;
            reg_file[17568] <= 8'h00;
            reg_file[17569] <= 8'h00;
            reg_file[17570] <= 8'h00;
            reg_file[17571] <= 8'h00;
            reg_file[17572] <= 8'h00;
            reg_file[17573] <= 8'h00;
            reg_file[17574] <= 8'h00;
            reg_file[17575] <= 8'h00;
            reg_file[17576] <= 8'h00;
            reg_file[17577] <= 8'h00;
            reg_file[17578] <= 8'h00;
            reg_file[17579] <= 8'h00;
            reg_file[17580] <= 8'h00;
            reg_file[17581] <= 8'h00;
            reg_file[17582] <= 8'h00;
            reg_file[17583] <= 8'h00;
            reg_file[17584] <= 8'h00;
            reg_file[17585] <= 8'h00;
            reg_file[17586] <= 8'h00;
            reg_file[17587] <= 8'h00;
            reg_file[17588] <= 8'h00;
            reg_file[17589] <= 8'h00;
            reg_file[17590] <= 8'h00;
            reg_file[17591] <= 8'h00;
            reg_file[17592] <= 8'h00;
            reg_file[17593] <= 8'h00;
            reg_file[17594] <= 8'h00;
            reg_file[17595] <= 8'h00;
            reg_file[17596] <= 8'h00;
            reg_file[17597] <= 8'h00;
            reg_file[17598] <= 8'h00;
            reg_file[17599] <= 8'h00;
            reg_file[17600] <= 8'h00;
            reg_file[17601] <= 8'h00;
            reg_file[17602] <= 8'h00;
            reg_file[17603] <= 8'h00;
            reg_file[17604] <= 8'h00;
            reg_file[17605] <= 8'h00;
            reg_file[17606] <= 8'h00;
            reg_file[17607] <= 8'h00;
            reg_file[17608] <= 8'h00;
            reg_file[17609] <= 8'h00;
            reg_file[17610] <= 8'h00;
            reg_file[17611] <= 8'h00;
            reg_file[17612] <= 8'h00;
            reg_file[17613] <= 8'h00;
            reg_file[17614] <= 8'h00;
            reg_file[17615] <= 8'h00;
            reg_file[17616] <= 8'h00;
            reg_file[17617] <= 8'h00;
            reg_file[17618] <= 8'h00;
            reg_file[17619] <= 8'h00;
            reg_file[17620] <= 8'h00;
            reg_file[17621] <= 8'h00;
            reg_file[17622] <= 8'h00;
            reg_file[17623] <= 8'h00;
            reg_file[17624] <= 8'h00;
            reg_file[17625] <= 8'h00;
            reg_file[17626] <= 8'h00;
            reg_file[17627] <= 8'h00;
            reg_file[17628] <= 8'h00;
            reg_file[17629] <= 8'h00;
            reg_file[17630] <= 8'h00;
            reg_file[17631] <= 8'h00;
            reg_file[17632] <= 8'h00;
            reg_file[17633] <= 8'h00;
            reg_file[17634] <= 8'h00;
            reg_file[17635] <= 8'h00;
            reg_file[17636] <= 8'h00;
            reg_file[17637] <= 8'h00;
            reg_file[17638] <= 8'h00;
            reg_file[17639] <= 8'h00;
            reg_file[17640] <= 8'h00;
            reg_file[17641] <= 8'h00;
            reg_file[17642] <= 8'h00;
            reg_file[17643] <= 8'h00;
            reg_file[17644] <= 8'h00;
            reg_file[17645] <= 8'h00;
            reg_file[17646] <= 8'h00;
            reg_file[17647] <= 8'h00;
            reg_file[17648] <= 8'h00;
            reg_file[17649] <= 8'h00;
            reg_file[17650] <= 8'h00;
            reg_file[17651] <= 8'h00;
            reg_file[17652] <= 8'h00;
            reg_file[17653] <= 8'h00;
            reg_file[17654] <= 8'h00;
            reg_file[17655] <= 8'h00;
            reg_file[17656] <= 8'h00;
            reg_file[17657] <= 8'h00;
            reg_file[17658] <= 8'h00;
            reg_file[17659] <= 8'h00;
            reg_file[17660] <= 8'h00;
            reg_file[17661] <= 8'h00;
            reg_file[17662] <= 8'h00;
            reg_file[17663] <= 8'h00;
            reg_file[17664] <= 8'h00;
            reg_file[17665] <= 8'h00;
            reg_file[17666] <= 8'h00;
            reg_file[17667] <= 8'h00;
            reg_file[17668] <= 8'h00;
            reg_file[17669] <= 8'h00;
            reg_file[17670] <= 8'h00;
            reg_file[17671] <= 8'h00;
            reg_file[17672] <= 8'h00;
            reg_file[17673] <= 8'h00;
            reg_file[17674] <= 8'h00;
            reg_file[17675] <= 8'h00;
            reg_file[17676] <= 8'h00;
            reg_file[17677] <= 8'h00;
            reg_file[17678] <= 8'h00;
            reg_file[17679] <= 8'h00;
            reg_file[17680] <= 8'h00;
            reg_file[17681] <= 8'h00;
            reg_file[17682] <= 8'h00;
            reg_file[17683] <= 8'h00;
            reg_file[17684] <= 8'h00;
            reg_file[17685] <= 8'h00;
            reg_file[17686] <= 8'h00;
            reg_file[17687] <= 8'h00;
            reg_file[17688] <= 8'h00;
            reg_file[17689] <= 8'h00;
            reg_file[17690] <= 8'h00;
            reg_file[17691] <= 8'h00;
            reg_file[17692] <= 8'h00;
            reg_file[17693] <= 8'h00;
            reg_file[17694] <= 8'h00;
            reg_file[17695] <= 8'h00;
            reg_file[17696] <= 8'h00;
            reg_file[17697] <= 8'h00;
            reg_file[17698] <= 8'h00;
            reg_file[17699] <= 8'h00;
            reg_file[17700] <= 8'h00;
            reg_file[17701] <= 8'h00;
            reg_file[17702] <= 8'h00;
            reg_file[17703] <= 8'h00;
            reg_file[17704] <= 8'h00;
            reg_file[17705] <= 8'h00;
            reg_file[17706] <= 8'h00;
            reg_file[17707] <= 8'h00;
            reg_file[17708] <= 8'h00;
            reg_file[17709] <= 8'h00;
            reg_file[17710] <= 8'h00;
            reg_file[17711] <= 8'h00;
            reg_file[17712] <= 8'h00;
            reg_file[17713] <= 8'h00;
            reg_file[17714] <= 8'h00;
            reg_file[17715] <= 8'h00;
            reg_file[17716] <= 8'h00;
            reg_file[17717] <= 8'h00;
            reg_file[17718] <= 8'h00;
            reg_file[17719] <= 8'h00;
            reg_file[17720] <= 8'h00;
            reg_file[17721] <= 8'h00;
            reg_file[17722] <= 8'h00;
            reg_file[17723] <= 8'h00;
            reg_file[17724] <= 8'h00;
            reg_file[17725] <= 8'h00;
            reg_file[17726] <= 8'h00;
            reg_file[17727] <= 8'h00;
            reg_file[17728] <= 8'h00;
            reg_file[17729] <= 8'h00;
            reg_file[17730] <= 8'h00;
            reg_file[17731] <= 8'h00;
            reg_file[17732] <= 8'h00;
            reg_file[17733] <= 8'h00;
            reg_file[17734] <= 8'h00;
            reg_file[17735] <= 8'h00;
            reg_file[17736] <= 8'h00;
            reg_file[17737] <= 8'h00;
            reg_file[17738] <= 8'h00;
            reg_file[17739] <= 8'h00;
            reg_file[17740] <= 8'h00;
            reg_file[17741] <= 8'h00;
            reg_file[17742] <= 8'h00;
            reg_file[17743] <= 8'h00;
            reg_file[17744] <= 8'h00;
            reg_file[17745] <= 8'h00;
            reg_file[17746] <= 8'h00;
            reg_file[17747] <= 8'h00;
            reg_file[17748] <= 8'h00;
            reg_file[17749] <= 8'h00;
            reg_file[17750] <= 8'h00;
            reg_file[17751] <= 8'h00;
            reg_file[17752] <= 8'h00;
            reg_file[17753] <= 8'h00;
            reg_file[17754] <= 8'h00;
            reg_file[17755] <= 8'h00;
            reg_file[17756] <= 8'h00;
            reg_file[17757] <= 8'h00;
            reg_file[17758] <= 8'h00;
            reg_file[17759] <= 8'h00;
            reg_file[17760] <= 8'h00;
            reg_file[17761] <= 8'h00;
            reg_file[17762] <= 8'h00;
            reg_file[17763] <= 8'h00;
            reg_file[17764] <= 8'h00;
            reg_file[17765] <= 8'h00;
            reg_file[17766] <= 8'h00;
            reg_file[17767] <= 8'h00;
            reg_file[17768] <= 8'h00;
            reg_file[17769] <= 8'h00;
            reg_file[17770] <= 8'h00;
            reg_file[17771] <= 8'h00;
            reg_file[17772] <= 8'h00;
            reg_file[17773] <= 8'h00;
            reg_file[17774] <= 8'h00;
            reg_file[17775] <= 8'h00;
            reg_file[17776] <= 8'h00;
            reg_file[17777] <= 8'h00;
            reg_file[17778] <= 8'h00;
            reg_file[17779] <= 8'h00;
            reg_file[17780] <= 8'h00;
            reg_file[17781] <= 8'h00;
            reg_file[17782] <= 8'h00;
            reg_file[17783] <= 8'h00;
            reg_file[17784] <= 8'h00;
            reg_file[17785] <= 8'h00;
            reg_file[17786] <= 8'h00;
            reg_file[17787] <= 8'h00;
            reg_file[17788] <= 8'h00;
            reg_file[17789] <= 8'h00;
            reg_file[17790] <= 8'h00;
            reg_file[17791] <= 8'h00;
            reg_file[17792] <= 8'h00;
            reg_file[17793] <= 8'h00;
            reg_file[17794] <= 8'h00;
            reg_file[17795] <= 8'h00;
            reg_file[17796] <= 8'h00;
            reg_file[17797] <= 8'h00;
            reg_file[17798] <= 8'h00;
            reg_file[17799] <= 8'h00;
            reg_file[17800] <= 8'h00;
            reg_file[17801] <= 8'h00;
            reg_file[17802] <= 8'h00;
            reg_file[17803] <= 8'h00;
            reg_file[17804] <= 8'h00;
            reg_file[17805] <= 8'h00;
            reg_file[17806] <= 8'h00;
            reg_file[17807] <= 8'h00;
            reg_file[17808] <= 8'h00;
            reg_file[17809] <= 8'h00;
            reg_file[17810] <= 8'h00;
            reg_file[17811] <= 8'h00;
            reg_file[17812] <= 8'h00;
            reg_file[17813] <= 8'h00;
            reg_file[17814] <= 8'h00;
            reg_file[17815] <= 8'h00;
            reg_file[17816] <= 8'h00;
            reg_file[17817] <= 8'h00;
            reg_file[17818] <= 8'h00;
            reg_file[17819] <= 8'h00;
            reg_file[17820] <= 8'h00;
            reg_file[17821] <= 8'h00;
            reg_file[17822] <= 8'h00;
            reg_file[17823] <= 8'h00;
            reg_file[17824] <= 8'h00;
            reg_file[17825] <= 8'h00;
            reg_file[17826] <= 8'h00;
            reg_file[17827] <= 8'h00;
            reg_file[17828] <= 8'h00;
            reg_file[17829] <= 8'h00;
            reg_file[17830] <= 8'h00;
            reg_file[17831] <= 8'h00;
            reg_file[17832] <= 8'h00;
            reg_file[17833] <= 8'h00;
            reg_file[17834] <= 8'h00;
            reg_file[17835] <= 8'h00;
            reg_file[17836] <= 8'h00;
            reg_file[17837] <= 8'h00;
            reg_file[17838] <= 8'h00;
            reg_file[17839] <= 8'h00;
            reg_file[17840] <= 8'h00;
            reg_file[17841] <= 8'h00;
            reg_file[17842] <= 8'h00;
            reg_file[17843] <= 8'h00;
            reg_file[17844] <= 8'h00;
            reg_file[17845] <= 8'h00;
            reg_file[17846] <= 8'h00;
            reg_file[17847] <= 8'h00;
            reg_file[17848] <= 8'h00;
            reg_file[17849] <= 8'h00;
            reg_file[17850] <= 8'h00;
            reg_file[17851] <= 8'h00;
            reg_file[17852] <= 8'h00;
            reg_file[17853] <= 8'h00;
            reg_file[17854] <= 8'h00;
            reg_file[17855] <= 8'h00;
            reg_file[17856] <= 8'h00;
            reg_file[17857] <= 8'h00;
            reg_file[17858] <= 8'h00;
            reg_file[17859] <= 8'h00;
            reg_file[17860] <= 8'h00;
            reg_file[17861] <= 8'h00;
            reg_file[17862] <= 8'h00;
            reg_file[17863] <= 8'h00;
            reg_file[17864] <= 8'h00;
            reg_file[17865] <= 8'h00;
            reg_file[17866] <= 8'h00;
            reg_file[17867] <= 8'h00;
            reg_file[17868] <= 8'h00;
            reg_file[17869] <= 8'h00;
            reg_file[17870] <= 8'h00;
            reg_file[17871] <= 8'h00;
            reg_file[17872] <= 8'h00;
            reg_file[17873] <= 8'h00;
            reg_file[17874] <= 8'h00;
            reg_file[17875] <= 8'h00;
            reg_file[17876] <= 8'h00;
            reg_file[17877] <= 8'h00;
            reg_file[17878] <= 8'h00;
            reg_file[17879] <= 8'h00;
            reg_file[17880] <= 8'h00;
            reg_file[17881] <= 8'h00;
            reg_file[17882] <= 8'h00;
            reg_file[17883] <= 8'h00;
            reg_file[17884] <= 8'h00;
            reg_file[17885] <= 8'h00;
            reg_file[17886] <= 8'h00;
            reg_file[17887] <= 8'h00;
            reg_file[17888] <= 8'h00;
            reg_file[17889] <= 8'h00;
            reg_file[17890] <= 8'h00;
            reg_file[17891] <= 8'h00;
            reg_file[17892] <= 8'h00;
            reg_file[17893] <= 8'h00;
            reg_file[17894] <= 8'h00;
            reg_file[17895] <= 8'h00;
            reg_file[17896] <= 8'h00;
            reg_file[17897] <= 8'h00;
            reg_file[17898] <= 8'h00;
            reg_file[17899] <= 8'h00;
            reg_file[17900] <= 8'h00;
            reg_file[17901] <= 8'h00;
            reg_file[17902] <= 8'h00;
            reg_file[17903] <= 8'h00;
            reg_file[17904] <= 8'h00;
            reg_file[17905] <= 8'h00;
            reg_file[17906] <= 8'h00;
            reg_file[17907] <= 8'h00;
            reg_file[17908] <= 8'h00;
            reg_file[17909] <= 8'h00;
            reg_file[17910] <= 8'h00;
            reg_file[17911] <= 8'h00;
            reg_file[17912] <= 8'h00;
            reg_file[17913] <= 8'h00;
            reg_file[17914] <= 8'h00;
            reg_file[17915] <= 8'h00;
            reg_file[17916] <= 8'h00;
            reg_file[17917] <= 8'h00;
            reg_file[17918] <= 8'h00;
            reg_file[17919] <= 8'h00;
            reg_file[17920] <= 8'h00;
            reg_file[17921] <= 8'h00;
            reg_file[17922] <= 8'h00;
            reg_file[17923] <= 8'h00;
            reg_file[17924] <= 8'h00;
            reg_file[17925] <= 8'h00;
            reg_file[17926] <= 8'h00;
            reg_file[17927] <= 8'h00;
            reg_file[17928] <= 8'h00;
            reg_file[17929] <= 8'h00;
            reg_file[17930] <= 8'h00;
            reg_file[17931] <= 8'h00;
            reg_file[17932] <= 8'h00;
            reg_file[17933] <= 8'h00;
            reg_file[17934] <= 8'h00;
            reg_file[17935] <= 8'h00;
            reg_file[17936] <= 8'h00;
            reg_file[17937] <= 8'h00;
            reg_file[17938] <= 8'h00;
            reg_file[17939] <= 8'h00;
            reg_file[17940] <= 8'h00;
            reg_file[17941] <= 8'h00;
            reg_file[17942] <= 8'h00;
            reg_file[17943] <= 8'h00;
            reg_file[17944] <= 8'h00;
            reg_file[17945] <= 8'h00;
            reg_file[17946] <= 8'h00;
            reg_file[17947] <= 8'h00;
            reg_file[17948] <= 8'h00;
            reg_file[17949] <= 8'h00;
            reg_file[17950] <= 8'h00;
            reg_file[17951] <= 8'h00;
            reg_file[17952] <= 8'h00;
            reg_file[17953] <= 8'h00;
            reg_file[17954] <= 8'h00;
            reg_file[17955] <= 8'h00;
            reg_file[17956] <= 8'h00;
            reg_file[17957] <= 8'h00;
            reg_file[17958] <= 8'h00;
            reg_file[17959] <= 8'h00;
            reg_file[17960] <= 8'h00;
            reg_file[17961] <= 8'h00;
            reg_file[17962] <= 8'h00;
            reg_file[17963] <= 8'h00;
            reg_file[17964] <= 8'h00;
            reg_file[17965] <= 8'h00;
            reg_file[17966] <= 8'h00;
            reg_file[17967] <= 8'h00;
            reg_file[17968] <= 8'h00;
            reg_file[17969] <= 8'h00;
            reg_file[17970] <= 8'h00;
            reg_file[17971] <= 8'h00;
            reg_file[17972] <= 8'h00;
            reg_file[17973] <= 8'h00;
            reg_file[17974] <= 8'h00;
            reg_file[17975] <= 8'h00;
            reg_file[17976] <= 8'h00;
            reg_file[17977] <= 8'h00;
            reg_file[17978] <= 8'h00;
            reg_file[17979] <= 8'h00;
            reg_file[17980] <= 8'h00;
            reg_file[17981] <= 8'h00;
            reg_file[17982] <= 8'h00;
            reg_file[17983] <= 8'h00;
            reg_file[17984] <= 8'h00;
            reg_file[17985] <= 8'h00;
            reg_file[17986] <= 8'h00;
            reg_file[17987] <= 8'h00;
            reg_file[17988] <= 8'h00;
            reg_file[17989] <= 8'h00;
            reg_file[17990] <= 8'h00;
            reg_file[17991] <= 8'h00;
            reg_file[17992] <= 8'h00;
            reg_file[17993] <= 8'h00;
            reg_file[17994] <= 8'h00;
            reg_file[17995] <= 8'h00;
            reg_file[17996] <= 8'h00;
            reg_file[17997] <= 8'h00;
            reg_file[17998] <= 8'h00;
            reg_file[17999] <= 8'h00;
            reg_file[18000] <= 8'h00;
            reg_file[18001] <= 8'h00;
            reg_file[18002] <= 8'h00;
            reg_file[18003] <= 8'h00;
            reg_file[18004] <= 8'h00;
            reg_file[18005] <= 8'h00;
            reg_file[18006] <= 8'h00;
            reg_file[18007] <= 8'h00;
            reg_file[18008] <= 8'h00;
            reg_file[18009] <= 8'h00;
            reg_file[18010] <= 8'h00;
            reg_file[18011] <= 8'h00;
            reg_file[18012] <= 8'h00;
            reg_file[18013] <= 8'h00;
            reg_file[18014] <= 8'h00;
            reg_file[18015] <= 8'h00;
            reg_file[18016] <= 8'h00;
            reg_file[18017] <= 8'h00;
            reg_file[18018] <= 8'h00;
            reg_file[18019] <= 8'h00;
            reg_file[18020] <= 8'h00;
            reg_file[18021] <= 8'h00;
            reg_file[18022] <= 8'h00;
            reg_file[18023] <= 8'h00;
            reg_file[18024] <= 8'h00;
            reg_file[18025] <= 8'h00;
            reg_file[18026] <= 8'h00;
            reg_file[18027] <= 8'h00;
            reg_file[18028] <= 8'h00;
            reg_file[18029] <= 8'h00;
            reg_file[18030] <= 8'h00;
            reg_file[18031] <= 8'h00;
            reg_file[18032] <= 8'h00;
            reg_file[18033] <= 8'h00;
            reg_file[18034] <= 8'h00;
            reg_file[18035] <= 8'h00;
            reg_file[18036] <= 8'h00;
            reg_file[18037] <= 8'h00;
            reg_file[18038] <= 8'h00;
            reg_file[18039] <= 8'h00;
            reg_file[18040] <= 8'h00;
            reg_file[18041] <= 8'h00;
            reg_file[18042] <= 8'h00;
            reg_file[18043] <= 8'h00;
            reg_file[18044] <= 8'h00;
            reg_file[18045] <= 8'h00;
            reg_file[18046] <= 8'h00;
            reg_file[18047] <= 8'h00;
            reg_file[18048] <= 8'h00;
            reg_file[18049] <= 8'h00;
            reg_file[18050] <= 8'h00;
            reg_file[18051] <= 8'h00;
            reg_file[18052] <= 8'h00;
            reg_file[18053] <= 8'h00;
            reg_file[18054] <= 8'h00;
            reg_file[18055] <= 8'h00;
            reg_file[18056] <= 8'h00;
            reg_file[18057] <= 8'h00;
            reg_file[18058] <= 8'h00;
            reg_file[18059] <= 8'h00;
            reg_file[18060] <= 8'h00;
            reg_file[18061] <= 8'h00;
            reg_file[18062] <= 8'h00;
            reg_file[18063] <= 8'h00;
            reg_file[18064] <= 8'h00;
            reg_file[18065] <= 8'h00;
            reg_file[18066] <= 8'h00;
            reg_file[18067] <= 8'h00;
            reg_file[18068] <= 8'h00;
            reg_file[18069] <= 8'h00;
            reg_file[18070] <= 8'h00;
            reg_file[18071] <= 8'h00;
            reg_file[18072] <= 8'h00;
            reg_file[18073] <= 8'h00;
            reg_file[18074] <= 8'h00;
            reg_file[18075] <= 8'h00;
            reg_file[18076] <= 8'h00;
            reg_file[18077] <= 8'h00;
            reg_file[18078] <= 8'h00;
            reg_file[18079] <= 8'h00;
            reg_file[18080] <= 8'h00;
            reg_file[18081] <= 8'h00;
            reg_file[18082] <= 8'h00;
            reg_file[18083] <= 8'h00;
            reg_file[18084] <= 8'h00;
            reg_file[18085] <= 8'h00;
            reg_file[18086] <= 8'h00;
            reg_file[18087] <= 8'h00;
            reg_file[18088] <= 8'h00;
            reg_file[18089] <= 8'h00;
            reg_file[18090] <= 8'h00;
            reg_file[18091] <= 8'h00;
            reg_file[18092] <= 8'h00;
            reg_file[18093] <= 8'h00;
            reg_file[18094] <= 8'h00;
            reg_file[18095] <= 8'h00;
            reg_file[18096] <= 8'h00;
            reg_file[18097] <= 8'h00;
            reg_file[18098] <= 8'h00;
            reg_file[18099] <= 8'h00;
            reg_file[18100] <= 8'h00;
            reg_file[18101] <= 8'h00;
            reg_file[18102] <= 8'h00;
            reg_file[18103] <= 8'h00;
            reg_file[18104] <= 8'h00;
            reg_file[18105] <= 8'h00;
            reg_file[18106] <= 8'h00;
            reg_file[18107] <= 8'h00;
            reg_file[18108] <= 8'h00;
            reg_file[18109] <= 8'h00;
            reg_file[18110] <= 8'h00;
            reg_file[18111] <= 8'h00;
            reg_file[18112] <= 8'h00;
            reg_file[18113] <= 8'h00;
            reg_file[18114] <= 8'h00;
            reg_file[18115] <= 8'h00;
            reg_file[18116] <= 8'h00;
            reg_file[18117] <= 8'h00;
            reg_file[18118] <= 8'h00;
            reg_file[18119] <= 8'h00;
            reg_file[18120] <= 8'h00;
            reg_file[18121] <= 8'h00;
            reg_file[18122] <= 8'h00;
            reg_file[18123] <= 8'h00;
            reg_file[18124] <= 8'h00;
            reg_file[18125] <= 8'h00;
            reg_file[18126] <= 8'h00;
            reg_file[18127] <= 8'h00;
            reg_file[18128] <= 8'h00;
            reg_file[18129] <= 8'h00;
            reg_file[18130] <= 8'h00;
            reg_file[18131] <= 8'h00;
            reg_file[18132] <= 8'h00;
            reg_file[18133] <= 8'h00;
            reg_file[18134] <= 8'h00;
            reg_file[18135] <= 8'h00;
            reg_file[18136] <= 8'h00;
            reg_file[18137] <= 8'h00;
            reg_file[18138] <= 8'h00;
            reg_file[18139] <= 8'h00;
            reg_file[18140] <= 8'h00;
            reg_file[18141] <= 8'h00;
            reg_file[18142] <= 8'h00;
            reg_file[18143] <= 8'h00;
            reg_file[18144] <= 8'h00;
            reg_file[18145] <= 8'h00;
            reg_file[18146] <= 8'h00;
            reg_file[18147] <= 8'h00;
            reg_file[18148] <= 8'h00;
            reg_file[18149] <= 8'h00;
            reg_file[18150] <= 8'h00;
            reg_file[18151] <= 8'h00;
            reg_file[18152] <= 8'h00;
            reg_file[18153] <= 8'h00;
            reg_file[18154] <= 8'h00;
            reg_file[18155] <= 8'h00;
            reg_file[18156] <= 8'h00;
            reg_file[18157] <= 8'h00;
            reg_file[18158] <= 8'h00;
            reg_file[18159] <= 8'h00;
            reg_file[18160] <= 8'h00;
            reg_file[18161] <= 8'h00;
            reg_file[18162] <= 8'h00;
            reg_file[18163] <= 8'h00;
            reg_file[18164] <= 8'h00;
            reg_file[18165] <= 8'h00;
            reg_file[18166] <= 8'h00;
            reg_file[18167] <= 8'h00;
            reg_file[18168] <= 8'h00;
            reg_file[18169] <= 8'h00;
            reg_file[18170] <= 8'h00;
            reg_file[18171] <= 8'h00;
            reg_file[18172] <= 8'h00;
            reg_file[18173] <= 8'h00;
            reg_file[18174] <= 8'h00;
            reg_file[18175] <= 8'h00;
            reg_file[18176] <= 8'h00;
            reg_file[18177] <= 8'h00;
            reg_file[18178] <= 8'h00;
            reg_file[18179] <= 8'h00;
            reg_file[18180] <= 8'h00;
            reg_file[18181] <= 8'h00;
            reg_file[18182] <= 8'h00;
            reg_file[18183] <= 8'h00;
            reg_file[18184] <= 8'h00;
            reg_file[18185] <= 8'h00;
            reg_file[18186] <= 8'h00;
            reg_file[18187] <= 8'h00;
            reg_file[18188] <= 8'h00;
            reg_file[18189] <= 8'h00;
            reg_file[18190] <= 8'h00;
            reg_file[18191] <= 8'h00;
            reg_file[18192] <= 8'h00;
            reg_file[18193] <= 8'h00;
            reg_file[18194] <= 8'h00;
            reg_file[18195] <= 8'h00;
            reg_file[18196] <= 8'h00;
            reg_file[18197] <= 8'h00;
            reg_file[18198] <= 8'h00;
            reg_file[18199] <= 8'h00;
            reg_file[18200] <= 8'h00;
            reg_file[18201] <= 8'h00;
            reg_file[18202] <= 8'h00;
            reg_file[18203] <= 8'h00;
            reg_file[18204] <= 8'h00;
            reg_file[18205] <= 8'h00;
            reg_file[18206] <= 8'h00;
            reg_file[18207] <= 8'h00;
            reg_file[18208] <= 8'h00;
            reg_file[18209] <= 8'h00;
            reg_file[18210] <= 8'h00;
            reg_file[18211] <= 8'h00;
            reg_file[18212] <= 8'h00;
            reg_file[18213] <= 8'h00;
            reg_file[18214] <= 8'h00;
            reg_file[18215] <= 8'h00;
            reg_file[18216] <= 8'h00;
            reg_file[18217] <= 8'h00;
            reg_file[18218] <= 8'h00;
            reg_file[18219] <= 8'h00;
            reg_file[18220] <= 8'h00;
            reg_file[18221] <= 8'h00;
            reg_file[18222] <= 8'h00;
            reg_file[18223] <= 8'h00;
            reg_file[18224] <= 8'h00;
            reg_file[18225] <= 8'h00;
            reg_file[18226] <= 8'h00;
            reg_file[18227] <= 8'h00;
            reg_file[18228] <= 8'h00;
            reg_file[18229] <= 8'h00;
            reg_file[18230] <= 8'h00;
            reg_file[18231] <= 8'h00;
            reg_file[18232] <= 8'h00;
            reg_file[18233] <= 8'h00;
            reg_file[18234] <= 8'h00;
            reg_file[18235] <= 8'h00;
            reg_file[18236] <= 8'h00;
            reg_file[18237] <= 8'h00;
            reg_file[18238] <= 8'h00;
            reg_file[18239] <= 8'h00;
            reg_file[18240] <= 8'h00;
            reg_file[18241] <= 8'h00;
            reg_file[18242] <= 8'h00;
            reg_file[18243] <= 8'h00;
            reg_file[18244] <= 8'h00;
            reg_file[18245] <= 8'h00;
            reg_file[18246] <= 8'h00;
            reg_file[18247] <= 8'h00;
            reg_file[18248] <= 8'h00;
            reg_file[18249] <= 8'h00;
            reg_file[18250] <= 8'h00;
            reg_file[18251] <= 8'h00;
            reg_file[18252] <= 8'h00;
            reg_file[18253] <= 8'h00;
            reg_file[18254] <= 8'h00;
            reg_file[18255] <= 8'h00;
            reg_file[18256] <= 8'h00;
            reg_file[18257] <= 8'h00;
            reg_file[18258] <= 8'h00;
            reg_file[18259] <= 8'h00;
            reg_file[18260] <= 8'h00;
            reg_file[18261] <= 8'h00;
            reg_file[18262] <= 8'h00;
            reg_file[18263] <= 8'h00;
            reg_file[18264] <= 8'h00;
            reg_file[18265] <= 8'h00;
            reg_file[18266] <= 8'h00;
            reg_file[18267] <= 8'h00;
            reg_file[18268] <= 8'h00;
            reg_file[18269] <= 8'h00;
            reg_file[18270] <= 8'h00;
            reg_file[18271] <= 8'h00;
            reg_file[18272] <= 8'h00;
            reg_file[18273] <= 8'h00;
            reg_file[18274] <= 8'h00;
            reg_file[18275] <= 8'h00;
            reg_file[18276] <= 8'h00;
            reg_file[18277] <= 8'h00;
            reg_file[18278] <= 8'h00;
            reg_file[18279] <= 8'h00;
            reg_file[18280] <= 8'h00;
            reg_file[18281] <= 8'h00;
            reg_file[18282] <= 8'h00;
            reg_file[18283] <= 8'h00;
            reg_file[18284] <= 8'h00;
            reg_file[18285] <= 8'h00;
            reg_file[18286] <= 8'h00;
            reg_file[18287] <= 8'h00;
            reg_file[18288] <= 8'h00;
            reg_file[18289] <= 8'h00;
            reg_file[18290] <= 8'h00;
            reg_file[18291] <= 8'h00;
            reg_file[18292] <= 8'h00;
            reg_file[18293] <= 8'h00;
            reg_file[18294] <= 8'h00;
            reg_file[18295] <= 8'h00;
            reg_file[18296] <= 8'h00;
            reg_file[18297] <= 8'h00;
            reg_file[18298] <= 8'h00;
            reg_file[18299] <= 8'h00;
            reg_file[18300] <= 8'h00;
            reg_file[18301] <= 8'h00;
            reg_file[18302] <= 8'h00;
            reg_file[18303] <= 8'h00;
            reg_file[18304] <= 8'h00;
            reg_file[18305] <= 8'h00;
            reg_file[18306] <= 8'h00;
            reg_file[18307] <= 8'h00;
            reg_file[18308] <= 8'h00;
            reg_file[18309] <= 8'h00;
            reg_file[18310] <= 8'h00;
            reg_file[18311] <= 8'h00;
            reg_file[18312] <= 8'h00;
            reg_file[18313] <= 8'h00;
            reg_file[18314] <= 8'h00;
            reg_file[18315] <= 8'h00;
            reg_file[18316] <= 8'h00;
            reg_file[18317] <= 8'h00;
            reg_file[18318] <= 8'h00;
            reg_file[18319] <= 8'h00;
            reg_file[18320] <= 8'h00;
            reg_file[18321] <= 8'h00;
            reg_file[18322] <= 8'h00;
            reg_file[18323] <= 8'h00;
            reg_file[18324] <= 8'h00;
            reg_file[18325] <= 8'h00;
            reg_file[18326] <= 8'h00;
            reg_file[18327] <= 8'h00;
            reg_file[18328] <= 8'h00;
            reg_file[18329] <= 8'h00;
            reg_file[18330] <= 8'h00;
            reg_file[18331] <= 8'h00;
            reg_file[18332] <= 8'h00;
            reg_file[18333] <= 8'h00;
            reg_file[18334] <= 8'h00;
            reg_file[18335] <= 8'h00;
            reg_file[18336] <= 8'h00;
            reg_file[18337] <= 8'h00;
            reg_file[18338] <= 8'h00;
            reg_file[18339] <= 8'h00;
            reg_file[18340] <= 8'h00;
            reg_file[18341] <= 8'h00;
            reg_file[18342] <= 8'h00;
            reg_file[18343] <= 8'h00;
            reg_file[18344] <= 8'h00;
            reg_file[18345] <= 8'h00;
            reg_file[18346] <= 8'h00;
            reg_file[18347] <= 8'h00;
            reg_file[18348] <= 8'h00;
            reg_file[18349] <= 8'h00;
            reg_file[18350] <= 8'h00;
            reg_file[18351] <= 8'h00;
            reg_file[18352] <= 8'h00;
            reg_file[18353] <= 8'h00;
            reg_file[18354] <= 8'h00;
            reg_file[18355] <= 8'h00;
            reg_file[18356] <= 8'h00;
            reg_file[18357] <= 8'h00;
            reg_file[18358] <= 8'h00;
            reg_file[18359] <= 8'h00;
            reg_file[18360] <= 8'h00;
            reg_file[18361] <= 8'h00;
            reg_file[18362] <= 8'h00;
            reg_file[18363] <= 8'h00;
            reg_file[18364] <= 8'h00;
            reg_file[18365] <= 8'h00;
            reg_file[18366] <= 8'h00;
            reg_file[18367] <= 8'h00;
            reg_file[18368] <= 8'h00;
            reg_file[18369] <= 8'h00;
            reg_file[18370] <= 8'h00;
            reg_file[18371] <= 8'h00;
            reg_file[18372] <= 8'h00;
            reg_file[18373] <= 8'h00;
            reg_file[18374] <= 8'h00;
            reg_file[18375] <= 8'h00;
            reg_file[18376] <= 8'h00;
            reg_file[18377] <= 8'h00;
            reg_file[18378] <= 8'h00;
            reg_file[18379] <= 8'h00;
            reg_file[18380] <= 8'h00;
            reg_file[18381] <= 8'h00;
            reg_file[18382] <= 8'h00;
            reg_file[18383] <= 8'h00;
            reg_file[18384] <= 8'h00;
            reg_file[18385] <= 8'h00;
            reg_file[18386] <= 8'h00;
            reg_file[18387] <= 8'h00;
            reg_file[18388] <= 8'h00;
            reg_file[18389] <= 8'h00;
            reg_file[18390] <= 8'h00;
            reg_file[18391] <= 8'h00;
            reg_file[18392] <= 8'h00;
            reg_file[18393] <= 8'h00;
            reg_file[18394] <= 8'h00;
            reg_file[18395] <= 8'h00;
            reg_file[18396] <= 8'h00;
            reg_file[18397] <= 8'h00;
            reg_file[18398] <= 8'h00;
            reg_file[18399] <= 8'h00;
            reg_file[18400] <= 8'h00;
            reg_file[18401] <= 8'h00;
            reg_file[18402] <= 8'h00;
            reg_file[18403] <= 8'h00;
            reg_file[18404] <= 8'h00;
            reg_file[18405] <= 8'h00;
            reg_file[18406] <= 8'h00;
            reg_file[18407] <= 8'h00;
            reg_file[18408] <= 8'h00;
            reg_file[18409] <= 8'h00;
            reg_file[18410] <= 8'h00;
            reg_file[18411] <= 8'h00;
            reg_file[18412] <= 8'h00;
            reg_file[18413] <= 8'h00;
            reg_file[18414] <= 8'h00;
            reg_file[18415] <= 8'h00;
            reg_file[18416] <= 8'h00;
            reg_file[18417] <= 8'h00;
            reg_file[18418] <= 8'h00;
            reg_file[18419] <= 8'h00;
            reg_file[18420] <= 8'h00;
            reg_file[18421] <= 8'h00;
            reg_file[18422] <= 8'h00;
            reg_file[18423] <= 8'h00;
            reg_file[18424] <= 8'h00;
            reg_file[18425] <= 8'h00;
            reg_file[18426] <= 8'h00;
            reg_file[18427] <= 8'h00;
            reg_file[18428] <= 8'h00;
            reg_file[18429] <= 8'h00;
            reg_file[18430] <= 8'h00;
            reg_file[18431] <= 8'h00;
            reg_file[18432] <= 8'h00;
            reg_file[18433] <= 8'h00;
            reg_file[18434] <= 8'h00;
            reg_file[18435] <= 8'h00;
            reg_file[18436] <= 8'h00;
            reg_file[18437] <= 8'h00;
            reg_file[18438] <= 8'h00;
            reg_file[18439] <= 8'h00;
            reg_file[18440] <= 8'h00;
            reg_file[18441] <= 8'h00;
            reg_file[18442] <= 8'h00;
            reg_file[18443] <= 8'h00;
            reg_file[18444] <= 8'h00;
            reg_file[18445] <= 8'h00;
            reg_file[18446] <= 8'h00;
            reg_file[18447] <= 8'h00;
            reg_file[18448] <= 8'h00;
            reg_file[18449] <= 8'h00;
            reg_file[18450] <= 8'h00;
            reg_file[18451] <= 8'h00;
            reg_file[18452] <= 8'h00;
            reg_file[18453] <= 8'h00;
            reg_file[18454] <= 8'h00;
            reg_file[18455] <= 8'h00;
            reg_file[18456] <= 8'h00;
            reg_file[18457] <= 8'h00;
            reg_file[18458] <= 8'h00;
            reg_file[18459] <= 8'h00;
            reg_file[18460] <= 8'h00;
            reg_file[18461] <= 8'h00;
            reg_file[18462] <= 8'h00;
            reg_file[18463] <= 8'h00;
            reg_file[18464] <= 8'h00;
            reg_file[18465] <= 8'h00;
            reg_file[18466] <= 8'h00;
            reg_file[18467] <= 8'h00;
            reg_file[18468] <= 8'h00;
            reg_file[18469] <= 8'h00;
            reg_file[18470] <= 8'h00;
            reg_file[18471] <= 8'h00;
            reg_file[18472] <= 8'h00;
            reg_file[18473] <= 8'h00;
            reg_file[18474] <= 8'h00;
            reg_file[18475] <= 8'h00;
            reg_file[18476] <= 8'h00;
            reg_file[18477] <= 8'h00;
            reg_file[18478] <= 8'h00;
            reg_file[18479] <= 8'h00;
            reg_file[18480] <= 8'h00;
            reg_file[18481] <= 8'h00;
            reg_file[18482] <= 8'h00;
            reg_file[18483] <= 8'h00;
            reg_file[18484] <= 8'h00;
            reg_file[18485] <= 8'h00;
            reg_file[18486] <= 8'h00;
            reg_file[18487] <= 8'h00;
            reg_file[18488] <= 8'h00;
            reg_file[18489] <= 8'h00;
            reg_file[18490] <= 8'h00;
            reg_file[18491] <= 8'h00;
            reg_file[18492] <= 8'h00;
            reg_file[18493] <= 8'h00;
            reg_file[18494] <= 8'h00;
            reg_file[18495] <= 8'h00;
            reg_file[18496] <= 8'h00;
            reg_file[18497] <= 8'h00;
            reg_file[18498] <= 8'h00;
            reg_file[18499] <= 8'h00;
            reg_file[18500] <= 8'h00;
            reg_file[18501] <= 8'h00;
            reg_file[18502] <= 8'h00;
            reg_file[18503] <= 8'h00;
            reg_file[18504] <= 8'h00;
            reg_file[18505] <= 8'h00;
            reg_file[18506] <= 8'h00;
            reg_file[18507] <= 8'h00;
            reg_file[18508] <= 8'h00;
            reg_file[18509] <= 8'h00;
            reg_file[18510] <= 8'h00;
            reg_file[18511] <= 8'h00;
            reg_file[18512] <= 8'h00;
            reg_file[18513] <= 8'h00;
            reg_file[18514] <= 8'h00;
            reg_file[18515] <= 8'h00;
            reg_file[18516] <= 8'h00;
            reg_file[18517] <= 8'h00;
            reg_file[18518] <= 8'h00;
            reg_file[18519] <= 8'h00;
            reg_file[18520] <= 8'h00;
            reg_file[18521] <= 8'h00;
            reg_file[18522] <= 8'h00;
            reg_file[18523] <= 8'h00;
            reg_file[18524] <= 8'h00;
            reg_file[18525] <= 8'h00;
            reg_file[18526] <= 8'h00;
            reg_file[18527] <= 8'h00;
            reg_file[18528] <= 8'h00;
            reg_file[18529] <= 8'h00;
            reg_file[18530] <= 8'h00;
            reg_file[18531] <= 8'h00;
            reg_file[18532] <= 8'h00;
            reg_file[18533] <= 8'h00;
            reg_file[18534] <= 8'h00;
            reg_file[18535] <= 8'h00;
            reg_file[18536] <= 8'h00;
            reg_file[18537] <= 8'h00;
            reg_file[18538] <= 8'h00;
            reg_file[18539] <= 8'h00;
            reg_file[18540] <= 8'h00;
            reg_file[18541] <= 8'h00;
            reg_file[18542] <= 8'h00;
            reg_file[18543] <= 8'h00;
            reg_file[18544] <= 8'h00;
            reg_file[18545] <= 8'h00;
            reg_file[18546] <= 8'h00;
            reg_file[18547] <= 8'h00;
            reg_file[18548] <= 8'h00;
            reg_file[18549] <= 8'h00;
            reg_file[18550] <= 8'h00;
            reg_file[18551] <= 8'h00;
            reg_file[18552] <= 8'h00;
            reg_file[18553] <= 8'h00;
            reg_file[18554] <= 8'h00;
            reg_file[18555] <= 8'h00;
            reg_file[18556] <= 8'h00;
            reg_file[18557] <= 8'h00;
            reg_file[18558] <= 8'h00;
            reg_file[18559] <= 8'h00;
            reg_file[18560] <= 8'h00;
            reg_file[18561] <= 8'h00;
            reg_file[18562] <= 8'h00;
            reg_file[18563] <= 8'h00;
            reg_file[18564] <= 8'h00;
            reg_file[18565] <= 8'h00;
            reg_file[18566] <= 8'h00;
            reg_file[18567] <= 8'h00;
            reg_file[18568] <= 8'h00;
            reg_file[18569] <= 8'h00;
            reg_file[18570] <= 8'h00;
            reg_file[18571] <= 8'h00;
            reg_file[18572] <= 8'h00;
            reg_file[18573] <= 8'h00;
            reg_file[18574] <= 8'h00;
            reg_file[18575] <= 8'h00;
            reg_file[18576] <= 8'h00;
            reg_file[18577] <= 8'h00;
            reg_file[18578] <= 8'h00;
            reg_file[18579] <= 8'h00;
            reg_file[18580] <= 8'h00;
            reg_file[18581] <= 8'h00;
            reg_file[18582] <= 8'h00;
            reg_file[18583] <= 8'h00;
            reg_file[18584] <= 8'h00;
            reg_file[18585] <= 8'h00;
            reg_file[18586] <= 8'h00;
            reg_file[18587] <= 8'h00;
            reg_file[18588] <= 8'h00;
            reg_file[18589] <= 8'h00;
            reg_file[18590] <= 8'h00;
            reg_file[18591] <= 8'h00;
            reg_file[18592] <= 8'h00;
            reg_file[18593] <= 8'h00;
            reg_file[18594] <= 8'h00;
            reg_file[18595] <= 8'h00;
            reg_file[18596] <= 8'h00;
            reg_file[18597] <= 8'h00;
            reg_file[18598] <= 8'h00;
            reg_file[18599] <= 8'h00;
            reg_file[18600] <= 8'h00;
            reg_file[18601] <= 8'h00;
            reg_file[18602] <= 8'h00;
            reg_file[18603] <= 8'h00;
            reg_file[18604] <= 8'h00;
            reg_file[18605] <= 8'h00;
            reg_file[18606] <= 8'h00;
            reg_file[18607] <= 8'h00;
            reg_file[18608] <= 8'h00;
            reg_file[18609] <= 8'h00;
            reg_file[18610] <= 8'h00;
            reg_file[18611] <= 8'h00;
            reg_file[18612] <= 8'h00;
            reg_file[18613] <= 8'h00;
            reg_file[18614] <= 8'h00;
            reg_file[18615] <= 8'h00;
            reg_file[18616] <= 8'hA4;
            reg_file[18617] <= 8'h01;
            reg_file[18618] <= 8'h00;
            reg_file[18619] <= 8'h80;
            reg_file[18620] <= 8'h00;
            reg_file[18621] <= 8'h00;
            reg_file[18622] <= 8'h00;
            reg_file[18623] <= 8'h00;
            reg_file[18624] <= 8'h00;
            reg_file[18625] <= 8'h00;
            reg_file[18626] <= 8'h00;
            reg_file[18627] <= 8'h00;
            reg_file[18628] <= 8'h00;
            reg_file[18629] <= 8'h00;
            reg_file[18630] <= 8'h00;
            reg_file[18631] <= 8'h00;
            reg_file[18632] <= 8'h00;
            reg_file[18633] <= 8'h00;
            reg_file[18634] <= 8'h00;
            reg_file[18635] <= 8'h00;
            reg_file[18636] <= 8'hB4;
            reg_file[18637] <= 8'h4B;
            reg_file[18638] <= 8'h00;
            reg_file[18639] <= 8'h80;
            reg_file[18640] <= 8'h1C;
            reg_file[18641] <= 8'h4C;
            reg_file[18642] <= 8'h00;
            reg_file[18643] <= 8'h80;
            reg_file[18644] <= 8'h84;
            reg_file[18645] <= 8'h4C;
            reg_file[18646] <= 8'h00;
            reg_file[18647] <= 8'h80;
            reg_file[18648] <= 8'h00;
            reg_file[18649] <= 8'h00;
            reg_file[18650] <= 8'h00;
            reg_file[18651] <= 8'h00;
            reg_file[18652] <= 8'h00;
            reg_file[18653] <= 8'h00;
            reg_file[18654] <= 8'h00;
            reg_file[18655] <= 8'h00;
            reg_file[18656] <= 8'h00;
            reg_file[18657] <= 8'h00;
            reg_file[18658] <= 8'h00;
            reg_file[18659] <= 8'h00;
            reg_file[18660] <= 8'h00;
            reg_file[18661] <= 8'h00;
            reg_file[18662] <= 8'h00;
            reg_file[18663] <= 8'h00;
            reg_file[18664] <= 8'h00;
            reg_file[18665] <= 8'h00;
            reg_file[18666] <= 8'h00;
            reg_file[18667] <= 8'h00;
            reg_file[18668] <= 8'h00;
            reg_file[18669] <= 8'h00;
            reg_file[18670] <= 8'h00;
            reg_file[18671] <= 8'h00;
            reg_file[18672] <= 8'h00;
            reg_file[18673] <= 8'h00;
            reg_file[18674] <= 8'h00;
            reg_file[18675] <= 8'h00;
            reg_file[18676] <= 8'h00;
            reg_file[18677] <= 8'h00;
            reg_file[18678] <= 8'h00;
            reg_file[18679] <= 8'h00;
            reg_file[18680] <= 8'h00;
            reg_file[18681] <= 8'h00;
            reg_file[18682] <= 8'h00;
            reg_file[18683] <= 8'h00;
            reg_file[18684] <= 8'h00;
            reg_file[18685] <= 8'h00;
            reg_file[18686] <= 8'h00;
            reg_file[18687] <= 8'h00;
            reg_file[18688] <= 8'h00;
            reg_file[18689] <= 8'h00;
            reg_file[18690] <= 8'h00;
            reg_file[18691] <= 8'h00;
            reg_file[18692] <= 8'h00;
            reg_file[18693] <= 8'h00;
            reg_file[18694] <= 8'h00;
            reg_file[18695] <= 8'h00;
            reg_file[18696] <= 8'h00;
            reg_file[18697] <= 8'h00;
            reg_file[18698] <= 8'h00;
            reg_file[18699] <= 8'h00;
            reg_file[18700] <= 8'h00;
            reg_file[18701] <= 8'h00;
            reg_file[18702] <= 8'h00;
            reg_file[18703] <= 8'h00;
            reg_file[18704] <= 8'h00;
            reg_file[18705] <= 8'h00;
            reg_file[18706] <= 8'h00;
            reg_file[18707] <= 8'h00;
            reg_file[18708] <= 8'h00;
            reg_file[18709] <= 8'h00;
            reg_file[18710] <= 8'h00;
            reg_file[18711] <= 8'h00;
            reg_file[18712] <= 8'h00;
            reg_file[18713] <= 8'h00;
            reg_file[18714] <= 8'h00;
            reg_file[18715] <= 8'h00;
            reg_file[18716] <= 8'h00;
            reg_file[18717] <= 8'h00;
            reg_file[18718] <= 8'h00;
            reg_file[18719] <= 8'h00;
            reg_file[18720] <= 8'h00;
            reg_file[18721] <= 8'h00;
            reg_file[18722] <= 8'h00;
            reg_file[18723] <= 8'h00;
            reg_file[18724] <= 8'h00;
            reg_file[18725] <= 8'h00;
            reg_file[18726] <= 8'h00;
            reg_file[18727] <= 8'h00;
            reg_file[18728] <= 8'h00;
            reg_file[18729] <= 8'h00;
            reg_file[18730] <= 8'h00;
            reg_file[18731] <= 8'h00;
            reg_file[18732] <= 8'h00;
            reg_file[18733] <= 8'h00;
            reg_file[18734] <= 8'h00;
            reg_file[18735] <= 8'h00;
            reg_file[18736] <= 8'h00;
            reg_file[18737] <= 8'h00;
            reg_file[18738] <= 8'h00;
            reg_file[18739] <= 8'h00;
            reg_file[18740] <= 8'h00;
            reg_file[18741] <= 8'h00;
            reg_file[18742] <= 8'h00;
            reg_file[18743] <= 8'h00;
            reg_file[18744] <= 8'h00;
            reg_file[18745] <= 8'h00;
            reg_file[18746] <= 8'h00;
            reg_file[18747] <= 8'h00;
            reg_file[18748] <= 8'h00;
            reg_file[18749] <= 8'h00;
            reg_file[18750] <= 8'h00;
            reg_file[18751] <= 8'h00;
            reg_file[18752] <= 8'h00;
            reg_file[18753] <= 8'h00;
            reg_file[18754] <= 8'h00;
            reg_file[18755] <= 8'h00;
            reg_file[18756] <= 8'h00;
            reg_file[18757] <= 8'h00;
            reg_file[18758] <= 8'h00;
            reg_file[18759] <= 8'h00;
            reg_file[18760] <= 8'h00;
            reg_file[18761] <= 8'h00;
            reg_file[18762] <= 8'h00;
            reg_file[18763] <= 8'h00;
            reg_file[18764] <= 8'h00;
            reg_file[18765] <= 8'h00;
            reg_file[18766] <= 8'h00;
            reg_file[18767] <= 8'h00;
            reg_file[18768] <= 8'h00;
            reg_file[18769] <= 8'h00;
            reg_file[18770] <= 8'h00;
            reg_file[18771] <= 8'h00;
            reg_file[18772] <= 8'h00;
            reg_file[18773] <= 8'h00;
            reg_file[18774] <= 8'h00;
            reg_file[18775] <= 8'h00;
            reg_file[18776] <= 8'h00;
            reg_file[18777] <= 8'h00;
            reg_file[18778] <= 8'h00;
            reg_file[18779] <= 8'h00;
            reg_file[18780] <= 8'h00;
            reg_file[18781] <= 8'h00;
            reg_file[18782] <= 8'h00;
            reg_file[18783] <= 8'h00;
            reg_file[18784] <= 8'h00;
            reg_file[18785] <= 8'h00;
            reg_file[18786] <= 8'h00;
            reg_file[18787] <= 8'h00;
            reg_file[18788] <= 8'h00;
            reg_file[18789] <= 8'h00;
            reg_file[18790] <= 8'h00;
            reg_file[18791] <= 8'h00;
            reg_file[18792] <= 8'h00;
            reg_file[18793] <= 8'h00;
            reg_file[18794] <= 8'h00;
            reg_file[18795] <= 8'h00;
            reg_file[18796] <= 8'h00;
            reg_file[18797] <= 8'h00;
            reg_file[18798] <= 8'h00;
            reg_file[18799] <= 8'h00;
            reg_file[18800] <= 8'h01;
            reg_file[18801] <= 8'h00;
            reg_file[18802] <= 8'h00;
            reg_file[18803] <= 8'h00;
            reg_file[18804] <= 8'h00;
            reg_file[18805] <= 8'h00;
            reg_file[18806] <= 8'h00;
            reg_file[18807] <= 8'h00;
            reg_file[18808] <= 8'h0E;
            reg_file[18809] <= 8'h33;
            reg_file[18810] <= 8'hCD;
            reg_file[18811] <= 8'hAB;
            reg_file[18812] <= 8'h34;
            reg_file[18813] <= 8'h12;
            reg_file[18814] <= 8'h6D;
            reg_file[18815] <= 8'hE6;
            reg_file[18816] <= 8'hEC;
            reg_file[18817] <= 8'hDE;
            reg_file[18818] <= 8'h05;
            reg_file[18819] <= 8'h00;
            reg_file[18820] <= 8'h0B;
            reg_file[18821] <= 8'h00;
            reg_file[18822] <= 8'h00;
            reg_file[18823] <= 8'h00;
            reg_file[18824] <= 8'h00;
            reg_file[18825] <= 8'h00;
            reg_file[18826] <= 8'h00;
            reg_file[18827] <= 8'h00;
            reg_file[18828] <= 8'h00;
            reg_file[18829] <= 8'h00;
            reg_file[18830] <= 8'h00;
            reg_file[18831] <= 8'h00;
            reg_file[18832] <= 8'h00;
            reg_file[18833] <= 8'h00;
            reg_file[18834] <= 8'h00;
            reg_file[18835] <= 8'h00;
            reg_file[18836] <= 8'h00;
            reg_file[18837] <= 8'h00;
            reg_file[18838] <= 8'h00;
            reg_file[18839] <= 8'h00;
            reg_file[18840] <= 8'h00;
            reg_file[18841] <= 8'h00;
            reg_file[18842] <= 8'h00;
            reg_file[18843] <= 8'h00;
            reg_file[18844] <= 8'h00;
            reg_file[18845] <= 8'h00;
            reg_file[18846] <= 8'h00;
            reg_file[18847] <= 8'h00;
            reg_file[18848] <= 8'h00;
            reg_file[18849] <= 8'h00;
            reg_file[18850] <= 8'h00;
            reg_file[18851] <= 8'h00;
            reg_file[18852] <= 8'h00;
            reg_file[18853] <= 8'h00;
            reg_file[18854] <= 8'h00;
            reg_file[18855] <= 8'h00;
            reg_file[18856] <= 8'h00;
            reg_file[18857] <= 8'h00;
            reg_file[18858] <= 8'h00;
            reg_file[18859] <= 8'h00;
            reg_file[18860] <= 8'h00;
            reg_file[18861] <= 8'h00;
            reg_file[18862] <= 8'h00;
            reg_file[18863] <= 8'h00;
            reg_file[18864] <= 8'h00;
            reg_file[18865] <= 8'h00;
            reg_file[18866] <= 8'h00;
            reg_file[18867] <= 8'h00;
            reg_file[18868] <= 8'h00;
            reg_file[18869] <= 8'h00;
            reg_file[18870] <= 8'h00;
            reg_file[18871] <= 8'h00;
            reg_file[18872] <= 8'h00;
            reg_file[18873] <= 8'h00;
            reg_file[18874] <= 8'h00;
            reg_file[18875] <= 8'h00;
            reg_file[18876] <= 8'h00;
            reg_file[18877] <= 8'h00;
            reg_file[18878] <= 8'h00;
            reg_file[18879] <= 8'h00;
            reg_file[18880] <= 8'h00;
            reg_file[18881] <= 8'h00;
            reg_file[18882] <= 8'h00;
            reg_file[18883] <= 8'h00;
            reg_file[18884] <= 8'h00;
            reg_file[18885] <= 8'h00;
            reg_file[18886] <= 8'h00;
            reg_file[18887] <= 8'h00;
            reg_file[18888] <= 8'h00;
            reg_file[18889] <= 8'h00;
            reg_file[18890] <= 8'h00;
            reg_file[18891] <= 8'h00;
            reg_file[18892] <= 8'h00;
            reg_file[18893] <= 8'h00;
            reg_file[18894] <= 8'h00;
            reg_file[18895] <= 8'h00;
            reg_file[18896] <= 8'h00;
            reg_file[18897] <= 8'h00;
            reg_file[18898] <= 8'h00;
            reg_file[18899] <= 8'h00;
            reg_file[18900] <= 8'h00;
            reg_file[18901] <= 8'h00;
            reg_file[18902] <= 8'h00;
            reg_file[18903] <= 8'h00;
            reg_file[18904] <= 8'h00;
            reg_file[18905] <= 8'h00;
            reg_file[18906] <= 8'h00;
            reg_file[18907] <= 8'h00;
            reg_file[18908] <= 8'h00;
            reg_file[18909] <= 8'h00;
            reg_file[18910] <= 8'h00;
            reg_file[18911] <= 8'h00;
            reg_file[18912] <= 8'h00;
            reg_file[18913] <= 8'h00;
            reg_file[18914] <= 8'h00;
            reg_file[18915] <= 8'h00;
            reg_file[18916] <= 8'h00;
            reg_file[18917] <= 8'h00;
            reg_file[18918] <= 8'h00;
            reg_file[18919] <= 8'h00;
            reg_file[18920] <= 8'h00;
            reg_file[18921] <= 8'h00;
            reg_file[18922] <= 8'h00;
            reg_file[18923] <= 8'h00;
            reg_file[18924] <= 8'h00;
            reg_file[18925] <= 8'h00;
            reg_file[18926] <= 8'h00;
            reg_file[18927] <= 8'h00;
            reg_file[18928] <= 8'h00;
            reg_file[18929] <= 8'h00;
            reg_file[18930] <= 8'h00;
            reg_file[18931] <= 8'h00;
            reg_file[18932] <= 8'h00;
            reg_file[18933] <= 8'h00;
            reg_file[18934] <= 8'h00;
            reg_file[18935] <= 8'h00;
            reg_file[18936] <= 8'h00;
            reg_file[18937] <= 8'h00;
            reg_file[18938] <= 8'h00;
            reg_file[18939] <= 8'h00;
            reg_file[18940] <= 8'h00;
            reg_file[18941] <= 8'h00;
            reg_file[18942] <= 8'h00;
            reg_file[18943] <= 8'h00;
            reg_file[18944] <= 8'h00;
            reg_file[18945] <= 8'h00;
            reg_file[18946] <= 8'h00;
            reg_file[18947] <= 8'h00;
            reg_file[18948] <= 8'h00;
            reg_file[18949] <= 8'h00;
            reg_file[18950] <= 8'h00;
            reg_file[18951] <= 8'h00;
            reg_file[18952] <= 8'h00;
            reg_file[18953] <= 8'h00;
            reg_file[18954] <= 8'h00;
            reg_file[18955] <= 8'h00;
            reg_file[18956] <= 8'h00;
            reg_file[18957] <= 8'h00;
            reg_file[18958] <= 8'h00;
            reg_file[18959] <= 8'h00;
            reg_file[18960] <= 8'h00;
            reg_file[18961] <= 8'h00;
            reg_file[18962] <= 8'h00;
            reg_file[18963] <= 8'h00;
            reg_file[18964] <= 8'h00;
            reg_file[18965] <= 8'h00;
            reg_file[18966] <= 8'h00;
            reg_file[18967] <= 8'h00;
            reg_file[18968] <= 8'h00;
            reg_file[18969] <= 8'h00;
            reg_file[18970] <= 8'h00;
            reg_file[18971] <= 8'h00;
            reg_file[18972] <= 8'h00;
            reg_file[18973] <= 8'h00;
            reg_file[18974] <= 8'h00;
            reg_file[18975] <= 8'h00;
            reg_file[18976] <= 8'h00;
            reg_file[18977] <= 8'h00;
            reg_file[18978] <= 8'h00;
            reg_file[18979] <= 8'h00;
            reg_file[18980] <= 8'h00;
            reg_file[18981] <= 8'h00;
            reg_file[18982] <= 8'h00;
            reg_file[18983] <= 8'h00;
            reg_file[18984] <= 8'h00;
            reg_file[18985] <= 8'h00;
            reg_file[18986] <= 8'h00;
            reg_file[18987] <= 8'h00;
            reg_file[18988] <= 8'h00;
            reg_file[18989] <= 8'h00;
            reg_file[18990] <= 8'h00;
            reg_file[18991] <= 8'h00;
            reg_file[18992] <= 8'h00;
            reg_file[18993] <= 8'h00;
            reg_file[18994] <= 8'h00;
            reg_file[18995] <= 8'h00;
            reg_file[18996] <= 8'h00;
            reg_file[18997] <= 8'h00;
            reg_file[18998] <= 8'h00;
            reg_file[18999] <= 8'h00;
            reg_file[19000] <= 8'h00;
            reg_file[19001] <= 8'h00;
            reg_file[19002] <= 8'h00;
            reg_file[19003] <= 8'h00;
            reg_file[19004] <= 8'h00;
            reg_file[19005] <= 8'h00;
            reg_file[19006] <= 8'h00;
            reg_file[19007] <= 8'h00;
            reg_file[19008] <= 8'h00;
            reg_file[19009] <= 8'h00;
            reg_file[19010] <= 8'h00;
            reg_file[19011] <= 8'h00;
            reg_file[19012] <= 8'h00;
            reg_file[19013] <= 8'h00;
            reg_file[19014] <= 8'h00;
            reg_file[19015] <= 8'h00;
            reg_file[19016] <= 8'h00;
            reg_file[19017] <= 8'h00;
            reg_file[19018] <= 8'h00;
            reg_file[19019] <= 8'h00;
            reg_file[19020] <= 8'h00;
            reg_file[19021] <= 8'h00;
            reg_file[19022] <= 8'h00;
            reg_file[19023] <= 8'h00;
            reg_file[19024] <= 8'h00;
            reg_file[19025] <= 8'h00;
            reg_file[19026] <= 8'h00;
            reg_file[19027] <= 8'h00;
            reg_file[19028] <= 8'h00;
            reg_file[19029] <= 8'h00;
            reg_file[19030] <= 8'h00;
            reg_file[19031] <= 8'h00;
            reg_file[19032] <= 8'h00;
            reg_file[19033] <= 8'h00;
            reg_file[19034] <= 8'h00;
            reg_file[19035] <= 8'h00;
            reg_file[19036] <= 8'h00;
            reg_file[19037] <= 8'h00;
            reg_file[19038] <= 8'h00;
            reg_file[19039] <= 8'h00;
            reg_file[19040] <= 8'h00;
            reg_file[19041] <= 8'h00;
            reg_file[19042] <= 8'h00;
            reg_file[19043] <= 8'h00;
            reg_file[19044] <= 8'h00;
            reg_file[19045] <= 8'h00;
            reg_file[19046] <= 8'h00;
            reg_file[19047] <= 8'h00;
            reg_file[19048] <= 8'h00;
            reg_file[19049] <= 8'h00;
            reg_file[19050] <= 8'h00;
            reg_file[19051] <= 8'h00;
            reg_file[19052] <= 8'h00;
            reg_file[19053] <= 8'h00;
            reg_file[19054] <= 8'h00;
            reg_file[19055] <= 8'h00;
            reg_file[19056] <= 8'h00;
            reg_file[19057] <= 8'h00;
            reg_file[19058] <= 8'h00;
            reg_file[19059] <= 8'h00;
            reg_file[19060] <= 8'h00;
            reg_file[19061] <= 8'h00;
            reg_file[19062] <= 8'h00;
            reg_file[19063] <= 8'h00;
            reg_file[19064] <= 8'h00;
            reg_file[19065] <= 8'h00;
            reg_file[19066] <= 8'h00;
            reg_file[19067] <= 8'h00;
            reg_file[19068] <= 8'h00;
            reg_file[19069] <= 8'h00;
            reg_file[19070] <= 8'h00;
            reg_file[19071] <= 8'h00;
            reg_file[19072] <= 8'h00;
            reg_file[19073] <= 8'h00;
            reg_file[19074] <= 8'h00;
            reg_file[19075] <= 8'h00;
            reg_file[19076] <= 8'h00;
            reg_file[19077] <= 8'h00;
            reg_file[19078] <= 8'h00;
            reg_file[19079] <= 8'h00;
            reg_file[19080] <= 8'h00;
            reg_file[19081] <= 8'h00;
            reg_file[19082] <= 8'h00;
            reg_file[19083] <= 8'h00;
            reg_file[19084] <= 8'h00;
            reg_file[19085] <= 8'h00;
            reg_file[19086] <= 8'h00;
            reg_file[19087] <= 8'h00;
            reg_file[19088] <= 8'h00;
            reg_file[19089] <= 8'h00;
            reg_file[19090] <= 8'h00;
            reg_file[19091] <= 8'h00;
            reg_file[19092] <= 8'h00;
            reg_file[19093] <= 8'h00;
            reg_file[19094] <= 8'h00;
            reg_file[19095] <= 8'h00;
            reg_file[19096] <= 8'h00;
            reg_file[19097] <= 8'h00;
            reg_file[19098] <= 8'h00;
            reg_file[19099] <= 8'h00;
            reg_file[19100] <= 8'h00;
            reg_file[19101] <= 8'h00;
            reg_file[19102] <= 8'h00;
            reg_file[19103] <= 8'h00;
            reg_file[19104] <= 8'h00;
            reg_file[19105] <= 8'h00;
            reg_file[19106] <= 8'h00;
            reg_file[19107] <= 8'h00;
            reg_file[19108] <= 8'h00;
            reg_file[19109] <= 8'h00;
            reg_file[19110] <= 8'h00;
            reg_file[19111] <= 8'h00;
            reg_file[19112] <= 8'h00;
            reg_file[19113] <= 8'h00;
            reg_file[19114] <= 8'h00;
            reg_file[19115] <= 8'h00;
            reg_file[19116] <= 8'h00;
            reg_file[19117] <= 8'h00;
            reg_file[19118] <= 8'h00;
            reg_file[19119] <= 8'h00;
            reg_file[19120] <= 8'h00;
            reg_file[19121] <= 8'h00;
            reg_file[19122] <= 8'h00;
            reg_file[19123] <= 8'h00;
            reg_file[19124] <= 8'h00;
            reg_file[19125] <= 8'h00;
            reg_file[19126] <= 8'h00;
            reg_file[19127] <= 8'h00;
            reg_file[19128] <= 8'h00;
            reg_file[19129] <= 8'h00;
            reg_file[19130] <= 8'h00;
            reg_file[19131] <= 8'h00;
            reg_file[19132] <= 8'h00;
            reg_file[19133] <= 8'h00;
            reg_file[19134] <= 8'h00;
            reg_file[19135] <= 8'h00;
            reg_file[19136] <= 8'h00;
            reg_file[19137] <= 8'h00;
            reg_file[19138] <= 8'h00;
            reg_file[19139] <= 8'h00;
            reg_file[19140] <= 8'h00;
            reg_file[19141] <= 8'h00;
            reg_file[19142] <= 8'h00;
            reg_file[19143] <= 8'h00;
            reg_file[19144] <= 8'h00;
            reg_file[19145] <= 8'h00;
            reg_file[19146] <= 8'h00;
            reg_file[19147] <= 8'h00;
            reg_file[19148] <= 8'h00;
            reg_file[19149] <= 8'h00;
            reg_file[19150] <= 8'h00;
            reg_file[19151] <= 8'h00;
            reg_file[19152] <= 8'h00;
            reg_file[19153] <= 8'h00;
            reg_file[19154] <= 8'h00;
            reg_file[19155] <= 8'h00;
            reg_file[19156] <= 8'h00;
            reg_file[19157] <= 8'h00;
            reg_file[19158] <= 8'h00;
            reg_file[19159] <= 8'h00;
            reg_file[19160] <= 8'h00;
            reg_file[19161] <= 8'h00;
            reg_file[19162] <= 8'h00;
            reg_file[19163] <= 8'h00;
            reg_file[19164] <= 8'h00;
            reg_file[19165] <= 8'h00;
            reg_file[19166] <= 8'h00;
            reg_file[19167] <= 8'h00;
            reg_file[19168] <= 8'h00;
            reg_file[19169] <= 8'h00;
            reg_file[19170] <= 8'h00;
            reg_file[19171] <= 8'h00;
            reg_file[19172] <= 8'h00;
            reg_file[19173] <= 8'h00;
            reg_file[19174] <= 8'h00;
            reg_file[19175] <= 8'h00;
            reg_file[19176] <= 8'h00;
            reg_file[19177] <= 8'h00;
            reg_file[19178] <= 8'h00;
            reg_file[19179] <= 8'h00;
            reg_file[19180] <= 8'h00;
            reg_file[19181] <= 8'h00;
            reg_file[19182] <= 8'h00;
            reg_file[19183] <= 8'h00;
            reg_file[19184] <= 8'h00;
            reg_file[19185] <= 8'h00;
            reg_file[19186] <= 8'h00;
            reg_file[19187] <= 8'h00;
            reg_file[19188] <= 8'h00;
            reg_file[19189] <= 8'h00;
            reg_file[19190] <= 8'h00;
            reg_file[19191] <= 8'h00;
            reg_file[19192] <= 8'h00;
            reg_file[19193] <= 8'h00;
            reg_file[19194] <= 8'h00;
            reg_file[19195] <= 8'h00;
            reg_file[19196] <= 8'h00;
            reg_file[19197] <= 8'h00;
            reg_file[19198] <= 8'h00;
            reg_file[19199] <= 8'h00;
            reg_file[19200] <= 8'h00;
            reg_file[19201] <= 8'h00;
            reg_file[19202] <= 8'h00;
            reg_file[19203] <= 8'h00;
            reg_file[19204] <= 8'h00;
            reg_file[19205] <= 8'h00;
            reg_file[19206] <= 8'h00;
            reg_file[19207] <= 8'h00;
            reg_file[19208] <= 8'h00;
            reg_file[19209] <= 8'h00;
            reg_file[19210] <= 8'h00;
            reg_file[19211] <= 8'h00;
            reg_file[19212] <= 8'h00;
            reg_file[19213] <= 8'h00;
            reg_file[19214] <= 8'h00;
            reg_file[19215] <= 8'h00;
            reg_file[19216] <= 8'h00;
            reg_file[19217] <= 8'h00;
            reg_file[19218] <= 8'h00;
            reg_file[19219] <= 8'h00;
            reg_file[19220] <= 8'h00;
            reg_file[19221] <= 8'h00;
            reg_file[19222] <= 8'h00;
            reg_file[19223] <= 8'h00;
            reg_file[19224] <= 8'h00;
            reg_file[19225] <= 8'h00;
            reg_file[19226] <= 8'h00;
            reg_file[19227] <= 8'h00;
            reg_file[19228] <= 8'h00;
            reg_file[19229] <= 8'h00;
            reg_file[19230] <= 8'h00;
            reg_file[19231] <= 8'h00;
            reg_file[19232] <= 8'h00;
            reg_file[19233] <= 8'h00;
            reg_file[19234] <= 8'h00;
            reg_file[19235] <= 8'h00;
            reg_file[19236] <= 8'h00;
            reg_file[19237] <= 8'h00;
            reg_file[19238] <= 8'h00;
            reg_file[19239] <= 8'h00;
            reg_file[19240] <= 8'h00;
            reg_file[19241] <= 8'h00;
            reg_file[19242] <= 8'h00;
            reg_file[19243] <= 8'h00;
            reg_file[19244] <= 8'h00;
            reg_file[19245] <= 8'h00;
            reg_file[19246] <= 8'h00;
            reg_file[19247] <= 8'h00;
            reg_file[19248] <= 8'h00;
            reg_file[19249] <= 8'h00;
            reg_file[19250] <= 8'h00;
            reg_file[19251] <= 8'h00;
            reg_file[19252] <= 8'h00;
            reg_file[19253] <= 8'h00;
            reg_file[19254] <= 8'h00;
            reg_file[19255] <= 8'h00;
            reg_file[19256] <= 8'h00;
            reg_file[19257] <= 8'h00;
            reg_file[19258] <= 8'h00;
            reg_file[19259] <= 8'h00;
            reg_file[19260] <= 8'h00;
            reg_file[19261] <= 8'h00;
            reg_file[19262] <= 8'h00;
            reg_file[19263] <= 8'h00;
            reg_file[19264] <= 8'h00;
            reg_file[19265] <= 8'h00;
            reg_file[19266] <= 8'h00;
            reg_file[19267] <= 8'h00;
            reg_file[19268] <= 8'h00;
            reg_file[19269] <= 8'h00;
            reg_file[19270] <= 8'h00;
            reg_file[19271] <= 8'h00;
            reg_file[19272] <= 8'h00;
            reg_file[19273] <= 8'h00;
            reg_file[19274] <= 8'h00;
            reg_file[19275] <= 8'h00;
            reg_file[19276] <= 8'h00;
            reg_file[19277] <= 8'h00;
            reg_file[19278] <= 8'h00;
            reg_file[19279] <= 8'h00;
            reg_file[19280] <= 8'h00;
            reg_file[19281] <= 8'h00;
            reg_file[19282] <= 8'h00;
            reg_file[19283] <= 8'h00;
            reg_file[19284] <= 8'h00;
            reg_file[19285] <= 8'h00;
            reg_file[19286] <= 8'h00;
            reg_file[19287] <= 8'h00;
            reg_file[19288] <= 8'h00;
            reg_file[19289] <= 8'h00;
            reg_file[19290] <= 8'h00;
            reg_file[19291] <= 8'h00;
            reg_file[19292] <= 8'h00;
            reg_file[19293] <= 8'h00;
            reg_file[19294] <= 8'h00;
            reg_file[19295] <= 8'h00;
            reg_file[19296] <= 8'h00;
            reg_file[19297] <= 8'h00;
            reg_file[19298] <= 8'h00;
            reg_file[19299] <= 8'h00;
            reg_file[19300] <= 8'h00;
            reg_file[19301] <= 8'h00;
            reg_file[19302] <= 8'h00;
            reg_file[19303] <= 8'h00;
            reg_file[19304] <= 8'h00;
            reg_file[19305] <= 8'h00;
            reg_file[19306] <= 8'h00;
            reg_file[19307] <= 8'h00;
            reg_file[19308] <= 8'h00;
            reg_file[19309] <= 8'h00;
            reg_file[19310] <= 8'h00;
            reg_file[19311] <= 8'h00;
            reg_file[19312] <= 8'h00;
            reg_file[19313] <= 8'h00;
            reg_file[19314] <= 8'h00;
            reg_file[19315] <= 8'h00;
            reg_file[19316] <= 8'h00;
            reg_file[19317] <= 8'h00;
            reg_file[19318] <= 8'h00;
            reg_file[19319] <= 8'h00;
            reg_file[19320] <= 8'h00;
            reg_file[19321] <= 8'h00;
            reg_file[19322] <= 8'h00;
            reg_file[19323] <= 8'h00;
            reg_file[19324] <= 8'h00;
            reg_file[19325] <= 8'h00;
            reg_file[19326] <= 8'h00;
            reg_file[19327] <= 8'h00;
            reg_file[19328] <= 8'h00;
            reg_file[19329] <= 8'h00;
            reg_file[19330] <= 8'h00;
            reg_file[19331] <= 8'h00;
            reg_file[19332] <= 8'h00;
            reg_file[19333] <= 8'h00;
            reg_file[19334] <= 8'h00;
            reg_file[19335] <= 8'h00;
            reg_file[19336] <= 8'h00;
            reg_file[19337] <= 8'h00;
            reg_file[19338] <= 8'h00;
            reg_file[19339] <= 8'h00;
            reg_file[19340] <= 8'h00;
            reg_file[19341] <= 8'h00;
            reg_file[19342] <= 8'h00;
            reg_file[19343] <= 8'h00;
            reg_file[19344] <= 8'h00;
            reg_file[19345] <= 8'h00;
            reg_file[19346] <= 8'h00;
            reg_file[19347] <= 8'h00;
            reg_file[19348] <= 8'h00;
            reg_file[19349] <= 8'h00;
            reg_file[19350] <= 8'h00;
            reg_file[19351] <= 8'h00;
            reg_file[19352] <= 8'h00;
            reg_file[19353] <= 8'h00;
            reg_file[19354] <= 8'h00;
            reg_file[19355] <= 8'h00;
            reg_file[19356] <= 8'h00;
            reg_file[19357] <= 8'h00;
            reg_file[19358] <= 8'h00;
            reg_file[19359] <= 8'h00;
            reg_file[19360] <= 8'h00;
            reg_file[19361] <= 8'h00;
            reg_file[19362] <= 8'h00;
            reg_file[19363] <= 8'h00;
            reg_file[19364] <= 8'h00;
            reg_file[19365] <= 8'h00;
            reg_file[19366] <= 8'h00;
            reg_file[19367] <= 8'h00;
            reg_file[19368] <= 8'h00;
            reg_file[19369] <= 8'h00;
            reg_file[19370] <= 8'h00;
            reg_file[19371] <= 8'h00;
            reg_file[19372] <= 8'h00;
            reg_file[19373] <= 8'h00;
            reg_file[19374] <= 8'h00;
            reg_file[19375] <= 8'h00;
            reg_file[19376] <= 8'h00;
            reg_file[19377] <= 8'h00;
            reg_file[19378] <= 8'h00;
            reg_file[19379] <= 8'h00;
            reg_file[19380] <= 8'h00;
            reg_file[19381] <= 8'h00;
            reg_file[19382] <= 8'h00;
            reg_file[19383] <= 8'h00;
            reg_file[19384] <= 8'h00;
            reg_file[19385] <= 8'h00;
            reg_file[19386] <= 8'h00;
            reg_file[19387] <= 8'h00;
            reg_file[19388] <= 8'h00;
            reg_file[19389] <= 8'h00;
            reg_file[19390] <= 8'h00;
            reg_file[19391] <= 8'h00;
            reg_file[19392] <= 8'h00;
            reg_file[19393] <= 8'h00;
            reg_file[19394] <= 8'h00;
            reg_file[19395] <= 8'h00;
            reg_file[19396] <= 8'h00;
            reg_file[19397] <= 8'h00;
            reg_file[19398] <= 8'h00;
            reg_file[19399] <= 8'h00;
            reg_file[19400] <= 8'h00;
            reg_file[19401] <= 8'h00;
            reg_file[19402] <= 8'h00;
            reg_file[19403] <= 8'h00;
            reg_file[19404] <= 8'h00;
            reg_file[19405] <= 8'h00;
            reg_file[19406] <= 8'h00;
            reg_file[19407] <= 8'h00;
            reg_file[19408] <= 8'h00;
            reg_file[19409] <= 8'h00;
            reg_file[19410] <= 8'h00;
            reg_file[19411] <= 8'h00;
            reg_file[19412] <= 8'h00;
            reg_file[19413] <= 8'h00;
            reg_file[19414] <= 8'h00;
            reg_file[19415] <= 8'h00;
            reg_file[19416] <= 8'h00;
            reg_file[19417] <= 8'h00;
            reg_file[19418] <= 8'h00;
            reg_file[19419] <= 8'h00;
            reg_file[19420] <= 8'h00;
            reg_file[19421] <= 8'h00;
            reg_file[19422] <= 8'h00;
            reg_file[19423] <= 8'h00;
            reg_file[19424] <= 8'h00;
            reg_file[19425] <= 8'h00;
            reg_file[19426] <= 8'h00;
            reg_file[19427] <= 8'h00;
            reg_file[19428] <= 8'h00;
            reg_file[19429] <= 8'h00;
            reg_file[19430] <= 8'h00;
            reg_file[19431] <= 8'h00;
            reg_file[19432] <= 8'h00;
            reg_file[19433] <= 8'h00;
            reg_file[19434] <= 8'h00;
            reg_file[19435] <= 8'h00;
            reg_file[19436] <= 8'h00;
            reg_file[19437] <= 8'h00;
            reg_file[19438] <= 8'h00;
            reg_file[19439] <= 8'h00;
            reg_file[19440] <= 8'h00;
            reg_file[19441] <= 8'h00;
            reg_file[19442] <= 8'h00;
            reg_file[19443] <= 8'h00;
            reg_file[19444] <= 8'h00;
            reg_file[19445] <= 8'h00;
            reg_file[19446] <= 8'h00;
            reg_file[19447] <= 8'h00;
            reg_file[19448] <= 8'h00;
            reg_file[19449] <= 8'h00;
            reg_file[19450] <= 8'h00;
            reg_file[19451] <= 8'h00;
            reg_file[19452] <= 8'h00;
            reg_file[19453] <= 8'h00;
            reg_file[19454] <= 8'h00;
            reg_file[19455] <= 8'h00;
            reg_file[19456] <= 8'h00;
            reg_file[19457] <= 8'h00;
            reg_file[19458] <= 8'h00;
            reg_file[19459] <= 8'h00;
            reg_file[19460] <= 8'h00;
            reg_file[19461] <= 8'h00;
            reg_file[19462] <= 8'h00;
            reg_file[19463] <= 8'h00;
            reg_file[19464] <= 8'h00;
            reg_file[19465] <= 8'h00;
            reg_file[19466] <= 8'h00;
            reg_file[19467] <= 8'h00;
            reg_file[19468] <= 8'h00;
            reg_file[19469] <= 8'h00;
            reg_file[19470] <= 8'h00;
            reg_file[19471] <= 8'h00;
            reg_file[19472] <= 8'h00;
            reg_file[19473] <= 8'h00;
            reg_file[19474] <= 8'h00;
            reg_file[19475] <= 8'h00;
            reg_file[19476] <= 8'h00;
            reg_file[19477] <= 8'h00;
            reg_file[19478] <= 8'h00;
            reg_file[19479] <= 8'h00;
            reg_file[19480] <= 8'h00;
            reg_file[19481] <= 8'h00;
            reg_file[19482] <= 8'h00;
            reg_file[19483] <= 8'h00;
            reg_file[19484] <= 8'h00;
            reg_file[19485] <= 8'h00;
            reg_file[19486] <= 8'h00;
            reg_file[19487] <= 8'h00;
            reg_file[19488] <= 8'h00;
            reg_file[19489] <= 8'h00;
            reg_file[19490] <= 8'h00;
            reg_file[19491] <= 8'h00;
            reg_file[19492] <= 8'h00;
            reg_file[19493] <= 8'h00;
            reg_file[19494] <= 8'h00;
            reg_file[19495] <= 8'h00;
            reg_file[19496] <= 8'h00;
            reg_file[19497] <= 8'h00;
            reg_file[19498] <= 8'h00;
            reg_file[19499] <= 8'h00;
            reg_file[19500] <= 8'h00;
            reg_file[19501] <= 8'h00;
            reg_file[19502] <= 8'h00;
            reg_file[19503] <= 8'h00;
            reg_file[19504] <= 8'h00;
            reg_file[19505] <= 8'h00;
            reg_file[19506] <= 8'h00;
            reg_file[19507] <= 8'h00;
            reg_file[19508] <= 8'h00;
            reg_file[19509] <= 8'h00;
            reg_file[19510] <= 8'h00;
            reg_file[19511] <= 8'h00;
            reg_file[19512] <= 8'h00;
            reg_file[19513] <= 8'h00;
            reg_file[19514] <= 8'h00;
            reg_file[19515] <= 8'h00;
            reg_file[19516] <= 8'h00;
            reg_file[19517] <= 8'h00;
            reg_file[19518] <= 8'h00;
            reg_file[19519] <= 8'h00;
            reg_file[19520] <= 8'h00;
            reg_file[19521] <= 8'h00;
            reg_file[19522] <= 8'h00;
            reg_file[19523] <= 8'h00;
            reg_file[19524] <= 8'h00;
            reg_file[19525] <= 8'h00;
            reg_file[19526] <= 8'h00;
            reg_file[19527] <= 8'h00;
            reg_file[19528] <= 8'h00;
            reg_file[19529] <= 8'h00;
            reg_file[19530] <= 8'h00;
            reg_file[19531] <= 8'h00;
            reg_file[19532] <= 8'h00;
            reg_file[19533] <= 8'h00;
            reg_file[19534] <= 8'h00;
            reg_file[19535] <= 8'h00;
            reg_file[19536] <= 8'h00;
            reg_file[19537] <= 8'h00;
            reg_file[19538] <= 8'h00;
            reg_file[19539] <= 8'h00;
            reg_file[19540] <= 8'h00;
            reg_file[19541] <= 8'h00;
            reg_file[19542] <= 8'h00;
            reg_file[19543] <= 8'h00;
            reg_file[19544] <= 8'h00;
            reg_file[19545] <= 8'h00;
            reg_file[19546] <= 8'h00;
            reg_file[19547] <= 8'h00;
            reg_file[19548] <= 8'h00;
            reg_file[19549] <= 8'h00;
            reg_file[19550] <= 8'h00;
            reg_file[19551] <= 8'h00;
            reg_file[19552] <= 8'h00;
            reg_file[19553] <= 8'h00;
            reg_file[19554] <= 8'h00;
            reg_file[19555] <= 8'h00;
            reg_file[19556] <= 8'h00;
            reg_file[19557] <= 8'h00;
            reg_file[19558] <= 8'h00;
            reg_file[19559] <= 8'h00;
            reg_file[19560] <= 8'h00;
            reg_file[19561] <= 8'h00;
            reg_file[19562] <= 8'h00;
            reg_file[19563] <= 8'h00;
            reg_file[19564] <= 8'h00;
            reg_file[19565] <= 8'h00;
            reg_file[19566] <= 8'h00;
            reg_file[19567] <= 8'h00;
            reg_file[19568] <= 8'h00;
            reg_file[19569] <= 8'h00;
            reg_file[19570] <= 8'h00;
            reg_file[19571] <= 8'h00;
            reg_file[19572] <= 8'h00;
            reg_file[19573] <= 8'h00;
            reg_file[19574] <= 8'h00;
            reg_file[19575] <= 8'h00;
            reg_file[19576] <= 8'h00;
            reg_file[19577] <= 8'h00;
            reg_file[19578] <= 8'h00;
            reg_file[19579] <= 8'h00;
            reg_file[19580] <= 8'h00;
            reg_file[19581] <= 8'h00;
            reg_file[19582] <= 8'h00;
            reg_file[19583] <= 8'h00;
            reg_file[19584] <= 8'h00;
            reg_file[19585] <= 8'h00;
            reg_file[19586] <= 8'h00;
            reg_file[19587] <= 8'h00;
            reg_file[19588] <= 8'h00;
            reg_file[19589] <= 8'h00;
            reg_file[19590] <= 8'h00;
            reg_file[19591] <= 8'h00;
            reg_file[19592] <= 8'h00;
            reg_file[19593] <= 8'h00;
            reg_file[19594] <= 8'h00;
            reg_file[19595] <= 8'h00;
            reg_file[19596] <= 8'h00;
            reg_file[19597] <= 8'h00;
            reg_file[19598] <= 8'h00;
            reg_file[19599] <= 8'h00;
            reg_file[19600] <= 8'h00;
            reg_file[19601] <= 8'h00;
            reg_file[19602] <= 8'h00;
            reg_file[19603] <= 8'h00;
            reg_file[19604] <= 8'h00;
            reg_file[19605] <= 8'h00;
            reg_file[19606] <= 8'h00;
            reg_file[19607] <= 8'h00;
            reg_file[19608] <= 8'h00;
            reg_file[19609] <= 8'h00;
            reg_file[19610] <= 8'h00;
            reg_file[19611] <= 8'h00;
            reg_file[19612] <= 8'h00;
            reg_file[19613] <= 8'h00;
            reg_file[19614] <= 8'h00;
            reg_file[19615] <= 8'h00;
            reg_file[19616] <= 8'h00;
            reg_file[19617] <= 8'h00;
            reg_file[19618] <= 8'h00;
            reg_file[19619] <= 8'h00;
            reg_file[19620] <= 8'h00;
            reg_file[19621] <= 8'h00;
            reg_file[19622] <= 8'h00;
            reg_file[19623] <= 8'h00;
            reg_file[19624] <= 8'h00;
            reg_file[19625] <= 8'h00;
            reg_file[19626] <= 8'h00;
            reg_file[19627] <= 8'h00;
            reg_file[19628] <= 8'h00;
            reg_file[19629] <= 8'h00;
            reg_file[19630] <= 8'h00;
            reg_file[19631] <= 8'h00;
            reg_file[19632] <= 8'h00;
            reg_file[19633] <= 8'h00;
            reg_file[19634] <= 8'h00;
            reg_file[19635] <= 8'h00;
            reg_file[19636] <= 8'h00;
            reg_file[19637] <= 8'h00;
            reg_file[19638] <= 8'h00;
            reg_file[19639] <= 8'h00;
            reg_file[19640] <= 8'h00;
            reg_file[19641] <= 8'h00;
            reg_file[19642] <= 8'h00;
            reg_file[19643] <= 8'h00;
            reg_file[19644] <= 8'h00;
            reg_file[19645] <= 8'h00;
            reg_file[19646] <= 8'h00;
            reg_file[19647] <= 8'h00;
            reg_file[19648] <= 8'h00;
            reg_file[19649] <= 8'h00;
            reg_file[19650] <= 8'h00;
            reg_file[19651] <= 8'h00;
            reg_file[19652] <= 8'h00;
            reg_file[19653] <= 8'h00;
            reg_file[19654] <= 8'h00;
            reg_file[19655] <= 8'h00;
            reg_file[19656] <= 8'h00;
            reg_file[19657] <= 8'h00;
            reg_file[19658] <= 8'h00;
            reg_file[19659] <= 8'h00;
            reg_file[19660] <= 8'h00;
            reg_file[19661] <= 8'h00;
            reg_file[19662] <= 8'h00;
            reg_file[19663] <= 8'h00;
            reg_file[19664] <= 8'h00;
            reg_file[19665] <= 8'h00;
            reg_file[19666] <= 8'h00;
            reg_file[19667] <= 8'h00;
            reg_file[19668] <= 8'h00;
            reg_file[19669] <= 8'h00;
            reg_file[19670] <= 8'h00;
            reg_file[19671] <= 8'h00;
            reg_file[19672] <= 8'h00;
            reg_file[19673] <= 8'h00;
            reg_file[19674] <= 8'h00;
            reg_file[19675] <= 8'h00;
            reg_file[19676] <= 8'h00;
            reg_file[19677] <= 8'h00;
            reg_file[19678] <= 8'h00;
            reg_file[19679] <= 8'h00;
            reg_file[19680] <= 8'h00;
            reg_file[19681] <= 8'h00;
            reg_file[19682] <= 8'h00;
            reg_file[19683] <= 8'h00;
            reg_file[19684] <= 8'h00;
            reg_file[19685] <= 8'h00;
            reg_file[19686] <= 8'h00;
            reg_file[19687] <= 8'h00;
            reg_file[19688] <= 8'h00;
            reg_file[19689] <= 8'h00;
            reg_file[19690] <= 8'h00;
            reg_file[19691] <= 8'h00;
            reg_file[19692] <= 8'h00;
            reg_file[19693] <= 8'h00;
            reg_file[19694] <= 8'h00;
            reg_file[19695] <= 8'h00;
            reg_file[19696] <= 8'hC8;
            reg_file[19697] <= 8'h48;
            reg_file[19698] <= 8'h00;
            reg_file[19699] <= 8'h80;
            reg_file[19700] <= 8'h00;
            reg_file[19701] <= 8'h00;
            reg_file[19702] <= 8'h00;
            reg_file[19703] <= 8'h00;
            reg_file[19704] <= 8'h7C;
            reg_file[19705] <= 8'h0F;
            reg_file[19706] <= 8'h97;
            reg_file[19707] <= 8'h1C;
            reg_file[19708] <= 8'h67;
            reg_file[19709] <= 8'hCB;
            reg_file[19710] <= 8'hB4;
            reg_file[19711] <= 8'h40;
            reg_file[19712] <= 8'h72;
            reg_file[19713] <= 8'h33;
            reg_file[19714] <= 8'hDC;
            reg_file[19715] <= 8'h80;
            reg_file[19716] <= 8'h1F;
            reg_file[19717] <= 8'hA3;
            reg_file[19718] <= 8'hB0;
            reg_file[19719] <= 8'h40;
            reg_file[19720] <= 8'hC8;
            reg_file[19721] <= 8'h48;
            reg_file[19722] <= 8'h00;
            reg_file[19723] <= 8'h80;
            reg_file[19724] <= 8'h00;
            reg_file[19725] <= 8'h00;
            reg_file[19726] <= 8'h00;
            reg_file[19727] <= 8'h00;
            reg_file[19728] <= 8'h00;
            reg_file[19729] <= 8'h00;
            reg_file[19730] <= 8'h00;
            reg_file[19731] <= 8'h00;
            reg_file[19732] <= 8'h00;
            reg_file[19733] <= 8'h00;
            reg_file[19734] <= 8'h00;
            reg_file[19735] <= 8'h00;
            reg_file[19736] <= 8'h00;
            reg_file[19737] <= 8'h00;
            reg_file[19738] <= 8'h00;
            reg_file[19739] <= 8'h00;
            reg_file[19740] <= 8'h00;
            reg_file[19741] <= 8'h00;
            reg_file[19742] <= 8'h00;
            reg_file[19743] <= 8'h00;
            reg_file[19744] <= 8'h00;
            reg_file[19745] <= 8'h00;
            reg_file[19746] <= 8'h00;
            reg_file[19747] <= 8'h00;
            reg_file[19748] <= 8'h00;
            reg_file[19749] <= 8'h00;
            reg_file[19750] <= 8'h00;
            reg_file[19751] <= 8'h00;
            reg_file[19752] <= 8'h00;
            reg_file[19753] <= 8'h00;
            reg_file[19754] <= 8'h00;
            reg_file[19755] <= 8'h00;
            reg_file[19756] <= 8'h00;
            reg_file[19757] <= 8'h00;
            reg_file[19758] <= 8'h00;
            reg_file[19759] <= 8'h00;
            reg_file[19760] <= 8'h00;
            reg_file[19761] <= 8'h00;
            reg_file[19762] <= 8'h00;
            reg_file[19763] <= 8'h00;
            reg_file[19764] <= 8'h00;
            reg_file[19765] <= 8'h00;
            reg_file[19766] <= 8'h00;
            reg_file[19767] <= 8'h00;
            reg_file[19768] <= 8'h00;
            reg_file[19769] <= 8'h00;
            reg_file[19770] <= 8'h00;
            reg_file[19771] <= 8'h00;
            reg_file[19772] <= 8'h00;
            reg_file[19773] <= 8'h00;
            reg_file[19774] <= 8'h00;
            reg_file[19775] <= 8'h00;
            reg_file[19776] <= 8'h00;
            reg_file[19777] <= 8'h00;
            reg_file[19778] <= 8'h00;
            reg_file[19779] <= 8'h00;
            reg_file[19780] <= 8'h00;
            reg_file[19781] <= 8'h00;
            reg_file[19782] <= 8'h00;
            reg_file[19783] <= 8'h00;
            reg_file[19784] <= 8'h00;
            reg_file[19785] <= 8'h00;
            reg_file[19786] <= 8'h00;
            reg_file[19787] <= 8'h00;
            reg_file[19788] <= 8'h00;
            reg_file[19789] <= 8'h00;
            reg_file[19790] <= 8'h00;
            reg_file[19791] <= 8'h00;
            reg_file[19792] <= 8'h00;
            reg_file[19793] <= 8'h00;
            reg_file[19794] <= 8'h00;
            reg_file[19795] <= 8'h00;
            reg_file[19796] <= 8'h00;
            reg_file[19797] <= 8'h00;
            reg_file[19798] <= 8'h00;
            reg_file[19799] <= 8'h00;
            reg_file[19800] <= 8'h00;
            reg_file[19801] <= 8'h00;
            reg_file[19802] <= 8'h00;
            reg_file[19803] <= 8'h00;
            reg_file[19804] <= 8'h00;
            reg_file[19805] <= 8'h00;
            reg_file[19806] <= 8'h00;
            reg_file[19807] <= 8'h00;
            reg_file[19808] <= 8'h00;
            reg_file[19809] <= 8'h00;
            reg_file[19810] <= 8'h00;
            reg_file[19811] <= 8'h00;
            reg_file[19812] <= 8'h00;
            reg_file[19813] <= 8'h00;
            reg_file[19814] <= 8'h00;
            reg_file[19815] <= 8'h00;
            reg_file[19816] <= 8'h00;
            reg_file[19817] <= 8'h00;
            reg_file[19818] <= 8'h00;
            reg_file[19819] <= 8'h00;
            reg_file[19820] <= 8'h00;
            reg_file[19821] <= 8'h00;
            reg_file[19822] <= 8'h00;
            reg_file[19823] <= 8'h00;
            reg_file[19824] <= 8'h00;
            reg_file[19825] <= 8'h00;
            reg_file[19826] <= 8'h00;
            reg_file[19827] <= 8'h00;
            reg_file[19828] <= 8'h00;
            reg_file[19829] <= 8'h00;
            reg_file[19830] <= 8'h00;
            reg_file[19831] <= 8'h00;
            reg_file[19832] <= 8'h00;
            reg_file[19833] <= 8'h00;
            reg_file[19834] <= 8'h00;
            reg_file[19835] <= 8'h00;
            reg_file[19836] <= 8'h00;
            reg_file[19837] <= 8'h00;
            reg_file[19838] <= 8'h00;
            reg_file[19839] <= 8'h00;
            reg_file[19840] <= 8'h00;
            reg_file[19841] <= 8'h00;
            reg_file[19842] <= 8'h00;
            reg_file[19843] <= 8'h00;
            reg_file[19844] <= 8'h00;
            reg_file[19845] <= 8'h00;
            reg_file[19846] <= 8'h00;
            reg_file[19847] <= 8'h00;
            reg_file[19848] <= 8'h00;
            reg_file[19849] <= 8'h00;
            reg_file[19850] <= 8'h00;
            reg_file[19851] <= 8'h00;
            reg_file[19852] <= 8'h00;
            reg_file[19853] <= 8'h00;
            reg_file[19854] <= 8'h00;
            reg_file[19855] <= 8'h00;
            reg_file[19856] <= 8'h00;
            reg_file[19857] <= 8'h00;
            reg_file[19858] <= 8'h00;
            reg_file[19859] <= 8'h00;
            reg_file[19860] <= 8'h00;
            reg_file[19861] <= 8'h00;
            reg_file[19862] <= 8'h00;
            reg_file[19863] <= 8'h00;
            reg_file[19864] <= 8'h00;
            reg_file[19865] <= 8'h00;
            reg_file[19866] <= 8'h00;
            reg_file[19867] <= 8'h00;
            reg_file[19868] <= 8'h00;
            reg_file[19869] <= 8'h00;
            reg_file[19870] <= 8'h00;
            reg_file[19871] <= 8'h00;
            reg_file[19872] <= 8'h00;
            reg_file[19873] <= 8'h00;
            reg_file[19874] <= 8'h00;
            reg_file[19875] <= 8'h00;
            reg_file[19876] <= 8'h00;
            reg_file[19877] <= 8'h00;
            reg_file[19878] <= 8'h00;
            reg_file[19879] <= 8'h00;
            reg_file[19880] <= 8'h00;
            reg_file[19881] <= 8'h00;
            reg_file[19882] <= 8'h00;
            reg_file[19883] <= 8'h00;
            reg_file[19884] <= 8'h00;
            reg_file[19885] <= 8'h00;
            reg_file[19886] <= 8'h00;
            reg_file[19887] <= 8'h00;
            reg_file[19888] <= 8'h00;
            reg_file[19889] <= 8'h00;
            reg_file[19890] <= 8'h00;
            reg_file[19891] <= 8'h00;
            reg_file[19892] <= 8'h00;
            reg_file[19893] <= 8'h00;
            reg_file[19894] <= 8'h00;
            reg_file[19895] <= 8'h00;
            reg_file[19896] <= 8'h00;
            reg_file[19897] <= 8'h00;
            reg_file[19898] <= 8'h00;
            reg_file[19899] <= 8'h00;
            reg_file[19900] <= 8'h00;
            reg_file[19901] <= 8'h00;
            reg_file[19902] <= 8'h00;
            reg_file[19903] <= 8'h00;
            reg_file[19904] <= 8'h00;
            reg_file[19905] <= 8'h00;
            reg_file[19906] <= 8'h00;
            reg_file[19907] <= 8'h00;
            reg_file[19908] <= 8'h00;
            reg_file[19909] <= 8'h00;
            reg_file[19910] <= 8'h00;
            reg_file[19911] <= 8'h00;
            reg_file[19912] <= 8'h00;
            reg_file[19913] <= 8'h00;
            reg_file[19914] <= 8'h00;
            reg_file[19915] <= 8'h00;
            reg_file[19916] <= 8'h00;
            reg_file[19917] <= 8'h00;
            reg_file[19918] <= 8'h00;
            reg_file[19919] <= 8'h00;
            reg_file[19920] <= 8'h00;
            reg_file[19921] <= 8'h00;
            reg_file[19922] <= 8'h00;
            reg_file[19923] <= 8'h00;
            reg_file[19924] <= 8'h00;
            reg_file[19925] <= 8'h00;
            reg_file[19926] <= 8'h00;
            reg_file[19927] <= 8'h00;
            reg_file[19928] <= 8'h00;
            reg_file[19929] <= 8'h00;
            reg_file[19930] <= 8'h00;
            reg_file[19931] <= 8'h00;
            reg_file[19932] <= 8'h00;
            reg_file[19933] <= 8'h00;
            reg_file[19934] <= 8'h00;
            reg_file[19935] <= 8'h00;
            reg_file[19936] <= 8'h00;
            reg_file[19937] <= 8'h00;
            reg_file[19938] <= 8'h00;
            reg_file[19939] <= 8'h00;
            reg_file[19940] <= 8'h00;
            reg_file[19941] <= 8'h00;
            reg_file[19942] <= 8'h00;
            reg_file[19943] <= 8'h00;
            reg_file[19944] <= 8'h00;
            reg_file[19945] <= 8'h00;
            reg_file[19946] <= 8'h00;
            reg_file[19947] <= 8'h00;
            reg_file[19948] <= 8'h00;
            reg_file[19949] <= 8'h00;
            reg_file[19950] <= 8'h00;
            reg_file[19951] <= 8'h00;
            reg_file[19952] <= 8'h00;
            reg_file[19953] <= 8'h00;
            reg_file[19954] <= 8'h00;
            reg_file[19955] <= 8'h00;
            reg_file[19956] <= 8'h00;
            reg_file[19957] <= 8'h00;
            reg_file[19958] <= 8'h00;
            reg_file[19959] <= 8'h00;
            reg_file[19960] <= 8'h00;
            reg_file[19961] <= 8'h00;
            reg_file[19962] <= 8'h00;
            reg_file[19963] <= 8'h00;
            reg_file[19964] <= 8'h00;
            reg_file[19965] <= 8'h00;
            reg_file[19966] <= 8'h00;
            reg_file[19967] <= 8'h00;
            reg_file[19968] <= 8'h00;
            reg_file[19969] <= 8'h00;
            reg_file[19970] <= 8'h00;
            reg_file[19971] <= 8'h00;
            reg_file[19972] <= 8'h00;
            reg_file[19973] <= 8'h00;
            reg_file[19974] <= 8'h00;
            reg_file[19975] <= 8'h00;
            reg_file[19976] <= 8'h00;
            reg_file[19977] <= 8'h00;
            reg_file[19978] <= 8'h00;
            reg_file[19979] <= 8'h00;
            reg_file[19980] <= 8'h00;
            reg_file[19981] <= 8'h00;
            reg_file[19982] <= 8'h00;
            reg_file[19983] <= 8'h00;
            reg_file[19984] <= 8'h00;
            reg_file[19985] <= 8'h00;
            reg_file[19986] <= 8'h00;
            reg_file[19987] <= 8'h00;
            reg_file[19988] <= 8'h00;
            reg_file[19989] <= 8'h00;
            reg_file[19990] <= 8'h00;
            reg_file[19991] <= 8'h00;
            reg_file[19992] <= 8'h00;
            reg_file[19993] <= 8'h00;
            reg_file[19994] <= 8'h00;
            reg_file[19995] <= 8'h00;
            reg_file[19996] <= 8'h00;
            reg_file[19997] <= 8'h00;
            reg_file[19998] <= 8'h00;
            reg_file[19999] <= 8'h00;
            reg_file[20000] <= 8'h00;
            reg_file[20001] <= 8'h00;
            reg_file[20002] <= 8'h00;
            reg_file[20003] <= 8'h00;
            reg_file[20004] <= 8'h00;
            reg_file[20005] <= 8'h00;
            reg_file[20006] <= 8'h00;
            reg_file[20007] <= 8'h00;
            reg_file[20008] <= 8'h00;
            reg_file[20009] <= 8'h00;
            reg_file[20010] <= 8'h00;
            reg_file[20011] <= 8'h00;
            reg_file[20012] <= 8'h00;
            reg_file[20013] <= 8'h00;
            reg_file[20014] <= 8'h00;
            reg_file[20015] <= 8'h00;
            reg_file[20016] <= 8'h00;
            reg_file[20017] <= 8'h00;
            reg_file[20018] <= 8'h00;
            reg_file[20019] <= 8'h00;
            reg_file[20020] <= 8'h00;
            reg_file[20021] <= 8'h00;
            reg_file[20022] <= 8'h00;
            reg_file[20023] <= 8'h00;
            reg_file[20024] <= 8'h00;
            reg_file[20025] <= 8'h00;
            reg_file[20026] <= 8'h00;
            reg_file[20027] <= 8'h00;
            reg_file[20028] <= 8'h00;
            reg_file[20029] <= 8'h00;
            reg_file[20030] <= 8'h00;
            reg_file[20031] <= 8'h00;
            reg_file[20032] <= 8'h00;
            reg_file[20033] <= 8'h00;
            reg_file[20034] <= 8'h00;
            reg_file[20035] <= 8'h00;
            reg_file[20036] <= 8'h00;
            reg_file[20037] <= 8'h00;
            reg_file[20038] <= 8'h00;
            reg_file[20039] <= 8'h00;
            reg_file[20040] <= 8'h00;
            reg_file[20041] <= 8'h00;
            reg_file[20042] <= 8'h00;
            reg_file[20043] <= 8'h00;
            reg_file[20044] <= 8'h00;
            reg_file[20045] <= 8'h00;
            reg_file[20046] <= 8'h00;
            reg_file[20047] <= 8'h00;
            reg_file[20048] <= 8'h00;
            reg_file[20049] <= 8'h00;
            reg_file[20050] <= 8'h00;
            reg_file[20051] <= 8'h00;
            reg_file[20052] <= 8'h00;
            reg_file[20053] <= 8'h00;
            reg_file[20054] <= 8'h00;
            reg_file[20055] <= 8'h00;
            reg_file[20056] <= 8'h00;
            reg_file[20057] <= 8'h00;
            reg_file[20058] <= 8'h00;
            reg_file[20059] <= 8'h00;
            reg_file[20060] <= 8'h00;
            reg_file[20061] <= 8'h00;
            reg_file[20062] <= 8'h00;
            reg_file[20063] <= 8'h00;
            reg_file[20064] <= 8'h00;
            reg_file[20065] <= 8'h00;
            reg_file[20066] <= 8'h00;
            reg_file[20067] <= 8'h00;
            reg_file[20068] <= 8'h00;
            reg_file[20069] <= 8'h00;
            reg_file[20070] <= 8'h00;
            reg_file[20071] <= 8'h00;
            reg_file[20072] <= 8'h00;
            reg_file[20073] <= 8'h00;
            reg_file[20074] <= 8'h00;
            reg_file[20075] <= 8'h00;
            reg_file[20076] <= 8'h00;
            reg_file[20077] <= 8'h00;
            reg_file[20078] <= 8'h00;
            reg_file[20079] <= 8'h00;
            reg_file[20080] <= 8'h00;
            reg_file[20081] <= 8'h00;
            reg_file[20082] <= 8'h00;
            reg_file[20083] <= 8'h00;
            reg_file[20084] <= 8'h00;
            reg_file[20085] <= 8'h00;
            reg_file[20086] <= 8'h00;
            reg_file[20087] <= 8'h00;
            reg_file[20088] <= 8'h00;
            reg_file[20089] <= 8'h00;
            reg_file[20090] <= 8'h00;
            reg_file[20091] <= 8'h00;
            reg_file[20092] <= 8'h00;
            reg_file[20093] <= 8'h00;
            reg_file[20094] <= 8'h00;
            reg_file[20095] <= 8'h00;
            reg_file[20096] <= 8'h00;
            reg_file[20097] <= 8'h00;
            reg_file[20098] <= 8'h00;
            reg_file[20099] <= 8'h00;
            reg_file[20100] <= 8'h00;
            reg_file[20101] <= 8'h00;
            reg_file[20102] <= 8'h00;
            reg_file[20103] <= 8'h00;
            reg_file[20104] <= 8'h00;
            reg_file[20105] <= 8'h00;
            reg_file[20106] <= 8'h00;
            reg_file[20107] <= 8'h00;
            reg_file[20108] <= 8'h00;
            reg_file[20109] <= 8'h00;
            reg_file[20110] <= 8'h00;
            reg_file[20111] <= 8'h00;
            reg_file[20112] <= 8'h00;
            reg_file[20113] <= 8'h00;
            reg_file[20114] <= 8'h00;
            reg_file[20115] <= 8'h00;
            reg_file[20116] <= 8'h00;
            reg_file[20117] <= 8'h00;
            reg_file[20118] <= 8'h00;
            reg_file[20119] <= 8'h00;
            reg_file[20120] <= 8'h00;
            reg_file[20121] <= 8'h00;
            reg_file[20122] <= 8'h00;
            reg_file[20123] <= 8'h00;
            reg_file[20124] <= 8'h00;
            reg_file[20125] <= 8'h00;
            reg_file[20126] <= 8'h00;
            reg_file[20127] <= 8'h00;
            reg_file[20128] <= 8'h00;
            reg_file[20129] <= 8'h00;
            reg_file[20130] <= 8'h00;
            reg_file[20131] <= 8'h00;
            reg_file[20132] <= 8'h00;
            reg_file[20133] <= 8'h00;
            reg_file[20134] <= 8'h00;
            reg_file[20135] <= 8'h00;
            reg_file[20136] <= 8'h00;
            reg_file[20137] <= 8'h00;
            reg_file[20138] <= 8'h00;
            reg_file[20139] <= 8'h00;
            reg_file[20140] <= 8'h00;
            reg_file[20141] <= 8'h00;
            reg_file[20142] <= 8'h00;
            reg_file[20143] <= 8'h00;
            reg_file[20144] <= 8'h00;
            reg_file[20145] <= 8'h00;
            reg_file[20146] <= 8'h00;
            reg_file[20147] <= 8'h00;
            reg_file[20148] <= 8'h00;
            reg_file[20149] <= 8'h00;
            reg_file[20150] <= 8'h00;
            reg_file[20151] <= 8'h00;
            reg_file[20152] <= 8'h00;
            reg_file[20153] <= 8'h00;
            reg_file[20154] <= 8'h00;
            reg_file[20155] <= 8'h00;
            reg_file[20156] <= 8'h00;
            reg_file[20157] <= 8'h00;
            reg_file[20158] <= 8'h00;
            reg_file[20159] <= 8'h00;
            reg_file[20160] <= 8'h00;
            reg_file[20161] <= 8'h00;
            reg_file[20162] <= 8'h00;
            reg_file[20163] <= 8'h00;
            reg_file[20164] <= 8'h00;
            reg_file[20165] <= 8'h00;
            reg_file[20166] <= 8'h00;
            reg_file[20167] <= 8'h00;
            reg_file[20168] <= 8'h00;
            reg_file[20169] <= 8'h00;
            reg_file[20170] <= 8'h00;
            reg_file[20171] <= 8'h00;
            reg_file[20172] <= 8'h00;
            reg_file[20173] <= 8'h00;
            reg_file[20174] <= 8'h00;
            reg_file[20175] <= 8'h00;
            reg_file[20176] <= 8'h00;
            reg_file[20177] <= 8'h00;
            reg_file[20178] <= 8'h00;
            reg_file[20179] <= 8'h00;
            reg_file[20180] <= 8'h00;
            reg_file[20181] <= 8'h00;
            reg_file[20182] <= 8'h00;
            reg_file[20183] <= 8'h00;
            reg_file[20184] <= 8'h00;
            reg_file[20185] <= 8'h00;
            reg_file[20186] <= 8'h00;
            reg_file[20187] <= 8'h00;
            reg_file[20188] <= 8'h00;
            reg_file[20189] <= 8'h00;
            reg_file[20190] <= 8'h00;
            reg_file[20191] <= 8'h00;
            reg_file[20192] <= 8'h00;
            reg_file[20193] <= 8'h00;
            reg_file[20194] <= 8'h00;
            reg_file[20195] <= 8'h00;
            reg_file[20196] <= 8'h00;
            reg_file[20197] <= 8'h00;
            reg_file[20198] <= 8'h00;
            reg_file[20199] <= 8'h00;
            reg_file[20200] <= 8'h00;
            reg_file[20201] <= 8'h00;
            reg_file[20202] <= 8'h00;
            reg_file[20203] <= 8'h00;
            reg_file[20204] <= 8'h00;
            reg_file[20205] <= 8'h00;
            reg_file[20206] <= 8'h00;
            reg_file[20207] <= 8'h00;
            reg_file[20208] <= 8'h00;
            reg_file[20209] <= 8'h00;
            reg_file[20210] <= 8'h00;
            reg_file[20211] <= 8'h00;
            reg_file[20212] <= 8'h00;
            reg_file[20213] <= 8'h00;
            reg_file[20214] <= 8'h00;
            reg_file[20215] <= 8'h00;
            reg_file[20216] <= 8'h00;
            reg_file[20217] <= 8'h00;
            reg_file[20218] <= 8'h00;
            reg_file[20219] <= 8'h00;
            reg_file[20220] <= 8'h00;
            reg_file[20221] <= 8'h00;
            reg_file[20222] <= 8'h00;
            reg_file[20223] <= 8'h00;
            reg_file[20224] <= 8'h00;
            reg_file[20225] <= 8'h00;
            reg_file[20226] <= 8'h00;
            reg_file[20227] <= 8'h00;
            reg_file[20228] <= 8'h00;
            reg_file[20229] <= 8'h00;
            reg_file[20230] <= 8'h00;
            reg_file[20231] <= 8'h00;
            reg_file[20232] <= 8'h00;
            reg_file[20233] <= 8'h00;
            reg_file[20234] <= 8'h00;
            reg_file[20235] <= 8'h00;
            reg_file[20236] <= 8'h00;
            reg_file[20237] <= 8'h00;
            reg_file[20238] <= 8'h00;
            reg_file[20239] <= 8'h00;
            reg_file[20240] <= 8'h00;
            reg_file[20241] <= 8'h00;
            reg_file[20242] <= 8'h00;
            reg_file[20243] <= 8'h00;
            reg_file[20244] <= 8'h00;
            reg_file[20245] <= 8'h00;
            reg_file[20246] <= 8'h00;
            reg_file[20247] <= 8'h00;
            reg_file[20248] <= 8'h00;
            reg_file[20249] <= 8'h00;
            reg_file[20250] <= 8'h00;
            reg_file[20251] <= 8'h00;
            reg_file[20252] <= 8'h00;
            reg_file[20253] <= 8'h00;
            reg_file[20254] <= 8'h00;
            reg_file[20255] <= 8'h00;
            reg_file[20256] <= 8'h00;
            reg_file[20257] <= 8'h00;
            reg_file[20258] <= 8'h00;
            reg_file[20259] <= 8'h00;
            reg_file[20260] <= 8'h00;
            reg_file[20261] <= 8'h00;
            reg_file[20262] <= 8'h00;
            reg_file[20263] <= 8'h00;
            reg_file[20264] <= 8'h00;
            reg_file[20265] <= 8'h00;
            reg_file[20266] <= 8'h00;
            reg_file[20267] <= 8'h00;
            reg_file[20268] <= 8'h00;
            reg_file[20269] <= 8'h00;
            reg_file[20270] <= 8'h00;
            reg_file[20271] <= 8'h00;
            reg_file[20272] <= 8'h00;
            reg_file[20273] <= 8'h00;
            reg_file[20274] <= 8'h00;
            reg_file[20275] <= 8'h00;
            reg_file[20276] <= 8'h00;
            reg_file[20277] <= 8'h00;
            reg_file[20278] <= 8'h00;
            reg_file[20279] <= 8'h00;
            reg_file[20280] <= 8'h00;
            reg_file[20281] <= 8'h00;
            reg_file[20282] <= 8'h00;
            reg_file[20283] <= 8'h00;
            reg_file[20284] <= 8'h00;
            reg_file[20285] <= 8'h00;
            reg_file[20286] <= 8'h00;
            reg_file[20287] <= 8'h00;
            reg_file[20288] <= 8'h00;
            reg_file[20289] <= 8'h00;
            reg_file[20290] <= 8'h00;
            reg_file[20291] <= 8'h00;
            reg_file[20292] <= 8'h00;
            reg_file[20293] <= 8'h00;
            reg_file[20294] <= 8'h00;
            reg_file[20295] <= 8'h00;
            reg_file[20296] <= 8'h00;
            reg_file[20297] <= 8'h00;
            reg_file[20298] <= 8'h00;
            reg_file[20299] <= 8'h00;
            reg_file[20300] <= 8'h00;
            reg_file[20301] <= 8'h00;
            reg_file[20302] <= 8'h00;
            reg_file[20303] <= 8'h00;
            reg_file[20304] <= 8'h00;
            reg_file[20305] <= 8'h00;
            reg_file[20306] <= 8'h00;
            reg_file[20307] <= 8'h00;
            reg_file[20308] <= 8'h00;
            reg_file[20309] <= 8'h00;
            reg_file[20310] <= 8'h00;
            reg_file[20311] <= 8'h00;
            reg_file[20312] <= 8'h00;
            reg_file[20313] <= 8'h00;
            reg_file[20314] <= 8'h00;
            reg_file[20315] <= 8'h00;
            reg_file[20316] <= 8'h00;
            reg_file[20317] <= 8'h00;
            reg_file[20318] <= 8'h00;
            reg_file[20319] <= 8'h00;
            reg_file[20320] <= 8'h00;
            reg_file[20321] <= 8'h00;
            reg_file[20322] <= 8'h00;
            reg_file[20323] <= 8'h00;
            reg_file[20324] <= 8'h00;
            reg_file[20325] <= 8'h00;
            reg_file[20326] <= 8'h00;
            reg_file[20327] <= 8'h00;
            reg_file[20328] <= 8'h00;
            reg_file[20329] <= 8'h00;
            reg_file[20330] <= 8'h00;
            reg_file[20331] <= 8'h00;
            reg_file[20332] <= 8'h00;
            reg_file[20333] <= 8'h00;
            reg_file[20334] <= 8'h00;
            reg_file[20335] <= 8'h00;
            reg_file[20336] <= 8'h00;
            reg_file[20337] <= 8'h00;
            reg_file[20338] <= 8'h00;
            reg_file[20339] <= 8'h00;
            reg_file[20340] <= 8'h00;
            reg_file[20341] <= 8'h00;
            reg_file[20342] <= 8'h00;
            reg_file[20343] <= 8'h00;
            reg_file[20344] <= 8'h00;
            reg_file[20345] <= 8'h00;
            reg_file[20346] <= 8'h00;
            reg_file[20347] <= 8'h00;
            reg_file[20348] <= 8'h00;
            reg_file[20349] <= 8'h00;
            reg_file[20350] <= 8'h00;
            reg_file[20351] <= 8'h00;
            reg_file[20352] <= 8'h00;
            reg_file[20353] <= 8'h00;
            reg_file[20354] <= 8'h00;
            reg_file[20355] <= 8'h00;
            reg_file[20356] <= 8'h00;
            reg_file[20357] <= 8'h00;
            reg_file[20358] <= 8'h00;
            reg_file[20359] <= 8'h00;
            reg_file[20360] <= 8'h00;
            reg_file[20361] <= 8'h00;
            reg_file[20362] <= 8'h00;
            reg_file[20363] <= 8'h00;
            reg_file[20364] <= 8'h00;
            reg_file[20365] <= 8'h00;
            reg_file[20366] <= 8'h00;
            reg_file[20367] <= 8'h00;
            reg_file[20368] <= 8'h00;
            reg_file[20369] <= 8'h00;
            reg_file[20370] <= 8'h00;
            reg_file[20371] <= 8'h00;
            reg_file[20372] <= 8'h00;
            reg_file[20373] <= 8'h00;
            reg_file[20374] <= 8'h00;
            reg_file[20375] <= 8'h00;
            reg_file[20376] <= 8'h00;
            reg_file[20377] <= 8'h00;
            reg_file[20378] <= 8'h00;
            reg_file[20379] <= 8'h00;
            reg_file[20380] <= 8'h00;
            reg_file[20381] <= 8'h00;
            reg_file[20382] <= 8'h00;
            reg_file[20383] <= 8'h00;
            reg_file[20384] <= 8'h00;
            reg_file[20385] <= 8'h00;
            reg_file[20386] <= 8'h00;
            reg_file[20387] <= 8'h00;
            reg_file[20388] <= 8'h00;
            reg_file[20389] <= 8'h00;
            reg_file[20390] <= 8'h00;
            reg_file[20391] <= 8'h00;
            reg_file[20392] <= 8'h00;
            reg_file[20393] <= 8'h00;
            reg_file[20394] <= 8'h00;
            reg_file[20395] <= 8'h00;
            reg_file[20396] <= 8'h00;
            reg_file[20397] <= 8'h00;
            reg_file[20398] <= 8'h00;
            reg_file[20399] <= 8'h00;
            reg_file[20400] <= 8'h00;
            reg_file[20401] <= 8'h00;
            reg_file[20402] <= 8'h00;
            reg_file[20403] <= 8'h00;
            reg_file[20404] <= 8'h00;
            reg_file[20405] <= 8'h00;
            reg_file[20406] <= 8'h00;
            reg_file[20407] <= 8'h00;
            reg_file[20408] <= 8'h00;
            reg_file[20409] <= 8'h00;
            reg_file[20410] <= 8'h00;
            reg_file[20411] <= 8'h00;
            reg_file[20412] <= 8'h00;
            reg_file[20413] <= 8'h00;
            reg_file[20414] <= 8'h00;
            reg_file[20415] <= 8'h00;
            reg_file[20416] <= 8'h00;
            reg_file[20417] <= 8'h00;
            reg_file[20418] <= 8'h00;
            reg_file[20419] <= 8'h00;
            reg_file[20420] <= 8'h00;
            reg_file[20421] <= 8'h00;
            reg_file[20422] <= 8'h00;
            reg_file[20423] <= 8'h00;
            reg_file[20424] <= 8'h00;
            reg_file[20425] <= 8'h00;
            reg_file[20426] <= 8'h00;
            reg_file[20427] <= 8'h00;
            reg_file[20428] <= 8'h00;
            reg_file[20429] <= 8'h00;
            reg_file[20430] <= 8'h00;
            reg_file[20431] <= 8'h00;
            reg_file[20432] <= 8'h00;
            reg_file[20433] <= 8'h00;
            reg_file[20434] <= 8'h00;
            reg_file[20435] <= 8'h00;
            reg_file[20436] <= 8'h00;
            reg_file[20437] <= 8'h00;
            reg_file[20438] <= 8'h00;
            reg_file[20439] <= 8'h00;
            reg_file[20440] <= 8'h00;
            reg_file[20441] <= 8'h00;
            reg_file[20442] <= 8'h00;
            reg_file[20443] <= 8'h00;
            reg_file[20444] <= 8'h00;
            reg_file[20445] <= 8'h00;
            reg_file[20446] <= 8'h00;
            reg_file[20447] <= 8'h00;
            reg_file[20448] <= 8'h00;
            reg_file[20449] <= 8'h00;
            reg_file[20450] <= 8'h00;
            reg_file[20451] <= 8'h00;
            reg_file[20452] <= 8'h00;
            reg_file[20453] <= 8'h00;
            reg_file[20454] <= 8'h00;
            reg_file[20455] <= 8'h00;
            reg_file[20456] <= 8'h00;
            reg_file[20457] <= 8'h00;
            reg_file[20458] <= 8'h00;
            reg_file[20459] <= 8'h00;
            reg_file[20460] <= 8'h00;
            reg_file[20461] <= 8'h00;
            reg_file[20462] <= 8'h00;
            reg_file[20463] <= 8'h00;
            reg_file[20464] <= 8'h00;
            reg_file[20465] <= 8'h00;
            reg_file[20466] <= 8'h00;
            reg_file[20467] <= 8'h00;
            reg_file[20468] <= 8'h00;
            reg_file[20469] <= 8'h00;
            reg_file[20470] <= 8'h00;
            reg_file[20471] <= 8'h00;
            reg_file[20472] <= 8'h00;
            reg_file[20473] <= 8'h00;
            reg_file[20474] <= 8'h00;
            reg_file[20475] <= 8'h00;
            reg_file[20476] <= 8'h00;
            reg_file[20477] <= 8'h00;
            reg_file[20478] <= 8'h00;
            reg_file[20479] <= 8'h00;
            reg_file[20480] <= 8'h00;
            reg_file[20481] <= 8'h00;
            reg_file[20482] <= 8'h00;
            reg_file[20483] <= 8'h00;
            reg_file[20484] <= 8'h00;
            reg_file[20485] <= 8'h00;
            reg_file[20486] <= 8'h00;
            reg_file[20487] <= 8'h00;
            reg_file[20488] <= 8'h00;
            reg_file[20489] <= 8'h00;
            reg_file[20490] <= 8'h00;
            reg_file[20491] <= 8'h00;
            reg_file[20492] <= 8'h00;
            reg_file[20493] <= 8'h00;
            reg_file[20494] <= 8'h00;
            reg_file[20495] <= 8'h00;
            reg_file[20496] <= 8'h00;
            reg_file[20497] <= 8'h00;
            reg_file[20498] <= 8'h00;
            reg_file[20499] <= 8'h00;
            reg_file[20500] <= 8'h00;
            reg_file[20501] <= 8'h00;
            reg_file[20502] <= 8'h00;
            reg_file[20503] <= 8'h00;
            reg_file[20504] <= 8'h00;
            reg_file[20505] <= 8'h00;
            reg_file[20506] <= 8'h00;
            reg_file[20507] <= 8'h00;
            reg_file[20508] <= 8'h00;
            reg_file[20509] <= 8'h00;
            reg_file[20510] <= 8'h00;
            reg_file[20511] <= 8'h00;
            reg_file[20512] <= 8'h00;
            reg_file[20513] <= 8'h00;
            reg_file[20514] <= 8'h00;
            reg_file[20515] <= 8'h00;
            reg_file[20516] <= 8'h00;
            reg_file[20517] <= 8'h00;
            reg_file[20518] <= 8'h00;
            reg_file[20519] <= 8'h00;
            reg_file[20520] <= 8'h00;
            reg_file[20521] <= 8'h00;
            reg_file[20522] <= 8'h00;
            reg_file[20523] <= 8'h00;
            reg_file[20524] <= 8'h00;
            reg_file[20525] <= 8'h00;
            reg_file[20526] <= 8'h00;
            reg_file[20527] <= 8'h00;
            reg_file[20528] <= 8'h00;
            reg_file[20529] <= 8'h00;
            reg_file[20530] <= 8'h00;
            reg_file[20531] <= 8'h00;
            reg_file[20532] <= 8'h00;
            reg_file[20533] <= 8'h00;
            reg_file[20534] <= 8'h00;
            reg_file[20535] <= 8'h00;
            reg_file[20536] <= 8'h00;
            reg_file[20537] <= 8'h00;
            reg_file[20538] <= 8'h00;
            reg_file[20539] <= 8'h00;
            reg_file[20540] <= 8'h00;
            reg_file[20541] <= 8'h00;
            reg_file[20542] <= 8'h00;
            reg_file[20543] <= 8'h00;
            reg_file[20544] <= 8'h00;
            reg_file[20545] <= 8'h00;
            reg_file[20546] <= 8'h00;
            reg_file[20547] <= 8'h00;
            reg_file[20548] <= 8'h00;
            reg_file[20549] <= 8'h00;
            reg_file[20550] <= 8'h00;
            reg_file[20551] <= 8'h00;
            reg_file[20552] <= 8'h00;
            reg_file[20553] <= 8'h00;
            reg_file[20554] <= 8'h00;
            reg_file[20555] <= 8'h00;
            reg_file[20556] <= 8'h00;
            reg_file[20557] <= 8'h00;
            reg_file[20558] <= 8'h00;
            reg_file[20559] <= 8'h00;
            reg_file[20560] <= 8'h00;
            reg_file[20561] <= 8'h00;
            reg_file[20562] <= 8'h00;
            reg_file[20563] <= 8'h00;
            reg_file[20564] <= 8'h00;
            reg_file[20565] <= 8'h00;
            reg_file[20566] <= 8'h00;
            reg_file[20567] <= 8'h00;
            reg_file[20568] <= 8'h00;
            reg_file[20569] <= 8'h00;
            reg_file[20570] <= 8'h00;
            reg_file[20571] <= 8'h00;
            reg_file[20572] <= 8'h00;
            reg_file[20573] <= 8'h00;
            reg_file[20574] <= 8'h00;
            reg_file[20575] <= 8'h00;
            reg_file[20576] <= 8'h00;
            reg_file[20577] <= 8'h00;
            reg_file[20578] <= 8'h00;
            reg_file[20579] <= 8'h00;
            reg_file[20580] <= 8'h00;
            reg_file[20581] <= 8'h00;
            reg_file[20582] <= 8'h00;
            reg_file[20583] <= 8'h00;
            reg_file[20584] <= 8'h00;
            reg_file[20585] <= 8'h00;
            reg_file[20586] <= 8'h00;
            reg_file[20587] <= 8'h00;
            reg_file[20588] <= 8'h00;
            reg_file[20589] <= 8'h00;
            reg_file[20590] <= 8'h00;
            reg_file[20591] <= 8'h00;
            reg_file[20592] <= 8'h00;
            reg_file[20593] <= 8'h00;
            reg_file[20594] <= 8'h00;
            reg_file[20595] <= 8'h00;
            reg_file[20596] <= 8'h00;
            reg_file[20597] <= 8'h00;
            reg_file[20598] <= 8'h00;
            reg_file[20599] <= 8'h00;
            reg_file[20600] <= 8'h00;
            reg_file[20601] <= 8'h00;
            reg_file[20602] <= 8'h00;
            reg_file[20603] <= 8'h00;
            reg_file[20604] <= 8'h00;
            reg_file[20605] <= 8'h00;
            reg_file[20606] <= 8'h00;
            reg_file[20607] <= 8'h00;
            reg_file[20608] <= 8'h00;
            reg_file[20609] <= 8'h00;
            reg_file[20610] <= 8'h00;
            reg_file[20611] <= 8'h00;
            reg_file[20612] <= 8'h00;
            reg_file[20613] <= 8'h00;
            reg_file[20614] <= 8'h00;
            reg_file[20615] <= 8'h00;
            reg_file[20616] <= 8'h00;
            reg_file[20617] <= 8'h00;
            reg_file[20618] <= 8'h00;
            reg_file[20619] <= 8'h00;
            reg_file[20620] <= 8'h00;
            reg_file[20621] <= 8'h00;
            reg_file[20622] <= 8'h00;
            reg_file[20623] <= 8'h00;
            reg_file[20624] <= 8'h00;
            reg_file[20625] <= 8'h00;
            reg_file[20626] <= 8'h00;
            reg_file[20627] <= 8'h00;
            reg_file[20628] <= 8'h00;
            reg_file[20629] <= 8'h00;
            reg_file[20630] <= 8'h00;
            reg_file[20631] <= 8'h00;
            reg_file[20632] <= 8'h00;
            reg_file[20633] <= 8'h00;
            reg_file[20634] <= 8'h00;
            reg_file[20635] <= 8'h00;
            reg_file[20636] <= 8'h00;
            reg_file[20637] <= 8'h00;
            reg_file[20638] <= 8'h00;
            reg_file[20639] <= 8'h00;
            reg_file[20640] <= 8'h00;
            reg_file[20641] <= 8'h00;
            reg_file[20642] <= 8'h00;
            reg_file[20643] <= 8'h00;
            reg_file[20644] <= 8'h00;
            reg_file[20645] <= 8'h00;
            reg_file[20646] <= 8'h00;
            reg_file[20647] <= 8'h00;
            reg_file[20648] <= 8'h00;
            reg_file[20649] <= 8'h00;
            reg_file[20650] <= 8'h00;
            reg_file[20651] <= 8'h00;
            reg_file[20652] <= 8'h00;
            reg_file[20653] <= 8'h00;
            reg_file[20654] <= 8'h00;
            reg_file[20655] <= 8'h00;
            reg_file[20656] <= 8'h00;
            reg_file[20657] <= 8'h00;
            reg_file[20658] <= 8'h00;
            reg_file[20659] <= 8'h00;
            reg_file[20660] <= 8'h00;
            reg_file[20661] <= 8'h00;
            reg_file[20662] <= 8'h00;
            reg_file[20663] <= 8'h00;
            reg_file[20664] <= 8'h00;
            reg_file[20665] <= 8'h00;
            reg_file[20666] <= 8'h00;
            reg_file[20667] <= 8'h00;
            reg_file[20668] <= 8'h00;
            reg_file[20669] <= 8'h00;
            reg_file[20670] <= 8'h00;
            reg_file[20671] <= 8'h00;
            reg_file[20672] <= 8'h00;
            reg_file[20673] <= 8'h00;
            reg_file[20674] <= 8'h00;
            reg_file[20675] <= 8'h00;
            reg_file[20676] <= 8'h00;
            reg_file[20677] <= 8'h00;
            reg_file[20678] <= 8'h00;
            reg_file[20679] <= 8'h00;
            reg_file[20680] <= 8'h00;
            reg_file[20681] <= 8'h00;
            reg_file[20682] <= 8'h00;
            reg_file[20683] <= 8'h00;
            reg_file[20684] <= 8'h00;
            reg_file[20685] <= 8'h00;
            reg_file[20686] <= 8'h00;
            reg_file[20687] <= 8'h00;
            reg_file[20688] <= 8'h00;
            reg_file[20689] <= 8'h00;
            reg_file[20690] <= 8'h00;
            reg_file[20691] <= 8'h00;
            reg_file[20692] <= 8'h00;
            reg_file[20693] <= 8'h00;
            reg_file[20694] <= 8'h00;
            reg_file[20695] <= 8'h00;
            reg_file[20696] <= 8'h00;
            reg_file[20697] <= 8'h00;
            reg_file[20698] <= 8'h00;
            reg_file[20699] <= 8'h00;
            reg_file[20700] <= 8'h00;
            reg_file[20701] <= 8'h00;
            reg_file[20702] <= 8'h00;
            reg_file[20703] <= 8'h00;
            reg_file[20704] <= 8'h00;
            reg_file[20705] <= 8'h00;
            reg_file[20706] <= 8'h00;
            reg_file[20707] <= 8'h00;
            reg_file[20708] <= 8'h00;
            reg_file[20709] <= 8'h00;
            reg_file[20710] <= 8'h00;
            reg_file[20711] <= 8'h00;
            reg_file[20712] <= 8'h00;
            reg_file[20713] <= 8'h00;
            reg_file[20714] <= 8'h00;
            reg_file[20715] <= 8'h00;
            reg_file[20716] <= 8'h00;
            reg_file[20717] <= 8'h00;
            reg_file[20718] <= 8'h00;
            reg_file[20719] <= 8'h00;
            reg_file[20720] <= 8'h00;
            reg_file[20721] <= 8'h00;
            reg_file[20722] <= 8'h00;
            reg_file[20723] <= 8'h00;
            reg_file[20724] <= 8'h00;
            reg_file[20725] <= 8'h00;
            reg_file[20726] <= 8'h00;
            reg_file[20727] <= 8'h00;
            reg_file[20728] <= 8'h00;
            reg_file[20729] <= 8'h00;
            reg_file[20730] <= 8'h00;
            reg_file[20731] <= 8'h00;
            reg_file[20732] <= 8'h00;
            reg_file[20733] <= 8'h00;
            reg_file[20734] <= 8'h00;
            reg_file[20735] <= 8'h00;
            reg_file[20736] <= 8'h00;
            reg_file[20737] <= 8'h00;
            reg_file[20738] <= 8'h00;
            reg_file[20739] <= 8'h00;
            reg_file[20740] <= 8'h00;
            reg_file[20741] <= 8'h00;
            reg_file[20742] <= 8'h00;
            reg_file[20743] <= 8'h00;
            reg_file[20744] <= 8'h00;
            reg_file[20745] <= 8'h00;
            reg_file[20746] <= 8'h00;
            reg_file[20747] <= 8'h00;
            reg_file[20748] <= 8'h00;
            reg_file[20749] <= 8'h00;
            reg_file[20750] <= 8'h00;
            reg_file[20751] <= 8'h00;
            reg_file[20752] <= 8'h00;
            reg_file[20753] <= 8'h00;
            reg_file[20754] <= 8'h00;
            reg_file[20755] <= 8'h00;
            reg_file[20756] <= 8'h00;
            reg_file[20757] <= 8'h00;
            reg_file[20758] <= 8'h00;
            reg_file[20759] <= 8'h00;
            reg_file[20760] <= 8'h00;
            reg_file[20761] <= 8'h00;
            reg_file[20762] <= 8'h00;
            reg_file[20763] <= 8'h00;
            reg_file[20764] <= 8'h00;
            reg_file[20765] <= 8'h00;
            reg_file[20766] <= 8'h00;
            reg_file[20767] <= 8'h00;
            reg_file[20768] <= 8'h00;
            reg_file[20769] <= 8'h00;
            reg_file[20770] <= 8'h00;
            reg_file[20771] <= 8'h00;
            reg_file[20772] <= 8'h00;
            reg_file[20773] <= 8'h00;
            reg_file[20774] <= 8'h00;
            reg_file[20775] <= 8'h00;
            reg_file[20776] <= 8'h00;
            reg_file[20777] <= 8'h00;
            reg_file[20778] <= 8'h00;
            reg_file[20779] <= 8'h00;
            reg_file[20780] <= 8'h00;
            reg_file[20781] <= 8'h00;
            reg_file[20782] <= 8'h00;
            reg_file[20783] <= 8'h00;
            reg_file[20784] <= 8'h00;
            reg_file[20785] <= 8'h00;
            reg_file[20786] <= 8'h00;
            reg_file[20787] <= 8'h00;
            reg_file[20788] <= 8'h00;
            reg_file[20789] <= 8'h00;
            reg_file[20790] <= 8'h00;
            reg_file[20791] <= 8'h00;
            reg_file[20792] <= 8'h00;
            reg_file[20793] <= 8'h00;
            reg_file[20794] <= 8'h00;
            reg_file[20795] <= 8'h00;
            reg_file[20796] <= 8'h00;
            reg_file[20797] <= 8'h00;
            reg_file[20798] <= 8'h00;
            reg_file[20799] <= 8'h00;
            reg_file[20800] <= 8'h00;
            reg_file[20801] <= 8'h00;
            reg_file[20802] <= 8'h00;
            reg_file[20803] <= 8'h00;
            reg_file[20804] <= 8'h00;
            reg_file[20805] <= 8'h00;
            reg_file[20806] <= 8'h00;
            reg_file[20807] <= 8'h00;
            reg_file[20808] <= 8'h00;
            reg_file[20809] <= 8'h00;
            reg_file[20810] <= 8'h00;
            reg_file[20811] <= 8'h00;
            reg_file[20812] <= 8'h00;
            reg_file[20813] <= 8'h00;
            reg_file[20814] <= 8'h00;
            reg_file[20815] <= 8'h00;
            reg_file[20816] <= 8'h00;
            reg_file[20817] <= 8'h00;
            reg_file[20818] <= 8'h00;
            reg_file[20819] <= 8'h00;
            reg_file[20820] <= 8'h00;
            reg_file[20821] <= 8'h00;
            reg_file[20822] <= 8'h00;
            reg_file[20823] <= 8'h00;
            reg_file[20824] <= 8'h00;
            reg_file[20825] <= 8'h00;
            reg_file[20826] <= 8'h00;
            reg_file[20827] <= 8'h00;
            reg_file[20828] <= 8'h00;
            reg_file[20829] <= 8'h00;
            reg_file[20830] <= 8'h00;
            reg_file[20831] <= 8'h00;
            reg_file[20832] <= 8'h00;
            reg_file[20833] <= 8'h00;
            reg_file[20834] <= 8'h00;
            reg_file[20835] <= 8'h00;
            reg_file[20836] <= 8'h00;
            reg_file[20837] <= 8'h00;
            reg_file[20838] <= 8'h00;
            reg_file[20839] <= 8'h00;
            reg_file[20840] <= 8'h00;
            reg_file[20841] <= 8'h00;
            reg_file[20842] <= 8'h00;
            reg_file[20843] <= 8'h00;
            reg_file[20844] <= 8'h00;
            reg_file[20845] <= 8'h00;
            reg_file[20846] <= 8'h00;
            reg_file[20847] <= 8'h00;
            reg_file[20848] <= 8'h00;
            reg_file[20849] <= 8'h00;
            reg_file[20850] <= 8'h00;
            reg_file[20851] <= 8'h00;
            reg_file[20852] <= 8'h00;
            reg_file[20853] <= 8'h00;
            reg_file[20854] <= 8'h00;
            reg_file[20855] <= 8'h00;
            reg_file[20856] <= 8'h00;
            reg_file[20857] <= 8'h00;
            reg_file[20858] <= 8'h00;
            reg_file[20859] <= 8'h00;
            reg_file[20860] <= 8'h00;
            reg_file[20861] <= 8'h00;
            reg_file[20862] <= 8'h00;
            reg_file[20863] <= 8'h00;
            reg_file[20864] <= 8'h00;
            reg_file[20865] <= 8'h00;
            reg_file[20866] <= 8'h00;
            reg_file[20867] <= 8'h00;
            reg_file[20868] <= 8'h00;
            reg_file[20869] <= 8'h00;
            reg_file[20870] <= 8'h00;
            reg_file[20871] <= 8'h00;
            reg_file[20872] <= 8'h00;
            reg_file[20873] <= 8'h00;
            reg_file[20874] <= 8'h00;
            reg_file[20875] <= 8'h00;
            reg_file[20876] <= 8'h00;
            reg_file[20877] <= 8'h00;
            reg_file[20878] <= 8'h00;
            reg_file[20879] <= 8'h00;
            reg_file[20880] <= 8'h00;
            reg_file[20881] <= 8'h00;
            reg_file[20882] <= 8'h00;
            reg_file[20883] <= 8'h00;
            reg_file[20884] <= 8'h00;
            reg_file[20885] <= 8'h00;
            reg_file[20886] <= 8'h00;
            reg_file[20887] <= 8'h00;
            reg_file[20888] <= 8'h00;
            reg_file[20889] <= 8'h00;
            reg_file[20890] <= 8'h00;
            reg_file[20891] <= 8'h00;
            reg_file[20892] <= 8'h00;
            reg_file[20893] <= 8'h00;
            reg_file[20894] <= 8'h00;
            reg_file[20895] <= 8'h00;
            reg_file[20896] <= 8'h00;
            reg_file[20897] <= 8'h00;
            reg_file[20898] <= 8'h00;
            reg_file[20899] <= 8'h00;
            reg_file[20900] <= 8'h00;
            reg_file[20901] <= 8'h00;
            reg_file[20902] <= 8'h00;
            reg_file[20903] <= 8'h00;
            reg_file[20904] <= 8'h00;
            reg_file[20905] <= 8'h00;
            reg_file[20906] <= 8'h00;
            reg_file[20907] <= 8'h00;
            reg_file[20908] <= 8'h00;
            reg_file[20909] <= 8'h00;
            reg_file[20910] <= 8'h00;
            reg_file[20911] <= 8'h00;
            reg_file[20912] <= 8'h00;
            reg_file[20913] <= 8'h00;
            reg_file[20914] <= 8'h00;
            reg_file[20915] <= 8'h00;
            reg_file[20916] <= 8'h00;
            reg_file[20917] <= 8'h00;
            reg_file[20918] <= 8'h00;
            reg_file[20919] <= 8'h00;
            reg_file[20920] <= 8'h00;
            reg_file[20921] <= 8'h00;
            reg_file[20922] <= 8'h00;
            reg_file[20923] <= 8'h00;
            reg_file[20924] <= 8'h00;
            reg_file[20925] <= 8'h00;
            reg_file[20926] <= 8'h00;
            reg_file[20927] <= 8'h00;
            reg_file[20928] <= 8'h00;
            reg_file[20929] <= 8'h00;
            reg_file[20930] <= 8'h00;
            reg_file[20931] <= 8'h00;
            reg_file[20932] <= 8'h00;
            reg_file[20933] <= 8'h00;
            reg_file[20934] <= 8'h00;
            reg_file[20935] <= 8'h00;
            reg_file[20936] <= 8'h00;
            reg_file[20937] <= 8'h00;
            reg_file[20938] <= 8'h00;
            reg_file[20939] <= 8'h00;
            reg_file[20940] <= 8'h00;
            reg_file[20941] <= 8'h00;
            reg_file[20942] <= 8'h00;
            reg_file[20943] <= 8'h00;
            reg_file[20944] <= 8'h00;
            reg_file[20945] <= 8'h00;
            reg_file[20946] <= 8'h00;
            reg_file[20947] <= 8'h00;
            reg_file[20948] <= 8'h00;
            reg_file[20949] <= 8'h00;
            reg_file[20950] <= 8'h00;
            reg_file[20951] <= 8'h00;
            reg_file[20952] <= 8'h00;
            reg_file[20953] <= 8'h00;
            reg_file[20954] <= 8'h00;
            reg_file[20955] <= 8'h00;
            reg_file[20956] <= 8'h00;
            reg_file[20957] <= 8'h00;
            reg_file[20958] <= 8'h00;
            reg_file[20959] <= 8'h00;
            reg_file[20960] <= 8'h00;
            reg_file[20961] <= 8'h00;
            reg_file[20962] <= 8'h00;
            reg_file[20963] <= 8'h00;
            reg_file[20964] <= 8'h00;
            reg_file[20965] <= 8'h00;
            reg_file[20966] <= 8'h00;
            reg_file[20967] <= 8'h00;
            reg_file[20968] <= 8'h00;
            reg_file[20969] <= 8'h00;
            reg_file[20970] <= 8'h00;
            reg_file[20971] <= 8'h00;
            reg_file[20972] <= 8'h00;
            reg_file[20973] <= 8'h00;
            reg_file[20974] <= 8'h00;
            reg_file[20975] <= 8'h00;
            reg_file[20976] <= 8'h00;
            reg_file[20977] <= 8'h00;
            reg_file[20978] <= 8'h00;
            reg_file[20979] <= 8'h00;
            reg_file[20980] <= 8'h00;
            reg_file[20981] <= 8'h00;
            reg_file[20982] <= 8'h00;
            reg_file[20983] <= 8'h00;
            reg_file[20984] <= 8'h00;
            reg_file[20985] <= 8'h00;
            reg_file[20986] <= 8'h00;
            reg_file[20987] <= 8'h00;
            reg_file[20988] <= 8'h00;
            reg_file[20989] <= 8'h00;
            reg_file[20990] <= 8'h00;
            reg_file[20991] <= 8'h00;
            reg_file[20992] <= 8'h00;
            reg_file[20993] <= 8'h00;
            reg_file[20994] <= 8'h00;
            reg_file[20995] <= 8'h00;
            reg_file[20996] <= 8'h00;
            reg_file[20997] <= 8'h00;
            reg_file[20998] <= 8'h00;
            reg_file[20999] <= 8'h00;
            reg_file[21000] <= 8'h00;
            reg_file[21001] <= 8'h00;
            reg_file[21002] <= 8'h00;
            reg_file[21003] <= 8'h00;
            reg_file[21004] <= 8'h00;
            reg_file[21005] <= 8'h00;
            reg_file[21006] <= 8'h00;
            reg_file[21007] <= 8'h00;
            reg_file[21008] <= 8'h00;
            reg_file[21009] <= 8'h00;
            reg_file[21010] <= 8'h00;
            reg_file[21011] <= 8'h00;
            reg_file[21012] <= 8'h00;
            reg_file[21013] <= 8'h00;
            reg_file[21014] <= 8'h00;
            reg_file[21015] <= 8'h00;
            reg_file[21016] <= 8'h00;
            reg_file[21017] <= 8'h00;
            reg_file[21018] <= 8'h00;
            reg_file[21019] <= 8'h00;
            reg_file[21020] <= 8'h00;
            reg_file[21021] <= 8'h00;
            reg_file[21022] <= 8'h00;
            reg_file[21023] <= 8'h00;
            reg_file[21024] <= 8'h00;
            reg_file[21025] <= 8'h00;
            reg_file[21026] <= 8'h00;
            reg_file[21027] <= 8'h00;
            reg_file[21028] <= 8'h00;
            reg_file[21029] <= 8'h00;
            reg_file[21030] <= 8'h00;
            reg_file[21031] <= 8'h00;
            reg_file[21032] <= 8'h00;
            reg_file[21033] <= 8'h00;
            reg_file[21034] <= 8'h00;
            reg_file[21035] <= 8'h00;
            reg_file[21036] <= 8'h00;
            reg_file[21037] <= 8'h00;
            reg_file[21038] <= 8'h00;
            reg_file[21039] <= 8'h00;
            reg_file[21040] <= 8'h00;
            reg_file[21041] <= 8'h00;
            reg_file[21042] <= 8'h00;
            reg_file[21043] <= 8'h00;
            reg_file[21044] <= 8'h00;
            reg_file[21045] <= 8'h00;
            reg_file[21046] <= 8'h00;
            reg_file[21047] <= 8'h00;
            reg_file[21048] <= 8'h00;
            reg_file[21049] <= 8'h00;
            reg_file[21050] <= 8'h00;
            reg_file[21051] <= 8'h00;
            reg_file[21052] <= 8'h00;
            reg_file[21053] <= 8'h00;
            reg_file[21054] <= 8'h00;
            reg_file[21055] <= 8'h00;
            reg_file[21056] <= 8'h00;
            reg_file[21057] <= 8'h00;
            reg_file[21058] <= 8'h00;
            reg_file[21059] <= 8'h00;
            reg_file[21060] <= 8'h00;
            reg_file[21061] <= 8'h00;
            reg_file[21062] <= 8'h00;
            reg_file[21063] <= 8'h00;
            reg_file[21064] <= 8'h00;
            reg_file[21065] <= 8'h00;
            reg_file[21066] <= 8'h00;
            reg_file[21067] <= 8'h00;
            reg_file[21068] <= 8'h00;
            reg_file[21069] <= 8'h00;
            reg_file[21070] <= 8'h00;
            reg_file[21071] <= 8'h00;
            reg_file[21072] <= 8'h00;
            reg_file[21073] <= 8'h00;
            reg_file[21074] <= 8'h00;
            reg_file[21075] <= 8'h00;
            reg_file[21076] <= 8'h00;
            reg_file[21077] <= 8'h00;
            reg_file[21078] <= 8'h00;
            reg_file[21079] <= 8'h00;
            reg_file[21080] <= 8'h00;
            reg_file[21081] <= 8'h00;
            reg_file[21082] <= 8'h00;
            reg_file[21083] <= 8'h00;
            reg_file[21084] <= 8'h00;
            reg_file[21085] <= 8'h00;
            reg_file[21086] <= 8'h00;
            reg_file[21087] <= 8'h00;
            reg_file[21088] <= 8'h00;
            reg_file[21089] <= 8'h00;
            reg_file[21090] <= 8'h00;
            reg_file[21091] <= 8'h00;
            reg_file[21092] <= 8'h00;
            reg_file[21093] <= 8'h00;
            reg_file[21094] <= 8'h00;
            reg_file[21095] <= 8'h00;
            reg_file[21096] <= 8'h00;
            reg_file[21097] <= 8'h00;
            reg_file[21098] <= 8'h00;
            reg_file[21099] <= 8'h00;
            reg_file[21100] <= 8'h00;
            reg_file[21101] <= 8'h00;
            reg_file[21102] <= 8'h00;
            reg_file[21103] <= 8'h00;
            reg_file[21104] <= 8'h00;
            reg_file[21105] <= 8'h00;
            reg_file[21106] <= 8'h00;
            reg_file[21107] <= 8'h00;
            reg_file[21108] <= 8'h00;
            reg_file[21109] <= 8'h00;
            reg_file[21110] <= 8'h00;
            reg_file[21111] <= 8'h00;
            reg_file[21112] <= 8'h00;
            reg_file[21113] <= 8'h00;
            reg_file[21114] <= 8'h00;
            reg_file[21115] <= 8'h00;
            reg_file[21116] <= 8'h00;
            reg_file[21117] <= 8'h00;
            reg_file[21118] <= 8'h00;
            reg_file[21119] <= 8'h00;
            reg_file[21120] <= 8'h00;
            reg_file[21121] <= 8'h00;
            reg_file[21122] <= 8'h00;
            reg_file[21123] <= 8'h00;
            reg_file[21124] <= 8'h00;
            reg_file[21125] <= 8'h00;
            reg_file[21126] <= 8'h00;
            reg_file[21127] <= 8'h00;
            reg_file[21128] <= 8'h00;
            reg_file[21129] <= 8'h00;
            reg_file[21130] <= 8'h00;
            reg_file[21131] <= 8'h00;
            reg_file[21132] <= 8'h00;
            reg_file[21133] <= 8'h00;
            reg_file[21134] <= 8'h00;
            reg_file[21135] <= 8'h00;
            reg_file[21136] <= 8'h00;
            reg_file[21137] <= 8'h00;
            reg_file[21138] <= 8'h00;
            reg_file[21139] <= 8'h00;
            reg_file[21140] <= 8'h00;
            reg_file[21141] <= 8'h00;
            reg_file[21142] <= 8'h00;
            reg_file[21143] <= 8'h00;
            reg_file[21144] <= 8'h00;
            reg_file[21145] <= 8'h00;
            reg_file[21146] <= 8'h00;
            reg_file[21147] <= 8'h00;
            reg_file[21148] <= 8'h00;
            reg_file[21149] <= 8'h00;
            reg_file[21150] <= 8'h00;
            reg_file[21151] <= 8'h00;
            reg_file[21152] <= 8'h00;
            reg_file[21153] <= 8'h00;
            reg_file[21154] <= 8'h00;
            reg_file[21155] <= 8'h00;
            reg_file[21156] <= 8'h00;
            reg_file[21157] <= 8'h00;
            reg_file[21158] <= 8'h00;
            reg_file[21159] <= 8'h00;
            reg_file[21160] <= 8'h00;
            reg_file[21161] <= 8'h00;
            reg_file[21162] <= 8'h00;
            reg_file[21163] <= 8'h00;
            reg_file[21164] <= 8'h00;
            reg_file[21165] <= 8'h00;
            reg_file[21166] <= 8'h00;
            reg_file[21167] <= 8'h00;
            reg_file[21168] <= 8'h00;
            reg_file[21169] <= 8'h00;
            reg_file[21170] <= 8'h00;
            reg_file[21171] <= 8'h00;
            reg_file[21172] <= 8'h00;
            reg_file[21173] <= 8'h00;
            reg_file[21174] <= 8'h00;
            reg_file[21175] <= 8'h00;
            reg_file[21176] <= 8'h00;
            reg_file[21177] <= 8'h00;
            reg_file[21178] <= 8'h00;
            reg_file[21179] <= 8'h00;
            reg_file[21180] <= 8'h00;
            reg_file[21181] <= 8'h00;
            reg_file[21182] <= 8'h00;
            reg_file[21183] <= 8'h00;
            reg_file[21184] <= 8'h00;
            reg_file[21185] <= 8'h00;
            reg_file[21186] <= 8'h00;
            reg_file[21187] <= 8'h00;
            reg_file[21188] <= 8'h00;
            reg_file[21189] <= 8'h00;
            reg_file[21190] <= 8'h00;
            reg_file[21191] <= 8'h00;
            reg_file[21192] <= 8'h00;
            reg_file[21193] <= 8'h00;
            reg_file[21194] <= 8'h00;
            reg_file[21195] <= 8'h00;
            reg_file[21196] <= 8'h00;
            reg_file[21197] <= 8'h00;
            reg_file[21198] <= 8'h00;
            reg_file[21199] <= 8'h00;
            reg_file[21200] <= 8'h00;
            reg_file[21201] <= 8'h00;
            reg_file[21202] <= 8'h00;
            reg_file[21203] <= 8'h00;
            reg_file[21204] <= 8'h00;
            reg_file[21205] <= 8'h00;
            reg_file[21206] <= 8'h00;
            reg_file[21207] <= 8'h00;
            reg_file[21208] <= 8'h00;
            reg_file[21209] <= 8'h00;
            reg_file[21210] <= 8'h00;
            reg_file[21211] <= 8'h00;
            reg_file[21212] <= 8'h00;
            reg_file[21213] <= 8'h00;
            reg_file[21214] <= 8'h00;
            reg_file[21215] <= 8'h00;
            reg_file[21216] <= 8'h00;
            reg_file[21217] <= 8'h00;
            reg_file[21218] <= 8'h00;
            reg_file[21219] <= 8'h00;
            reg_file[21220] <= 8'h00;
            reg_file[21221] <= 8'h00;
            reg_file[21222] <= 8'h00;
            reg_file[21223] <= 8'h00;
            reg_file[21224] <= 8'h00;
            reg_file[21225] <= 8'h00;
            reg_file[21226] <= 8'h00;
            reg_file[21227] <= 8'h00;
            reg_file[21228] <= 8'h00;
            reg_file[21229] <= 8'h00;
            reg_file[21230] <= 8'h00;
            reg_file[21231] <= 8'h00;
            reg_file[21232] <= 8'h00;
            reg_file[21233] <= 8'h00;
            reg_file[21234] <= 8'h00;
            reg_file[21235] <= 8'h00;
            reg_file[21236] <= 8'h00;
            reg_file[21237] <= 8'h00;
            reg_file[21238] <= 8'h00;
            reg_file[21239] <= 8'h00;
            reg_file[21240] <= 8'h00;
            reg_file[21241] <= 8'h00;
            reg_file[21242] <= 8'h00;
            reg_file[21243] <= 8'h00;
            reg_file[21244] <= 8'h00;
            reg_file[21245] <= 8'h00;
            reg_file[21246] <= 8'h00;
            reg_file[21247] <= 8'h00;
            reg_file[21248] <= 8'h00;
            reg_file[21249] <= 8'h00;
            reg_file[21250] <= 8'h00;
            reg_file[21251] <= 8'h00;
            reg_file[21252] <= 8'h00;
            reg_file[21253] <= 8'h00;
            reg_file[21254] <= 8'h00;
            reg_file[21255] <= 8'h00;
            reg_file[21256] <= 8'h00;
            reg_file[21257] <= 8'h00;
            reg_file[21258] <= 8'h00;
            reg_file[21259] <= 8'h00;
            reg_file[21260] <= 8'h00;
            reg_file[21261] <= 8'h00;
            reg_file[21262] <= 8'h00;
            reg_file[21263] <= 8'h00;
            reg_file[21264] <= 8'h00;
            reg_file[21265] <= 8'h00;
            reg_file[21266] <= 8'h00;
            reg_file[21267] <= 8'h00;
            reg_file[21268] <= 8'h00;
            reg_file[21269] <= 8'h00;
            reg_file[21270] <= 8'h00;
            reg_file[21271] <= 8'h00;
            reg_file[21272] <= 8'h00;
            reg_file[21273] <= 8'h00;
            reg_file[21274] <= 8'h00;
            reg_file[21275] <= 8'h00;
            reg_file[21276] <= 8'h00;
            reg_file[21277] <= 8'h00;
            reg_file[21278] <= 8'h00;
            reg_file[21279] <= 8'h00;
            reg_file[21280] <= 8'h00;
            reg_file[21281] <= 8'h00;
            reg_file[21282] <= 8'h00;
            reg_file[21283] <= 8'h00;
            reg_file[21284] <= 8'h00;
            reg_file[21285] <= 8'h00;
            reg_file[21286] <= 8'h00;
            reg_file[21287] <= 8'h00;
            reg_file[21288] <= 8'h00;
            reg_file[21289] <= 8'h00;
            reg_file[21290] <= 8'h00;
            reg_file[21291] <= 8'h00;
            reg_file[21292] <= 8'h00;
            reg_file[21293] <= 8'h00;
            reg_file[21294] <= 8'h00;
            reg_file[21295] <= 8'h00;
            reg_file[21296] <= 8'h00;
            reg_file[21297] <= 8'h00;
            reg_file[21298] <= 8'h00;
            reg_file[21299] <= 8'h00;
            reg_file[21300] <= 8'h00;
            reg_file[21301] <= 8'h00;
            reg_file[21302] <= 8'h00;
            reg_file[21303] <= 8'h00;
            reg_file[21304] <= 8'h00;
            reg_file[21305] <= 8'h00;
            reg_file[21306] <= 8'h00;
            reg_file[21307] <= 8'h00;
            reg_file[21308] <= 8'h00;
            reg_file[21309] <= 8'h00;
            reg_file[21310] <= 8'h00;
            reg_file[21311] <= 8'h00;
            reg_file[21312] <= 8'h00;
            reg_file[21313] <= 8'h00;
            reg_file[21314] <= 8'h00;
            reg_file[21315] <= 8'h00;
            reg_file[21316] <= 8'h00;
            reg_file[21317] <= 8'h00;
            reg_file[21318] <= 8'h00;
            reg_file[21319] <= 8'h00;
            reg_file[21320] <= 8'h00;
            reg_file[21321] <= 8'h00;
            reg_file[21322] <= 8'h00;
            reg_file[21323] <= 8'h00;
            reg_file[21324] <= 8'h00;
            reg_file[21325] <= 8'h00;
            reg_file[21326] <= 8'h00;
            reg_file[21327] <= 8'h00;
            reg_file[21328] <= 8'h00;
            reg_file[21329] <= 8'h00;
            reg_file[21330] <= 8'h00;
            reg_file[21331] <= 8'h00;
            reg_file[21332] <= 8'h00;
            reg_file[21333] <= 8'h00;
            reg_file[21334] <= 8'h00;
            reg_file[21335] <= 8'h00;
            reg_file[21336] <= 8'h00;
            reg_file[21337] <= 8'h00;
            reg_file[21338] <= 8'h00;
            reg_file[21339] <= 8'h00;
            reg_file[21340] <= 8'h00;
            reg_file[21341] <= 8'h00;
            reg_file[21342] <= 8'h00;
            reg_file[21343] <= 8'h00;
            reg_file[21344] <= 8'h00;
            reg_file[21345] <= 8'h00;
            reg_file[21346] <= 8'h00;
            reg_file[21347] <= 8'h00;
            reg_file[21348] <= 8'h00;
            reg_file[21349] <= 8'h00;
            reg_file[21350] <= 8'h00;
            reg_file[21351] <= 8'h00;
            reg_file[21352] <= 8'h00;
            reg_file[21353] <= 8'h00;
            reg_file[21354] <= 8'h00;
            reg_file[21355] <= 8'h00;
            reg_file[21356] <= 8'h00;
            reg_file[21357] <= 8'h00;
            reg_file[21358] <= 8'h00;
            reg_file[21359] <= 8'h00;
            reg_file[21360] <= 8'h00;
            reg_file[21361] <= 8'h00;
            reg_file[21362] <= 8'h00;
            reg_file[21363] <= 8'h00;
            reg_file[21364] <= 8'h00;
            reg_file[21365] <= 8'h00;
            reg_file[21366] <= 8'h00;
            reg_file[21367] <= 8'h00;
            reg_file[21368] <= 8'h00;
            reg_file[21369] <= 8'h00;
            reg_file[21370] <= 8'h00;
            reg_file[21371] <= 8'h00;
            reg_file[21372] <= 8'h00;
            reg_file[21373] <= 8'h00;
            reg_file[21374] <= 8'h00;
            reg_file[21375] <= 8'h00;
            reg_file[21376] <= 8'h00;
            reg_file[21377] <= 8'h00;
            reg_file[21378] <= 8'h00;
            reg_file[21379] <= 8'h00;
            reg_file[21380] <= 8'h00;
            reg_file[21381] <= 8'h00;
            reg_file[21382] <= 8'h00;
            reg_file[21383] <= 8'h00;
            reg_file[21384] <= 8'h00;
            reg_file[21385] <= 8'h00;
            reg_file[21386] <= 8'h00;
            reg_file[21387] <= 8'h00;
            reg_file[21388] <= 8'h00;
            reg_file[21389] <= 8'h00;
            reg_file[21390] <= 8'h00;
            reg_file[21391] <= 8'h00;
            reg_file[21392] <= 8'h00;
            reg_file[21393] <= 8'h00;
            reg_file[21394] <= 8'h00;
            reg_file[21395] <= 8'h00;
            reg_file[21396] <= 8'h00;
            reg_file[21397] <= 8'h00;
            reg_file[21398] <= 8'h00;
            reg_file[21399] <= 8'h00;
            reg_file[21400] <= 8'h00;
            reg_file[21401] <= 8'h00;
            reg_file[21402] <= 8'h00;
            reg_file[21403] <= 8'h00;
            reg_file[21404] <= 8'h00;
            reg_file[21405] <= 8'h00;
            reg_file[21406] <= 8'h00;
            reg_file[21407] <= 8'h00;
            reg_file[21408] <= 8'h00;
            reg_file[21409] <= 8'h00;
            reg_file[21410] <= 8'h00;
            reg_file[21411] <= 8'h00;
            reg_file[21412] <= 8'h00;
            reg_file[21413] <= 8'h00;
            reg_file[21414] <= 8'h00;
            reg_file[21415] <= 8'h00;
            reg_file[21416] <= 8'h00;
            reg_file[21417] <= 8'h00;
            reg_file[21418] <= 8'h00;
            reg_file[21419] <= 8'h00;
            reg_file[21420] <= 8'h00;
            reg_file[21421] <= 8'h00;
            reg_file[21422] <= 8'h00;
            reg_file[21423] <= 8'h00;
            reg_file[21424] <= 8'h00;
            reg_file[21425] <= 8'h00;
            reg_file[21426] <= 8'h00;
            reg_file[21427] <= 8'h00;
            reg_file[21428] <= 8'h00;
            reg_file[21429] <= 8'h00;
            reg_file[21430] <= 8'h00;
            reg_file[21431] <= 8'h00;
            reg_file[21432] <= 8'h00;
            reg_file[21433] <= 8'h00;
            reg_file[21434] <= 8'h00;
            reg_file[21435] <= 8'h00;
            reg_file[21436] <= 8'h00;
            reg_file[21437] <= 8'h00;
            reg_file[21438] <= 8'h00;
            reg_file[21439] <= 8'h00;
            reg_file[21440] <= 8'h00;
            reg_file[21441] <= 8'h00;
            reg_file[21442] <= 8'h00;
            reg_file[21443] <= 8'h00;
            reg_file[21444] <= 8'h00;
            reg_file[21445] <= 8'h00;
            reg_file[21446] <= 8'h00;
            reg_file[21447] <= 8'h00;
            reg_file[21448] <= 8'h00;
            reg_file[21449] <= 8'h00;
            reg_file[21450] <= 8'h00;
            reg_file[21451] <= 8'h00;
            reg_file[21452] <= 8'h00;
            reg_file[21453] <= 8'h00;
            reg_file[21454] <= 8'h00;
            reg_file[21455] <= 8'h00;
            reg_file[21456] <= 8'h00;
            reg_file[21457] <= 8'h00;
            reg_file[21458] <= 8'h00;
            reg_file[21459] <= 8'h00;
            reg_file[21460] <= 8'h00;
            reg_file[21461] <= 8'h00;
            reg_file[21462] <= 8'h00;
            reg_file[21463] <= 8'h00;
            reg_file[21464] <= 8'h00;
            reg_file[21465] <= 8'h00;
            reg_file[21466] <= 8'h00;
            reg_file[21467] <= 8'h00;
            reg_file[21468] <= 8'h00;
            reg_file[21469] <= 8'h00;
            reg_file[21470] <= 8'h00;
            reg_file[21471] <= 8'h00;
            reg_file[21472] <= 8'h00;
            reg_file[21473] <= 8'h00;
            reg_file[21474] <= 8'h00;
            reg_file[21475] <= 8'h00;
            reg_file[21476] <= 8'h00;
            reg_file[21477] <= 8'h00;
            reg_file[21478] <= 8'h00;
            reg_file[21479] <= 8'h00;
            reg_file[21480] <= 8'h00;
            reg_file[21481] <= 8'h00;
            reg_file[21482] <= 8'h00;
            reg_file[21483] <= 8'h00;
            reg_file[21484] <= 8'h00;
            reg_file[21485] <= 8'h00;
            reg_file[21486] <= 8'h00;
            reg_file[21487] <= 8'h00;
            reg_file[21488] <= 8'h00;
            reg_file[21489] <= 8'h00;
            reg_file[21490] <= 8'h00;
            reg_file[21491] <= 8'h00;
            reg_file[21492] <= 8'h00;
            reg_file[21493] <= 8'h00;
            reg_file[21494] <= 8'h00;
            reg_file[21495] <= 8'h00;
            reg_file[21496] <= 8'h00;
            reg_file[21497] <= 8'h00;
            reg_file[21498] <= 8'h00;
            reg_file[21499] <= 8'h00;
            reg_file[21500] <= 8'h00;
            reg_file[21501] <= 8'h00;
            reg_file[21502] <= 8'h00;
            reg_file[21503] <= 8'h00;
            reg_file[21504] <= 8'h00;
            reg_file[21505] <= 8'h00;
            reg_file[21506] <= 8'h00;
            reg_file[21507] <= 8'h00;
            reg_file[21508] <= 8'h00;
            reg_file[21509] <= 8'h00;
            reg_file[21510] <= 8'h00;
            reg_file[21511] <= 8'h00;
            reg_file[21512] <= 8'h00;
            reg_file[21513] <= 8'h00;
            reg_file[21514] <= 8'h00;
            reg_file[21515] <= 8'h00;
            reg_file[21516] <= 8'h00;
            reg_file[21517] <= 8'h00;
            reg_file[21518] <= 8'h00;
            reg_file[21519] <= 8'h00;
            reg_file[21520] <= 8'h00;
            reg_file[21521] <= 8'h00;
            reg_file[21522] <= 8'h00;
            reg_file[21523] <= 8'h00;
            reg_file[21524] <= 8'h00;
            reg_file[21525] <= 8'h00;
            reg_file[21526] <= 8'h00;
            reg_file[21527] <= 8'h00;
            reg_file[21528] <= 8'h00;
            reg_file[21529] <= 8'h00;
            reg_file[21530] <= 8'h00;
            reg_file[21531] <= 8'h00;
            reg_file[21532] <= 8'h00;
            reg_file[21533] <= 8'h00;
            reg_file[21534] <= 8'h00;
            reg_file[21535] <= 8'h00;
            reg_file[21536] <= 8'h00;
            reg_file[21537] <= 8'h00;
            reg_file[21538] <= 8'h00;
            reg_file[21539] <= 8'h00;
            reg_file[21540] <= 8'h00;
            reg_file[21541] <= 8'h00;
            reg_file[21542] <= 8'h00;
            reg_file[21543] <= 8'h00;
            reg_file[21544] <= 8'h00;
            reg_file[21545] <= 8'h00;
            reg_file[21546] <= 8'h00;
            reg_file[21547] <= 8'h00;
            reg_file[21548] <= 8'h00;
            reg_file[21549] <= 8'h00;
            reg_file[21550] <= 8'h00;
            reg_file[21551] <= 8'h00;
            reg_file[21552] <= 8'h00;
            reg_file[21553] <= 8'h00;
            reg_file[21554] <= 8'h00;
            reg_file[21555] <= 8'h00;
            reg_file[21556] <= 8'h00;
            reg_file[21557] <= 8'h00;
            reg_file[21558] <= 8'h00;
            reg_file[21559] <= 8'h00;
            reg_file[21560] <= 8'h00;
            reg_file[21561] <= 8'h00;
            reg_file[21562] <= 8'h00;
            reg_file[21563] <= 8'h00;
            reg_file[21564] <= 8'h00;
            reg_file[21565] <= 8'h00;
            reg_file[21566] <= 8'h00;
            reg_file[21567] <= 8'h00;
            reg_file[21568] <= 8'h00;
            reg_file[21569] <= 8'h00;
            reg_file[21570] <= 8'h00;
            reg_file[21571] <= 8'h00;
            reg_file[21572] <= 8'h00;
            reg_file[21573] <= 8'h00;
            reg_file[21574] <= 8'h00;
            reg_file[21575] <= 8'h00;
            reg_file[21576] <= 8'h00;
            reg_file[21577] <= 8'h00;
            reg_file[21578] <= 8'h00;
            reg_file[21579] <= 8'h00;
            reg_file[21580] <= 8'h00;
            reg_file[21581] <= 8'h00;
            reg_file[21582] <= 8'h00;
            reg_file[21583] <= 8'h00;
            reg_file[21584] <= 8'h00;
            reg_file[21585] <= 8'h00;
            reg_file[21586] <= 8'h00;
            reg_file[21587] <= 8'h00;
            reg_file[21588] <= 8'h00;
            reg_file[21589] <= 8'h00;
            reg_file[21590] <= 8'h00;
            reg_file[21591] <= 8'h00;
            reg_file[21592] <= 8'h00;
            reg_file[21593] <= 8'h00;
            reg_file[21594] <= 8'h00;
            reg_file[21595] <= 8'h00;
            reg_file[21596] <= 8'h00;
            reg_file[21597] <= 8'h00;
            reg_file[21598] <= 8'h00;
            reg_file[21599] <= 8'h00;
            reg_file[21600] <= 8'h00;
            reg_file[21601] <= 8'h00;
            reg_file[21602] <= 8'h00;
            reg_file[21603] <= 8'h00;
            reg_file[21604] <= 8'h00;
            reg_file[21605] <= 8'h00;
            reg_file[21606] <= 8'h00;
            reg_file[21607] <= 8'h00;
            reg_file[21608] <= 8'h00;
            reg_file[21609] <= 8'h00;
            reg_file[21610] <= 8'h00;
            reg_file[21611] <= 8'h00;
            reg_file[21612] <= 8'h00;
            reg_file[21613] <= 8'h00;
            reg_file[21614] <= 8'h00;
            reg_file[21615] <= 8'h00;
            reg_file[21616] <= 8'h00;
            reg_file[21617] <= 8'h00;
            reg_file[21618] <= 8'h00;
            reg_file[21619] <= 8'h00;
            reg_file[21620] <= 8'h00;
            reg_file[21621] <= 8'h00;
            reg_file[21622] <= 8'h00;
            reg_file[21623] <= 8'h00;
            reg_file[21624] <= 8'h00;
            reg_file[21625] <= 8'h00;
            reg_file[21626] <= 8'h00;
            reg_file[21627] <= 8'h00;
            reg_file[21628] <= 8'h00;
            reg_file[21629] <= 8'h00;
            reg_file[21630] <= 8'h00;
            reg_file[21631] <= 8'h00;
            reg_file[21632] <= 8'h00;
            reg_file[21633] <= 8'h00;
            reg_file[21634] <= 8'h00;
            reg_file[21635] <= 8'h00;
            reg_file[21636] <= 8'h00;
            reg_file[21637] <= 8'h00;
            reg_file[21638] <= 8'h00;
            reg_file[21639] <= 8'h00;
            reg_file[21640] <= 8'h00;
            reg_file[21641] <= 8'h00;
            reg_file[21642] <= 8'h00;
            reg_file[21643] <= 8'h00;
            reg_file[21644] <= 8'h00;
            reg_file[21645] <= 8'h00;
            reg_file[21646] <= 8'h00;
            reg_file[21647] <= 8'h00;
            reg_file[21648] <= 8'h00;
            reg_file[21649] <= 8'h00;
            reg_file[21650] <= 8'h00;
            reg_file[21651] <= 8'h00;
            reg_file[21652] <= 8'h00;
            reg_file[21653] <= 8'h00;
            reg_file[21654] <= 8'h00;
            reg_file[21655] <= 8'h00;
            reg_file[21656] <= 8'h00;
            reg_file[21657] <= 8'h00;
            reg_file[21658] <= 8'h00;
            reg_file[21659] <= 8'h00;
            reg_file[21660] <= 8'h00;
            reg_file[21661] <= 8'h00;
            reg_file[21662] <= 8'h00;
            reg_file[21663] <= 8'h00;
            reg_file[21664] <= 8'h00;
            reg_file[21665] <= 8'h00;
            reg_file[21666] <= 8'h00;
            reg_file[21667] <= 8'h00;
            reg_file[21668] <= 8'h00;
            reg_file[21669] <= 8'h00;
            reg_file[21670] <= 8'h00;
            reg_file[21671] <= 8'h00;
            reg_file[21672] <= 8'h00;
            reg_file[21673] <= 8'h00;
            reg_file[21674] <= 8'h00;
            reg_file[21675] <= 8'h00;
            reg_file[21676] <= 8'h00;
            reg_file[21677] <= 8'h00;
            reg_file[21678] <= 8'h00;
            reg_file[21679] <= 8'h00;
            reg_file[21680] <= 8'h00;
            reg_file[21681] <= 8'h00;
            reg_file[21682] <= 8'h00;
            reg_file[21683] <= 8'h00;
            reg_file[21684] <= 8'h00;
            reg_file[21685] <= 8'h00;
            reg_file[21686] <= 8'h00;
            reg_file[21687] <= 8'h00;
            reg_file[21688] <= 8'h00;
            reg_file[21689] <= 8'h00;
            reg_file[21690] <= 8'h00;
            reg_file[21691] <= 8'h00;
            reg_file[21692] <= 8'h00;
            reg_file[21693] <= 8'h00;
            reg_file[21694] <= 8'h00;
            reg_file[21695] <= 8'h00;
            reg_file[21696] <= 8'h00;
            reg_file[21697] <= 8'h00;
            reg_file[21698] <= 8'h00;
            reg_file[21699] <= 8'h00;
            reg_file[21700] <= 8'h00;
            reg_file[21701] <= 8'h00;
            reg_file[21702] <= 8'h00;
            reg_file[21703] <= 8'h00;
            reg_file[21704] <= 8'h00;
            reg_file[21705] <= 8'h00;
            reg_file[21706] <= 8'h00;
            reg_file[21707] <= 8'h00;
            reg_file[21708] <= 8'h00;
            reg_file[21709] <= 8'h00;
            reg_file[21710] <= 8'h00;
            reg_file[21711] <= 8'h00;
            reg_file[21712] <= 8'h00;
            reg_file[21713] <= 8'h00;
            reg_file[21714] <= 8'h00;
            reg_file[21715] <= 8'h00;
            reg_file[21716] <= 8'h00;
            reg_file[21717] <= 8'h00;
            reg_file[21718] <= 8'h00;
            reg_file[21719] <= 8'h00;
            reg_file[21720] <= 8'h00;
            reg_file[21721] <= 8'h00;
            reg_file[21722] <= 8'h00;
            reg_file[21723] <= 8'h00;
            reg_file[21724] <= 8'h00;
            reg_file[21725] <= 8'h00;
            reg_file[21726] <= 8'h00;
            reg_file[21727] <= 8'h00;
            reg_file[21728] <= 8'h00;
            reg_file[21729] <= 8'h00;
            reg_file[21730] <= 8'h00;
            reg_file[21731] <= 8'h00;
            reg_file[21732] <= 8'h00;
            reg_file[21733] <= 8'h00;
            reg_file[21734] <= 8'h00;
            reg_file[21735] <= 8'h00;
            reg_file[21736] <= 8'h00;
            reg_file[21737] <= 8'h00;
            reg_file[21738] <= 8'h00;
            reg_file[21739] <= 8'h00;
            reg_file[21740] <= 8'h00;
            reg_file[21741] <= 8'h00;
            reg_file[21742] <= 8'h00;
            reg_file[21743] <= 8'h00;
            reg_file[21744] <= 8'h00;
            reg_file[21745] <= 8'h00;
            reg_file[21746] <= 8'h00;
            reg_file[21747] <= 8'h00;
            reg_file[21748] <= 8'h00;
            reg_file[21749] <= 8'h00;
            reg_file[21750] <= 8'h00;
            reg_file[21751] <= 8'h00;
            reg_file[21752] <= 8'h00;
            reg_file[21753] <= 8'h00;
            reg_file[21754] <= 8'h00;
            reg_file[21755] <= 8'h00;
            reg_file[21756] <= 8'h00;
            reg_file[21757] <= 8'h00;
            reg_file[21758] <= 8'h00;
            reg_file[21759] <= 8'h00;
            reg_file[21760] <= 8'h00;
            reg_file[21761] <= 8'h00;
            reg_file[21762] <= 8'h00;
            reg_file[21763] <= 8'h00;
            reg_file[21764] <= 8'h00;
            reg_file[21765] <= 8'h00;
            reg_file[21766] <= 8'h00;
            reg_file[21767] <= 8'h00;
            reg_file[21768] <= 8'h00;
            reg_file[21769] <= 8'h00;
            reg_file[21770] <= 8'h00;
            reg_file[21771] <= 8'h00;
            reg_file[21772] <= 8'h00;
            reg_file[21773] <= 8'h00;
            reg_file[21774] <= 8'h00;
            reg_file[21775] <= 8'h00;
            reg_file[21776] <= 8'h00;
            reg_file[21777] <= 8'h00;
            reg_file[21778] <= 8'h00;
            reg_file[21779] <= 8'h00;
            reg_file[21780] <= 8'h00;
            reg_file[21781] <= 8'h00;
            reg_file[21782] <= 8'h00;
            reg_file[21783] <= 8'h00;
            reg_file[21784] <= 8'h00;
            reg_file[21785] <= 8'h00;
            reg_file[21786] <= 8'h00;
            reg_file[21787] <= 8'h00;
            reg_file[21788] <= 8'h00;
            reg_file[21789] <= 8'h00;
            reg_file[21790] <= 8'h00;
            reg_file[21791] <= 8'h00;
            reg_file[21792] <= 8'h00;
            reg_file[21793] <= 8'h00;
            reg_file[21794] <= 8'h00;
            reg_file[21795] <= 8'h00;
            reg_file[21796] <= 8'h00;
            reg_file[21797] <= 8'h00;
            reg_file[21798] <= 8'h00;
            reg_file[21799] <= 8'h00;
            reg_file[21800] <= 8'h00;
            reg_file[21801] <= 8'h00;
            reg_file[21802] <= 8'h00;
            reg_file[21803] <= 8'h00;
            reg_file[21804] <= 8'h00;
            reg_file[21805] <= 8'h00;
            reg_file[21806] <= 8'h00;
            reg_file[21807] <= 8'h00;
            reg_file[21808] <= 8'h00;
            reg_file[21809] <= 8'h00;
            reg_file[21810] <= 8'h00;
            reg_file[21811] <= 8'h00;
            reg_file[21812] <= 8'h00;
            reg_file[21813] <= 8'h00;
            reg_file[21814] <= 8'h00;
            reg_file[21815] <= 8'h00;
            reg_file[21816] <= 8'h00;
            reg_file[21817] <= 8'h00;
            reg_file[21818] <= 8'h00;
            reg_file[21819] <= 8'h00;
            reg_file[21820] <= 8'h00;
            reg_file[21821] <= 8'h00;
            reg_file[21822] <= 8'h00;
            reg_file[21823] <= 8'h00;
            reg_file[21824] <= 8'h00;
            reg_file[21825] <= 8'h00;
            reg_file[21826] <= 8'h00;
            reg_file[21827] <= 8'h00;
            reg_file[21828] <= 8'h00;
            reg_file[21829] <= 8'h00;
            reg_file[21830] <= 8'h00;
            reg_file[21831] <= 8'h00;
            reg_file[21832] <= 8'h00;
            reg_file[21833] <= 8'h00;
            reg_file[21834] <= 8'h00;
            reg_file[21835] <= 8'h00;
            reg_file[21836] <= 8'h00;
            reg_file[21837] <= 8'h00;
            reg_file[21838] <= 8'h00;
            reg_file[21839] <= 8'h00;
            reg_file[21840] <= 8'h00;
            reg_file[21841] <= 8'h00;
            reg_file[21842] <= 8'h00;
            reg_file[21843] <= 8'h00;
            reg_file[21844] <= 8'h00;
            reg_file[21845] <= 8'h00;
            reg_file[21846] <= 8'h00;
            reg_file[21847] <= 8'h00;
            reg_file[21848] <= 8'h00;
            reg_file[21849] <= 8'h00;
            reg_file[21850] <= 8'h00;
            reg_file[21851] <= 8'h00;
            reg_file[21852] <= 8'h00;
            reg_file[21853] <= 8'h00;
            reg_file[21854] <= 8'h00;
            reg_file[21855] <= 8'h00;
            reg_file[21856] <= 8'h00;
            reg_file[21857] <= 8'h00;
            reg_file[21858] <= 8'h00;
            reg_file[21859] <= 8'h00;
            reg_file[21860] <= 8'h00;
            reg_file[21861] <= 8'h00;
            reg_file[21862] <= 8'h00;
            reg_file[21863] <= 8'h00;
            reg_file[21864] <= 8'h00;
            reg_file[21865] <= 8'h00;
            reg_file[21866] <= 8'h00;
            reg_file[21867] <= 8'h00;
            reg_file[21868] <= 8'h00;
            reg_file[21869] <= 8'h00;
            reg_file[21870] <= 8'h00;
            reg_file[21871] <= 8'h00;
            reg_file[21872] <= 8'h00;
            reg_file[21873] <= 8'h00;
            reg_file[21874] <= 8'h00;
            reg_file[21875] <= 8'h00;
            reg_file[21876] <= 8'h00;
            reg_file[21877] <= 8'h00;
            reg_file[21878] <= 8'h00;
            reg_file[21879] <= 8'h00;
            reg_file[21880] <= 8'h00;
            reg_file[21881] <= 8'h00;
            reg_file[21882] <= 8'h00;
            reg_file[21883] <= 8'h00;
            reg_file[21884] <= 8'h00;
            reg_file[21885] <= 8'h00;
            reg_file[21886] <= 8'h00;
            reg_file[21887] <= 8'h00;
            reg_file[21888] <= 8'h00;
            reg_file[21889] <= 8'h00;
            reg_file[21890] <= 8'h00;
            reg_file[21891] <= 8'h00;
            reg_file[21892] <= 8'h00;
            reg_file[21893] <= 8'h00;
            reg_file[21894] <= 8'h00;
            reg_file[21895] <= 8'h00;
            reg_file[21896] <= 8'h00;
            reg_file[21897] <= 8'h00;
            reg_file[21898] <= 8'h00;
            reg_file[21899] <= 8'h00;
            reg_file[21900] <= 8'h00;
            reg_file[21901] <= 8'h00;
            reg_file[21902] <= 8'h00;
            reg_file[21903] <= 8'h00;
            reg_file[21904] <= 8'h00;
            reg_file[21905] <= 8'h00;
            reg_file[21906] <= 8'h00;
            reg_file[21907] <= 8'h00;
            reg_file[21908] <= 8'h00;
            reg_file[21909] <= 8'h00;
            reg_file[21910] <= 8'h00;
            reg_file[21911] <= 8'h00;
            reg_file[21912] <= 8'h00;
            reg_file[21913] <= 8'h00;
            reg_file[21914] <= 8'h00;
            reg_file[21915] <= 8'h00;
            reg_file[21916] <= 8'h00;
            reg_file[21917] <= 8'h00;
            reg_file[21918] <= 8'h00;
            reg_file[21919] <= 8'h00;
            reg_file[21920] <= 8'h00;
            reg_file[21921] <= 8'h00;
            reg_file[21922] <= 8'h00;
            reg_file[21923] <= 8'h00;
            reg_file[21924] <= 8'h00;
            reg_file[21925] <= 8'h00;
            reg_file[21926] <= 8'h00;
            reg_file[21927] <= 8'h00;
            reg_file[21928] <= 8'h00;
            reg_file[21929] <= 8'h00;
            reg_file[21930] <= 8'h00;
            reg_file[21931] <= 8'h00;
            reg_file[21932] <= 8'h00;
            reg_file[21933] <= 8'h00;
            reg_file[21934] <= 8'h00;
            reg_file[21935] <= 8'h00;
            reg_file[21936] <= 8'h00;
            reg_file[21937] <= 8'h00;
            reg_file[21938] <= 8'h00;
            reg_file[21939] <= 8'h00;
            reg_file[21940] <= 8'h00;
            reg_file[21941] <= 8'h00;
            reg_file[21942] <= 8'h00;
            reg_file[21943] <= 8'h00;
            reg_file[21944] <= 8'h00;
            reg_file[21945] <= 8'h00;
            reg_file[21946] <= 8'h00;
            reg_file[21947] <= 8'h00;
            reg_file[21948] <= 8'h00;
            reg_file[21949] <= 8'h00;
            reg_file[21950] <= 8'h00;
            reg_file[21951] <= 8'h00;
            reg_file[21952] <= 8'h00;
            reg_file[21953] <= 8'h00;
            reg_file[21954] <= 8'h00;
            reg_file[21955] <= 8'h00;
            reg_file[21956] <= 8'h00;
            reg_file[21957] <= 8'h00;
            reg_file[21958] <= 8'h00;
            reg_file[21959] <= 8'h00;
            reg_file[21960] <= 8'h00;
            reg_file[21961] <= 8'h00;
            reg_file[21962] <= 8'h00;
            reg_file[21963] <= 8'h00;
            reg_file[21964] <= 8'h00;
            reg_file[21965] <= 8'h00;
            reg_file[21966] <= 8'h00;
            reg_file[21967] <= 8'h00;
            reg_file[21968] <= 8'h00;
            reg_file[21969] <= 8'h00;
            reg_file[21970] <= 8'h00;
            reg_file[21971] <= 8'h00;
            reg_file[21972] <= 8'h00;
            reg_file[21973] <= 8'h00;
            reg_file[21974] <= 8'h00;
            reg_file[21975] <= 8'h00;
            reg_file[21976] <= 8'h00;
            reg_file[21977] <= 8'h00;
            reg_file[21978] <= 8'h00;
            reg_file[21979] <= 8'h00;
            reg_file[21980] <= 8'h00;
            reg_file[21981] <= 8'h00;
            reg_file[21982] <= 8'h00;
            reg_file[21983] <= 8'h00;
            reg_file[21984] <= 8'h00;
            reg_file[21985] <= 8'h00;
            reg_file[21986] <= 8'h00;
            reg_file[21987] <= 8'h00;
            reg_file[21988] <= 8'h00;
            reg_file[21989] <= 8'h00;
            reg_file[21990] <= 8'h00;
            reg_file[21991] <= 8'h00;
            reg_file[21992] <= 8'h00;
            reg_file[21993] <= 8'h00;
            reg_file[21994] <= 8'h00;
            reg_file[21995] <= 8'h00;
            reg_file[21996] <= 8'h00;
            reg_file[21997] <= 8'h00;
            reg_file[21998] <= 8'h00;
            reg_file[21999] <= 8'h00;
            reg_file[22000] <= 8'h00;
            reg_file[22001] <= 8'h00;
            reg_file[22002] <= 8'h00;
            reg_file[22003] <= 8'h00;
            reg_file[22004] <= 8'h00;
            reg_file[22005] <= 8'h00;
            reg_file[22006] <= 8'h00;
            reg_file[22007] <= 8'h00;
            reg_file[22008] <= 8'h00;
            reg_file[22009] <= 8'h00;
            reg_file[22010] <= 8'h00;
            reg_file[22011] <= 8'h00;
            reg_file[22012] <= 8'h00;
            reg_file[22013] <= 8'h00;
            reg_file[22014] <= 8'h00;
            reg_file[22015] <= 8'h00;
            reg_file[22016] <= 8'h00;
            reg_file[22017] <= 8'h00;
            reg_file[22018] <= 8'h00;
            reg_file[22019] <= 8'h00;
            reg_file[22020] <= 8'h00;
            reg_file[22021] <= 8'h00;
            reg_file[22022] <= 8'h00;
            reg_file[22023] <= 8'h00;
            reg_file[22024] <= 8'h00;
            reg_file[22025] <= 8'h00;
            reg_file[22026] <= 8'h00;
            reg_file[22027] <= 8'h00;
            reg_file[22028] <= 8'h00;
            reg_file[22029] <= 8'h00;
            reg_file[22030] <= 8'h00;
            reg_file[22031] <= 8'h00;
            reg_file[22032] <= 8'h00;
            reg_file[22033] <= 8'h00;
            reg_file[22034] <= 8'h00;
            reg_file[22035] <= 8'h00;
            reg_file[22036] <= 8'h00;
            reg_file[22037] <= 8'h00;
            reg_file[22038] <= 8'h00;
            reg_file[22039] <= 8'h00;
            reg_file[22040] <= 8'h00;
            reg_file[22041] <= 8'h00;
            reg_file[22042] <= 8'h00;
            reg_file[22043] <= 8'h00;
            reg_file[22044] <= 8'h00;
            reg_file[22045] <= 8'h00;
            reg_file[22046] <= 8'h00;
            reg_file[22047] <= 8'h00;
            reg_file[22048] <= 8'h00;
            reg_file[22049] <= 8'h00;
            reg_file[22050] <= 8'h00;
            reg_file[22051] <= 8'h00;
            reg_file[22052] <= 8'h00;
            reg_file[22053] <= 8'h00;
            reg_file[22054] <= 8'h00;
            reg_file[22055] <= 8'h00;
            reg_file[22056] <= 8'h00;
            reg_file[22057] <= 8'h00;
            reg_file[22058] <= 8'h00;
            reg_file[22059] <= 8'h00;
            reg_file[22060] <= 8'h00;
            reg_file[22061] <= 8'h00;
            reg_file[22062] <= 8'h00;
            reg_file[22063] <= 8'h00;
            reg_file[22064] <= 8'h00;
            reg_file[22065] <= 8'h00;
            reg_file[22066] <= 8'h00;
            reg_file[22067] <= 8'h00;
            reg_file[22068] <= 8'h00;
            reg_file[22069] <= 8'h00;
            reg_file[22070] <= 8'h00;
            reg_file[22071] <= 8'h00;
            reg_file[22072] <= 8'h00;
            reg_file[22073] <= 8'h00;
            reg_file[22074] <= 8'h00;
            reg_file[22075] <= 8'h00;
            reg_file[22076] <= 8'h00;
            reg_file[22077] <= 8'h00;
            reg_file[22078] <= 8'h00;
            reg_file[22079] <= 8'h00;
            reg_file[22080] <= 8'h00;
            reg_file[22081] <= 8'h00;
            reg_file[22082] <= 8'h00;
            reg_file[22083] <= 8'h00;
            reg_file[22084] <= 8'h00;
            reg_file[22085] <= 8'h00;
            reg_file[22086] <= 8'h00;
            reg_file[22087] <= 8'h00;
            reg_file[22088] <= 8'h00;
            reg_file[22089] <= 8'h00;
            reg_file[22090] <= 8'h00;
            reg_file[22091] <= 8'h00;
            reg_file[22092] <= 8'h00;
            reg_file[22093] <= 8'h00;
            reg_file[22094] <= 8'h00;
            reg_file[22095] <= 8'h00;
            reg_file[22096] <= 8'h00;
            reg_file[22097] <= 8'h00;
            reg_file[22098] <= 8'h00;
            reg_file[22099] <= 8'h00;
            reg_file[22100] <= 8'h00;
            reg_file[22101] <= 8'h00;
            reg_file[22102] <= 8'h00;
            reg_file[22103] <= 8'h00;
            reg_file[22104] <= 8'h00;
            reg_file[22105] <= 8'h00;
            reg_file[22106] <= 8'h00;
            reg_file[22107] <= 8'h00;
            reg_file[22108] <= 8'h00;
            reg_file[22109] <= 8'h00;
            reg_file[22110] <= 8'h00;
            reg_file[22111] <= 8'h00;
            reg_file[22112] <= 8'h00;
            reg_file[22113] <= 8'h00;
            reg_file[22114] <= 8'h00;
            reg_file[22115] <= 8'h00;
            reg_file[22116] <= 8'h00;
            reg_file[22117] <= 8'h00;
            reg_file[22118] <= 8'h00;
            reg_file[22119] <= 8'h00;
            reg_file[22120] <= 8'h00;
            reg_file[22121] <= 8'h00;
            reg_file[22122] <= 8'h00;
            reg_file[22123] <= 8'h00;
            reg_file[22124] <= 8'h00;
            reg_file[22125] <= 8'h00;
            reg_file[22126] <= 8'h00;
            reg_file[22127] <= 8'h00;
            reg_file[22128] <= 8'h00;
            reg_file[22129] <= 8'h00;
            reg_file[22130] <= 8'h00;
            reg_file[22131] <= 8'h00;
            reg_file[22132] <= 8'h00;
            reg_file[22133] <= 8'h00;
            reg_file[22134] <= 8'h00;
            reg_file[22135] <= 8'h00;
            reg_file[22136] <= 8'h00;
            reg_file[22137] <= 8'h00;
            reg_file[22138] <= 8'h00;
            reg_file[22139] <= 8'h00;
            reg_file[22140] <= 8'h00;
            reg_file[22141] <= 8'h00;
            reg_file[22142] <= 8'h00;
            reg_file[22143] <= 8'h00;
            reg_file[22144] <= 8'h00;
            reg_file[22145] <= 8'h00;
            reg_file[22146] <= 8'h00;
            reg_file[22147] <= 8'h00;
            reg_file[22148] <= 8'h00;
            reg_file[22149] <= 8'h00;
            reg_file[22150] <= 8'h00;
            reg_file[22151] <= 8'h00;
            reg_file[22152] <= 8'h00;
            reg_file[22153] <= 8'h00;
            reg_file[22154] <= 8'h00;
            reg_file[22155] <= 8'h00;
            reg_file[22156] <= 8'h00;
            reg_file[22157] <= 8'h00;
            reg_file[22158] <= 8'h00;
            reg_file[22159] <= 8'h00;
            reg_file[22160] <= 8'h00;
            reg_file[22161] <= 8'h00;
            reg_file[22162] <= 8'h00;
            reg_file[22163] <= 8'h00;
            reg_file[22164] <= 8'h00;
            reg_file[22165] <= 8'h00;
            reg_file[22166] <= 8'h00;
            reg_file[22167] <= 8'h00;
            reg_file[22168] <= 8'h00;
            reg_file[22169] <= 8'h00;
            reg_file[22170] <= 8'h00;
            reg_file[22171] <= 8'h00;
            reg_file[22172] <= 8'h00;
            reg_file[22173] <= 8'h00;
            reg_file[22174] <= 8'h00;
            reg_file[22175] <= 8'h00;
            reg_file[22176] <= 8'h00;
            reg_file[22177] <= 8'h00;
            reg_file[22178] <= 8'h00;
            reg_file[22179] <= 8'h00;
            reg_file[22180] <= 8'h00;
            reg_file[22181] <= 8'h00;
            reg_file[22182] <= 8'h00;
            reg_file[22183] <= 8'h00;
            reg_file[22184] <= 8'h00;
            reg_file[22185] <= 8'h00;
            reg_file[22186] <= 8'h00;
            reg_file[22187] <= 8'h00;
            reg_file[22188] <= 8'h00;
            reg_file[22189] <= 8'h00;
            reg_file[22190] <= 8'h00;
            reg_file[22191] <= 8'h00;
            reg_file[22192] <= 8'h00;
            reg_file[22193] <= 8'h00;
            reg_file[22194] <= 8'h00;
            reg_file[22195] <= 8'h00;
            reg_file[22196] <= 8'h00;
            reg_file[22197] <= 8'h00;
            reg_file[22198] <= 8'h00;
            reg_file[22199] <= 8'h00;
            reg_file[22200] <= 8'h00;
            reg_file[22201] <= 8'h00;
            reg_file[22202] <= 8'h00;
            reg_file[22203] <= 8'h00;
            reg_file[22204] <= 8'h00;
            reg_file[22205] <= 8'h00;
            reg_file[22206] <= 8'h00;
            reg_file[22207] <= 8'h00;
            reg_file[22208] <= 8'h00;
            reg_file[22209] <= 8'h00;
            reg_file[22210] <= 8'h00;
            reg_file[22211] <= 8'h00;
            reg_file[22212] <= 8'h00;
            reg_file[22213] <= 8'h00;
            reg_file[22214] <= 8'h00;
            reg_file[22215] <= 8'h00;
            reg_file[22216] <= 8'h00;
            reg_file[22217] <= 8'h00;
            reg_file[22218] <= 8'h00;
            reg_file[22219] <= 8'h00;
            reg_file[22220] <= 8'h00;
            reg_file[22221] <= 8'h00;
            reg_file[22222] <= 8'h00;
            reg_file[22223] <= 8'h00;
            reg_file[22224] <= 8'h00;
            reg_file[22225] <= 8'h00;
            reg_file[22226] <= 8'h00;
            reg_file[22227] <= 8'h00;
            reg_file[22228] <= 8'h00;
            reg_file[22229] <= 8'h00;
            reg_file[22230] <= 8'h00;
            reg_file[22231] <= 8'h00;
            reg_file[22232] <= 8'h00;
            reg_file[22233] <= 8'h00;
            reg_file[22234] <= 8'h00;
            reg_file[22235] <= 8'h00;
            reg_file[22236] <= 8'h00;
            reg_file[22237] <= 8'h00;
            reg_file[22238] <= 8'h00;
            reg_file[22239] <= 8'h00;
            reg_file[22240] <= 8'h00;
            reg_file[22241] <= 8'h00;
            reg_file[22242] <= 8'h00;
            reg_file[22243] <= 8'h00;
            reg_file[22244] <= 8'h00;
            reg_file[22245] <= 8'h00;
            reg_file[22246] <= 8'h00;
            reg_file[22247] <= 8'h00;
            reg_file[22248] <= 8'h00;
            reg_file[22249] <= 8'h00;
            reg_file[22250] <= 8'h00;
            reg_file[22251] <= 8'h00;
            reg_file[22252] <= 8'h00;
            reg_file[22253] <= 8'h00;
            reg_file[22254] <= 8'h00;
            reg_file[22255] <= 8'h00;
            reg_file[22256] <= 8'h00;
            reg_file[22257] <= 8'h00;
            reg_file[22258] <= 8'h00;
            reg_file[22259] <= 8'h00;
            reg_file[22260] <= 8'h00;
            reg_file[22261] <= 8'h00;
            reg_file[22262] <= 8'h00;
            reg_file[22263] <= 8'h00;
            reg_file[22264] <= 8'h00;
            reg_file[22265] <= 8'h00;
            reg_file[22266] <= 8'h00;
            reg_file[22267] <= 8'h00;
            reg_file[22268] <= 8'h00;
            reg_file[22269] <= 8'h00;
            reg_file[22270] <= 8'h00;
            reg_file[22271] <= 8'h00;
            reg_file[22272] <= 8'h00;
            reg_file[22273] <= 8'h00;
            reg_file[22274] <= 8'h00;
            reg_file[22275] <= 8'h00;
            reg_file[22276] <= 8'h00;
            reg_file[22277] <= 8'h00;
            reg_file[22278] <= 8'h00;
            reg_file[22279] <= 8'h00;
            reg_file[22280] <= 8'h00;
            reg_file[22281] <= 8'h00;
            reg_file[22282] <= 8'h00;
            reg_file[22283] <= 8'h00;
            reg_file[22284] <= 8'h00;
            reg_file[22285] <= 8'h00;
            reg_file[22286] <= 8'h00;
            reg_file[22287] <= 8'h00;
            reg_file[22288] <= 8'h00;
            reg_file[22289] <= 8'h00;
            reg_file[22290] <= 8'h00;
            reg_file[22291] <= 8'h00;
            reg_file[22292] <= 8'h00;
            reg_file[22293] <= 8'h00;
            reg_file[22294] <= 8'h00;
            reg_file[22295] <= 8'h00;
            reg_file[22296] <= 8'h00;
            reg_file[22297] <= 8'h00;
            reg_file[22298] <= 8'h00;
            reg_file[22299] <= 8'h00;
            reg_file[22300] <= 8'h00;
            reg_file[22301] <= 8'h00;
            reg_file[22302] <= 8'h00;
            reg_file[22303] <= 8'h00;
            reg_file[22304] <= 8'h00;
            reg_file[22305] <= 8'h00;
            reg_file[22306] <= 8'h00;
            reg_file[22307] <= 8'h00;
            reg_file[22308] <= 8'h00;
            reg_file[22309] <= 8'h00;
            reg_file[22310] <= 8'h00;
            reg_file[22311] <= 8'h00;
            reg_file[22312] <= 8'h00;
            reg_file[22313] <= 8'h00;
            reg_file[22314] <= 8'h00;
            reg_file[22315] <= 8'h00;
            reg_file[22316] <= 8'h00;
            reg_file[22317] <= 8'h00;
            reg_file[22318] <= 8'h00;
            reg_file[22319] <= 8'h00;
            reg_file[22320] <= 8'h00;
            reg_file[22321] <= 8'h00;
            reg_file[22322] <= 8'h00;
            reg_file[22323] <= 8'h00;
            reg_file[22324] <= 8'h00;
            reg_file[22325] <= 8'h00;
            reg_file[22326] <= 8'h00;
            reg_file[22327] <= 8'h00;
            reg_file[22328] <= 8'h00;
            reg_file[22329] <= 8'h00;
            reg_file[22330] <= 8'h00;
            reg_file[22331] <= 8'h00;
            reg_file[22332] <= 8'h00;
            reg_file[22333] <= 8'h00;
            reg_file[22334] <= 8'h00;
            reg_file[22335] <= 8'h00;
            reg_file[22336] <= 8'h00;
            reg_file[22337] <= 8'h00;
            reg_file[22338] <= 8'h00;
            reg_file[22339] <= 8'h00;
            reg_file[22340] <= 8'h00;
            reg_file[22341] <= 8'h00;
            reg_file[22342] <= 8'h00;
            reg_file[22343] <= 8'h00;
            reg_file[22344] <= 8'h00;
            reg_file[22345] <= 8'h00;
            reg_file[22346] <= 8'h00;
            reg_file[22347] <= 8'h00;
            reg_file[22348] <= 8'h00;
            reg_file[22349] <= 8'h00;
            reg_file[22350] <= 8'h00;
            reg_file[22351] <= 8'h00;
            reg_file[22352] <= 8'h00;
            reg_file[22353] <= 8'h00;
            reg_file[22354] <= 8'h00;
            reg_file[22355] <= 8'h00;
            reg_file[22356] <= 8'h00;
            reg_file[22357] <= 8'h00;
            reg_file[22358] <= 8'h00;
            reg_file[22359] <= 8'h00;
            reg_file[22360] <= 8'h00;
            reg_file[22361] <= 8'h00;
            reg_file[22362] <= 8'h00;
            reg_file[22363] <= 8'h00;
            reg_file[22364] <= 8'h00;
            reg_file[22365] <= 8'h00;
            reg_file[22366] <= 8'h00;
            reg_file[22367] <= 8'h00;
            reg_file[22368] <= 8'h00;
            reg_file[22369] <= 8'h00;
            reg_file[22370] <= 8'h00;
            reg_file[22371] <= 8'h00;
            reg_file[22372] <= 8'h00;
            reg_file[22373] <= 8'h00;
            reg_file[22374] <= 8'h00;
            reg_file[22375] <= 8'h00;
            reg_file[22376] <= 8'h00;
            reg_file[22377] <= 8'h00;
            reg_file[22378] <= 8'h00;
            reg_file[22379] <= 8'h00;
            reg_file[22380] <= 8'h00;
            reg_file[22381] <= 8'h00;
            reg_file[22382] <= 8'h00;
            reg_file[22383] <= 8'h00;
            reg_file[22384] <= 8'h00;
            reg_file[22385] <= 8'h00;
            reg_file[22386] <= 8'h00;
            reg_file[22387] <= 8'h00;
            reg_file[22388] <= 8'h00;
            reg_file[22389] <= 8'h00;
            reg_file[22390] <= 8'h00;
            reg_file[22391] <= 8'h00;
            reg_file[22392] <= 8'h00;
            reg_file[22393] <= 8'h00;
            reg_file[22394] <= 8'h00;
            reg_file[22395] <= 8'h00;
            reg_file[22396] <= 8'h00;
            reg_file[22397] <= 8'h00;
            reg_file[22398] <= 8'h00;
            reg_file[22399] <= 8'h00;
            reg_file[22400] <= 8'h00;
            reg_file[22401] <= 8'h00;
            reg_file[22402] <= 8'h00;
            reg_file[22403] <= 8'h00;
            reg_file[22404] <= 8'h00;
            reg_file[22405] <= 8'h00;
            reg_file[22406] <= 8'h00;
            reg_file[22407] <= 8'h00;
            reg_file[22408] <= 8'h00;
            reg_file[22409] <= 8'h00;
            reg_file[22410] <= 8'h00;
            reg_file[22411] <= 8'h00;
            reg_file[22412] <= 8'h00;
            reg_file[22413] <= 8'h00;
            reg_file[22414] <= 8'h00;
            reg_file[22415] <= 8'h00;
            reg_file[22416] <= 8'h00;
            reg_file[22417] <= 8'h00;
            reg_file[22418] <= 8'h00;
            reg_file[22419] <= 8'h00;
            reg_file[22420] <= 8'h00;
            reg_file[22421] <= 8'h00;
            reg_file[22422] <= 8'h00;
            reg_file[22423] <= 8'h00;
            reg_file[22424] <= 8'h00;
            reg_file[22425] <= 8'h00;
            reg_file[22426] <= 8'h00;
            reg_file[22427] <= 8'h00;
            reg_file[22428] <= 8'h00;
            reg_file[22429] <= 8'h00;
            reg_file[22430] <= 8'h00;
            reg_file[22431] <= 8'h00;
            reg_file[22432] <= 8'h00;
            reg_file[22433] <= 8'h00;
            reg_file[22434] <= 8'h00;
            reg_file[22435] <= 8'h00;
            reg_file[22436] <= 8'h00;
            reg_file[22437] <= 8'h00;
            reg_file[22438] <= 8'h00;
            reg_file[22439] <= 8'h00;
            reg_file[22440] <= 8'h00;
            reg_file[22441] <= 8'h00;
            reg_file[22442] <= 8'h00;
            reg_file[22443] <= 8'h00;
            reg_file[22444] <= 8'h00;
            reg_file[22445] <= 8'h00;
            reg_file[22446] <= 8'h00;
            reg_file[22447] <= 8'h00;
            reg_file[22448] <= 8'h00;
            reg_file[22449] <= 8'h00;
            reg_file[22450] <= 8'h00;
            reg_file[22451] <= 8'h00;
            reg_file[22452] <= 8'h00;
            reg_file[22453] <= 8'h00;
            reg_file[22454] <= 8'h00;
            reg_file[22455] <= 8'h00;
            reg_file[22456] <= 8'h00;
            reg_file[22457] <= 8'h00;
            reg_file[22458] <= 8'h00;
            reg_file[22459] <= 8'h00;
            reg_file[22460] <= 8'h00;
            reg_file[22461] <= 8'h00;
            reg_file[22462] <= 8'h00;
            reg_file[22463] <= 8'h00;
            reg_file[22464] <= 8'h00;
            reg_file[22465] <= 8'h00;
            reg_file[22466] <= 8'h00;
            reg_file[22467] <= 8'h00;
            reg_file[22468] <= 8'h00;
            reg_file[22469] <= 8'h00;
            reg_file[22470] <= 8'h00;
            reg_file[22471] <= 8'h00;
            reg_file[22472] <= 8'h00;
            reg_file[22473] <= 8'h00;
            reg_file[22474] <= 8'h00;
            reg_file[22475] <= 8'h00;
            reg_file[22476] <= 8'h00;
            reg_file[22477] <= 8'h00;
            reg_file[22478] <= 8'h00;
            reg_file[22479] <= 8'h00;
            reg_file[22480] <= 8'h00;
            reg_file[22481] <= 8'h00;
            reg_file[22482] <= 8'h00;
            reg_file[22483] <= 8'h00;
            reg_file[22484] <= 8'h00;
            reg_file[22485] <= 8'h00;
            reg_file[22486] <= 8'h00;
            reg_file[22487] <= 8'h00;
            reg_file[22488] <= 8'h00;
            reg_file[22489] <= 8'h00;
            reg_file[22490] <= 8'h00;
            reg_file[22491] <= 8'h00;
            reg_file[22492] <= 8'h00;
            reg_file[22493] <= 8'h00;
            reg_file[22494] <= 8'h00;
            reg_file[22495] <= 8'h00;
            reg_file[22496] <= 8'h00;
            reg_file[22497] <= 8'h00;
            reg_file[22498] <= 8'h00;
            reg_file[22499] <= 8'h00;
            reg_file[22500] <= 8'h00;
            reg_file[22501] <= 8'h00;
            reg_file[22502] <= 8'h00;
            reg_file[22503] <= 8'h00;
            reg_file[22504] <= 8'h00;
            reg_file[22505] <= 8'h00;
            reg_file[22506] <= 8'h00;
            reg_file[22507] <= 8'h00;
            reg_file[22508] <= 8'h00;
            reg_file[22509] <= 8'h00;
            reg_file[22510] <= 8'h00;
            reg_file[22511] <= 8'h00;
            reg_file[22512] <= 8'h00;
            reg_file[22513] <= 8'h00;
            reg_file[22514] <= 8'h00;
            reg_file[22515] <= 8'h00;
            reg_file[22516] <= 8'h00;
            reg_file[22517] <= 8'h00;
            reg_file[22518] <= 8'h00;
            reg_file[22519] <= 8'h00;
            reg_file[22520] <= 8'h00;
            reg_file[22521] <= 8'h00;
            reg_file[22522] <= 8'h00;
            reg_file[22523] <= 8'h00;
            reg_file[22524] <= 8'h00;
            reg_file[22525] <= 8'h00;
            reg_file[22526] <= 8'h00;
            reg_file[22527] <= 8'h00;
            reg_file[22528] <= 8'h00;
            reg_file[22529] <= 8'h00;
            reg_file[22530] <= 8'h00;
            reg_file[22531] <= 8'h00;
            reg_file[22532] <= 8'h00;
            reg_file[22533] <= 8'h00;
            reg_file[22534] <= 8'h00;
            reg_file[22535] <= 8'h00;
            reg_file[22536] <= 8'h00;
            reg_file[22537] <= 8'h00;
            reg_file[22538] <= 8'h00;
            reg_file[22539] <= 8'h00;
            reg_file[22540] <= 8'h00;
            reg_file[22541] <= 8'h00;
            reg_file[22542] <= 8'h00;
            reg_file[22543] <= 8'h00;
            reg_file[22544] <= 8'h00;
            reg_file[22545] <= 8'h00;
            reg_file[22546] <= 8'h00;
            reg_file[22547] <= 8'h00;
            reg_file[22548] <= 8'h00;
            reg_file[22549] <= 8'h00;
            reg_file[22550] <= 8'h00;
            reg_file[22551] <= 8'h00;
            reg_file[22552] <= 8'h00;
            reg_file[22553] <= 8'h00;
            reg_file[22554] <= 8'h00;
            reg_file[22555] <= 8'h00;
            reg_file[22556] <= 8'h00;
            reg_file[22557] <= 8'h00;
            reg_file[22558] <= 8'h00;
            reg_file[22559] <= 8'h00;
            reg_file[22560] <= 8'h00;
            reg_file[22561] <= 8'h00;
            reg_file[22562] <= 8'h00;
            reg_file[22563] <= 8'h00;
            reg_file[22564] <= 8'h00;
            reg_file[22565] <= 8'h00;
            reg_file[22566] <= 8'h00;
            reg_file[22567] <= 8'h00;
            reg_file[22568] <= 8'h00;
            reg_file[22569] <= 8'h00;
            reg_file[22570] <= 8'h00;
            reg_file[22571] <= 8'h00;
            reg_file[22572] <= 8'h00;
            reg_file[22573] <= 8'h00;
            reg_file[22574] <= 8'h00;
            reg_file[22575] <= 8'h00;
            reg_file[22576] <= 8'h00;
            reg_file[22577] <= 8'h00;
            reg_file[22578] <= 8'h00;
            reg_file[22579] <= 8'h00;
            reg_file[22580] <= 8'h00;
            reg_file[22581] <= 8'h00;
            reg_file[22582] <= 8'h00;
            reg_file[22583] <= 8'h00;
            reg_file[22584] <= 8'h00;
            reg_file[22585] <= 8'h00;
            reg_file[22586] <= 8'h00;
            reg_file[22587] <= 8'h00;
            reg_file[22588] <= 8'h00;
            reg_file[22589] <= 8'h00;
            reg_file[22590] <= 8'h00;
            reg_file[22591] <= 8'h00;
            reg_file[22592] <= 8'h00;
            reg_file[22593] <= 8'h00;
            reg_file[22594] <= 8'h00;
            reg_file[22595] <= 8'h00;
            reg_file[22596] <= 8'h00;
            reg_file[22597] <= 8'h00;
            reg_file[22598] <= 8'h00;
            reg_file[22599] <= 8'h00;
            reg_file[22600] <= 8'h00;
            reg_file[22601] <= 8'h00;
            reg_file[22602] <= 8'h00;
            reg_file[22603] <= 8'h00;
            reg_file[22604] <= 8'h00;
            reg_file[22605] <= 8'h00;
            reg_file[22606] <= 8'h00;
            reg_file[22607] <= 8'h00;
            reg_file[22608] <= 8'h00;
            reg_file[22609] <= 8'h00;
            reg_file[22610] <= 8'h00;
            reg_file[22611] <= 8'h00;
            reg_file[22612] <= 8'h00;
            reg_file[22613] <= 8'h00;
            reg_file[22614] <= 8'h00;
            reg_file[22615] <= 8'h00;
            reg_file[22616] <= 8'h00;
            reg_file[22617] <= 8'h00;
            reg_file[22618] <= 8'h00;
            reg_file[22619] <= 8'h00;
            reg_file[22620] <= 8'h00;
            reg_file[22621] <= 8'h00;
            reg_file[22622] <= 8'h00;
            reg_file[22623] <= 8'h00;
            reg_file[22624] <= 8'h00;
            reg_file[22625] <= 8'h00;
            reg_file[22626] <= 8'h00;
            reg_file[22627] <= 8'h00;
            reg_file[22628] <= 8'h00;
            reg_file[22629] <= 8'h00;
            reg_file[22630] <= 8'h00;
            reg_file[22631] <= 8'h00;
            reg_file[22632] <= 8'h00;
            reg_file[22633] <= 8'h00;
            reg_file[22634] <= 8'h00;
            reg_file[22635] <= 8'h00;
            reg_file[22636] <= 8'h00;
            reg_file[22637] <= 8'h00;
            reg_file[22638] <= 8'h00;
            reg_file[22639] <= 8'h00;
            reg_file[22640] <= 8'h00;
            reg_file[22641] <= 8'h00;
            reg_file[22642] <= 8'h00;
            reg_file[22643] <= 8'h00;
            reg_file[22644] <= 8'h00;
            reg_file[22645] <= 8'h00;
            reg_file[22646] <= 8'h00;
            reg_file[22647] <= 8'h00;
            reg_file[22648] <= 8'h00;
            reg_file[22649] <= 8'h00;
            reg_file[22650] <= 8'h00;
            reg_file[22651] <= 8'h00;
            reg_file[22652] <= 8'h00;
            reg_file[22653] <= 8'h00;
            reg_file[22654] <= 8'h00;
            reg_file[22655] <= 8'h00;
            reg_file[22656] <= 8'h00;
            reg_file[22657] <= 8'h00;
            reg_file[22658] <= 8'h00;
            reg_file[22659] <= 8'h00;
            reg_file[22660] <= 8'h00;
            reg_file[22661] <= 8'h00;
            reg_file[22662] <= 8'h00;
            reg_file[22663] <= 8'h00;
            reg_file[22664] <= 8'h00;
            reg_file[22665] <= 8'h00;
            reg_file[22666] <= 8'h00;
            reg_file[22667] <= 8'h00;
            reg_file[22668] <= 8'h00;
            reg_file[22669] <= 8'h00;
            reg_file[22670] <= 8'h00;
            reg_file[22671] <= 8'h00;
            reg_file[22672] <= 8'h00;
            reg_file[22673] <= 8'h00;
            reg_file[22674] <= 8'h00;
            reg_file[22675] <= 8'h00;
            reg_file[22676] <= 8'h00;
            reg_file[22677] <= 8'h00;
            reg_file[22678] <= 8'h00;
            reg_file[22679] <= 8'h00;
            reg_file[22680] <= 8'h00;
            reg_file[22681] <= 8'h00;
            reg_file[22682] <= 8'h00;
            reg_file[22683] <= 8'h00;
            reg_file[22684] <= 8'h00;
            reg_file[22685] <= 8'h00;
            reg_file[22686] <= 8'h00;
            reg_file[22687] <= 8'h00;
            reg_file[22688] <= 8'h00;
            reg_file[22689] <= 8'h00;
            reg_file[22690] <= 8'h00;
            reg_file[22691] <= 8'h00;
            reg_file[22692] <= 8'h00;
            reg_file[22693] <= 8'h00;
            reg_file[22694] <= 8'h00;
            reg_file[22695] <= 8'h00;
            reg_file[22696] <= 8'h00;
            reg_file[22697] <= 8'h00;
            reg_file[22698] <= 8'h00;
            reg_file[22699] <= 8'h00;
            reg_file[22700] <= 8'h00;
            reg_file[22701] <= 8'h00;
            reg_file[22702] <= 8'h00;
            reg_file[22703] <= 8'h00;
            reg_file[22704] <= 8'h00;
            reg_file[22705] <= 8'h00;
            reg_file[22706] <= 8'h00;
            reg_file[22707] <= 8'h00;
            reg_file[22708] <= 8'h00;
            reg_file[22709] <= 8'h00;
            reg_file[22710] <= 8'h00;
            reg_file[22711] <= 8'h00;
            reg_file[22712] <= 8'h00;
            reg_file[22713] <= 8'h00;
            reg_file[22714] <= 8'h00;
            reg_file[22715] <= 8'h00;
            reg_file[22716] <= 8'h00;
            reg_file[22717] <= 8'h00;
            reg_file[22718] <= 8'h00;
            reg_file[22719] <= 8'h00;
            reg_file[22720] <= 8'h00;
            reg_file[22721] <= 8'h00;
            reg_file[22722] <= 8'h00;
            reg_file[22723] <= 8'h00;
            reg_file[22724] <= 8'h00;
            reg_file[22725] <= 8'h00;
            reg_file[22726] <= 8'h00;
            reg_file[22727] <= 8'h00;
            reg_file[22728] <= 8'h00;
            reg_file[22729] <= 8'h00;
            reg_file[22730] <= 8'h00;
            reg_file[22731] <= 8'h00;
            reg_file[22732] <= 8'h00;
            reg_file[22733] <= 8'h00;
            reg_file[22734] <= 8'h00;
            reg_file[22735] <= 8'h00;
            reg_file[22736] <= 8'h00;
            reg_file[22737] <= 8'h00;
            reg_file[22738] <= 8'h00;
            reg_file[22739] <= 8'h00;
            reg_file[22740] <= 8'h00;
            reg_file[22741] <= 8'h00;
            reg_file[22742] <= 8'h00;
            reg_file[22743] <= 8'h00;
            reg_file[22744] <= 8'h00;
            reg_file[22745] <= 8'h00;
            reg_file[22746] <= 8'h00;
            reg_file[22747] <= 8'h00;
            reg_file[22748] <= 8'h00;
            reg_file[22749] <= 8'h00;
            reg_file[22750] <= 8'h00;
            reg_file[22751] <= 8'h00;
            reg_file[22752] <= 8'h00;
            reg_file[22753] <= 8'h00;
            reg_file[22754] <= 8'h00;
            reg_file[22755] <= 8'h00;
            reg_file[22756] <= 8'h00;
            reg_file[22757] <= 8'h00;
            reg_file[22758] <= 8'h00;
            reg_file[22759] <= 8'h00;
            reg_file[22760] <= 8'h00;
            reg_file[22761] <= 8'h00;
            reg_file[22762] <= 8'h00;
            reg_file[22763] <= 8'h00;
            reg_file[22764] <= 8'h00;
            reg_file[22765] <= 8'h00;
            reg_file[22766] <= 8'h00;
            reg_file[22767] <= 8'h00;
            reg_file[22768] <= 8'h00;
            reg_file[22769] <= 8'h00;
            reg_file[22770] <= 8'h00;
            reg_file[22771] <= 8'h00;
            reg_file[22772] <= 8'h00;
            reg_file[22773] <= 8'h00;
            reg_file[22774] <= 8'h00;
            reg_file[22775] <= 8'h00;
            reg_file[22776] <= 8'h00;
            reg_file[22777] <= 8'h00;
            reg_file[22778] <= 8'h00;
            reg_file[22779] <= 8'h00;
            reg_file[22780] <= 8'h00;
            reg_file[22781] <= 8'h00;
            reg_file[22782] <= 8'h00;
            reg_file[22783] <= 8'h00;
            reg_file[22784] <= 8'h00;
            reg_file[22785] <= 8'h00;
            reg_file[22786] <= 8'h00;
            reg_file[22787] <= 8'h00;
            reg_file[22788] <= 8'h00;
            reg_file[22789] <= 8'h00;
            reg_file[22790] <= 8'h00;
            reg_file[22791] <= 8'h00;
            reg_file[22792] <= 8'h00;
            reg_file[22793] <= 8'h00;
            reg_file[22794] <= 8'h00;
            reg_file[22795] <= 8'h00;
            reg_file[22796] <= 8'h00;
            reg_file[22797] <= 8'h00;
            reg_file[22798] <= 8'h00;
            reg_file[22799] <= 8'h00;
            reg_file[22800] <= 8'h00;
            reg_file[22801] <= 8'h00;
            reg_file[22802] <= 8'h00;
            reg_file[22803] <= 8'h00;
            reg_file[22804] <= 8'h00;
            reg_file[22805] <= 8'h00;
            reg_file[22806] <= 8'h00;
            reg_file[22807] <= 8'h00;
            reg_file[22808] <= 8'h00;
            reg_file[22809] <= 8'h00;
            reg_file[22810] <= 8'h00;
            reg_file[22811] <= 8'h00;
            reg_file[22812] <= 8'h00;
            reg_file[22813] <= 8'h00;
            reg_file[22814] <= 8'h00;
            reg_file[22815] <= 8'h00;
            reg_file[22816] <= 8'h00;
            reg_file[22817] <= 8'h00;
            reg_file[22818] <= 8'h00;
            reg_file[22819] <= 8'h00;
            reg_file[22820] <= 8'h00;
            reg_file[22821] <= 8'h00;
            reg_file[22822] <= 8'h00;
            reg_file[22823] <= 8'h00;
            reg_file[22824] <= 8'h00;
            reg_file[22825] <= 8'h00;
            reg_file[22826] <= 8'h00;
            reg_file[22827] <= 8'h00;
            reg_file[22828] <= 8'h00;
            reg_file[22829] <= 8'h00;
            reg_file[22830] <= 8'h00;
            reg_file[22831] <= 8'h00;
            reg_file[22832] <= 8'h00;
            reg_file[22833] <= 8'h00;
            reg_file[22834] <= 8'h00;
            reg_file[22835] <= 8'h00;
            reg_file[22836] <= 8'h00;
            reg_file[22837] <= 8'h00;
            reg_file[22838] <= 8'h00;
            reg_file[22839] <= 8'h00;
            reg_file[22840] <= 8'h00;
            reg_file[22841] <= 8'h00;
            reg_file[22842] <= 8'h00;
            reg_file[22843] <= 8'h00;
            reg_file[22844] <= 8'h00;
            reg_file[22845] <= 8'h00;
            reg_file[22846] <= 8'h00;
            reg_file[22847] <= 8'h00;
            reg_file[22848] <= 8'h00;
            reg_file[22849] <= 8'h00;
            reg_file[22850] <= 8'h00;
            reg_file[22851] <= 8'h00;
            reg_file[22852] <= 8'h00;
            reg_file[22853] <= 8'h00;
            reg_file[22854] <= 8'h00;
            reg_file[22855] <= 8'h00;
            reg_file[22856] <= 8'h00;
            reg_file[22857] <= 8'h00;
            reg_file[22858] <= 8'h00;
            reg_file[22859] <= 8'h00;
            reg_file[22860] <= 8'h00;
            reg_file[22861] <= 8'h00;
            reg_file[22862] <= 8'h00;
            reg_file[22863] <= 8'h00;
            reg_file[22864] <= 8'h00;
            reg_file[22865] <= 8'h00;
            reg_file[22866] <= 8'h00;
            reg_file[22867] <= 8'h00;
            reg_file[22868] <= 8'h00;
            reg_file[22869] <= 8'h00;
            reg_file[22870] <= 8'h00;
            reg_file[22871] <= 8'h00;
            reg_file[22872] <= 8'h00;
            reg_file[22873] <= 8'h00;
            reg_file[22874] <= 8'h00;
            reg_file[22875] <= 8'h00;
            reg_file[22876] <= 8'h00;
            reg_file[22877] <= 8'h00;
            reg_file[22878] <= 8'h00;
            reg_file[22879] <= 8'h00;
            reg_file[22880] <= 8'h00;
            reg_file[22881] <= 8'h00;
            reg_file[22882] <= 8'h00;
            reg_file[22883] <= 8'h00;
            reg_file[22884] <= 8'h00;
            reg_file[22885] <= 8'h00;
            reg_file[22886] <= 8'h00;
            reg_file[22887] <= 8'h00;
            reg_file[22888] <= 8'h00;
            reg_file[22889] <= 8'h00;
            reg_file[22890] <= 8'h00;
            reg_file[22891] <= 8'h00;
            reg_file[22892] <= 8'h00;
            reg_file[22893] <= 8'h00;
            reg_file[22894] <= 8'h00;
            reg_file[22895] <= 8'h00;
            reg_file[22896] <= 8'h00;
            reg_file[22897] <= 8'h00;
            reg_file[22898] <= 8'h00;
            reg_file[22899] <= 8'h00;
            reg_file[22900] <= 8'h00;
            reg_file[22901] <= 8'h00;
            reg_file[22902] <= 8'h00;
            reg_file[22903] <= 8'h00;
            reg_file[22904] <= 8'h00;
            reg_file[22905] <= 8'h00;
            reg_file[22906] <= 8'h00;
            reg_file[22907] <= 8'h00;
            reg_file[22908] <= 8'h00;
            reg_file[22909] <= 8'h00;
            reg_file[22910] <= 8'h00;
            reg_file[22911] <= 8'h00;
            reg_file[22912] <= 8'h00;
            reg_file[22913] <= 8'h00;
            reg_file[22914] <= 8'h00;
            reg_file[22915] <= 8'h00;
            reg_file[22916] <= 8'h00;
            reg_file[22917] <= 8'h00;
            reg_file[22918] <= 8'h00;
            reg_file[22919] <= 8'h00;
            reg_file[22920] <= 8'h00;
            reg_file[22921] <= 8'h00;
            reg_file[22922] <= 8'h00;
            reg_file[22923] <= 8'h00;
            reg_file[22924] <= 8'h00;
            reg_file[22925] <= 8'h00;
            reg_file[22926] <= 8'h00;
            reg_file[22927] <= 8'h00;
            reg_file[22928] <= 8'h00;
            reg_file[22929] <= 8'h00;
            reg_file[22930] <= 8'h00;
            reg_file[22931] <= 8'h00;
            reg_file[22932] <= 8'h00;
            reg_file[22933] <= 8'h00;
            reg_file[22934] <= 8'h00;
            reg_file[22935] <= 8'h00;
            reg_file[22936] <= 8'h00;
            reg_file[22937] <= 8'h00;
            reg_file[22938] <= 8'h00;
            reg_file[22939] <= 8'h00;
            reg_file[22940] <= 8'h00;
            reg_file[22941] <= 8'h00;
            reg_file[22942] <= 8'h00;
            reg_file[22943] <= 8'h00;
            reg_file[22944] <= 8'h00;
            reg_file[22945] <= 8'h00;
            reg_file[22946] <= 8'h00;
            reg_file[22947] <= 8'h00;
            reg_file[22948] <= 8'h00;
            reg_file[22949] <= 8'h00;
            reg_file[22950] <= 8'h00;
            reg_file[22951] <= 8'h00;
            reg_file[22952] <= 8'h00;
            reg_file[22953] <= 8'h00;
            reg_file[22954] <= 8'h00;
            reg_file[22955] <= 8'h00;
            reg_file[22956] <= 8'h00;
            reg_file[22957] <= 8'h00;
            reg_file[22958] <= 8'h00;
            reg_file[22959] <= 8'h00;
            reg_file[22960] <= 8'h00;
            reg_file[22961] <= 8'h00;
            reg_file[22962] <= 8'h00;
            reg_file[22963] <= 8'h00;
            reg_file[22964] <= 8'h00;
            reg_file[22965] <= 8'h00;
            reg_file[22966] <= 8'h00;
            reg_file[22967] <= 8'h00;
            reg_file[22968] <= 8'h00;
            reg_file[22969] <= 8'h00;
            reg_file[22970] <= 8'h00;
            reg_file[22971] <= 8'h00;
            reg_file[22972] <= 8'h00;
            reg_file[22973] <= 8'h00;
            reg_file[22974] <= 8'h00;
            reg_file[22975] <= 8'h00;
            reg_file[22976] <= 8'h00;
            reg_file[22977] <= 8'h00;
            reg_file[22978] <= 8'h00;
            reg_file[22979] <= 8'h00;
            reg_file[22980] <= 8'h00;
            reg_file[22981] <= 8'h00;
            reg_file[22982] <= 8'h00;
            reg_file[22983] <= 8'h00;
            reg_file[22984] <= 8'h00;
            reg_file[22985] <= 8'h00;
            reg_file[22986] <= 8'h00;
            reg_file[22987] <= 8'h00;
            reg_file[22988] <= 8'h00;
            reg_file[22989] <= 8'h00;
            reg_file[22990] <= 8'h00;
            reg_file[22991] <= 8'h00;
            reg_file[22992] <= 8'h00;
            reg_file[22993] <= 8'h00;
            reg_file[22994] <= 8'h00;
            reg_file[22995] <= 8'h00;
            reg_file[22996] <= 8'h00;
            reg_file[22997] <= 8'h00;
            reg_file[22998] <= 8'h00;
            reg_file[22999] <= 8'h00;
            reg_file[23000] <= 8'h00;
            reg_file[23001] <= 8'h00;
            reg_file[23002] <= 8'h00;
            reg_file[23003] <= 8'h00;
            reg_file[23004] <= 8'h00;
            reg_file[23005] <= 8'h00;
            reg_file[23006] <= 8'h00;
            reg_file[23007] <= 8'h00;
            reg_file[23008] <= 8'h00;
            reg_file[23009] <= 8'h00;
            reg_file[23010] <= 8'h00;
            reg_file[23011] <= 8'h00;
            reg_file[23012] <= 8'h00;
            reg_file[23013] <= 8'h00;
            reg_file[23014] <= 8'h00;
            reg_file[23015] <= 8'h00;
            reg_file[23016] <= 8'h00;
            reg_file[23017] <= 8'h00;
            reg_file[23018] <= 8'h00;
            reg_file[23019] <= 8'h00;
            reg_file[23020] <= 8'h00;
            reg_file[23021] <= 8'h00;
            reg_file[23022] <= 8'h00;
            reg_file[23023] <= 8'h00;
            reg_file[23024] <= 8'h00;
            reg_file[23025] <= 8'h00;
            reg_file[23026] <= 8'h00;
            reg_file[23027] <= 8'h00;
            reg_file[23028] <= 8'h00;
            reg_file[23029] <= 8'h00;
            reg_file[23030] <= 8'h00;
            reg_file[23031] <= 8'h00;
            reg_file[23032] <= 8'h00;
            reg_file[23033] <= 8'h00;
            reg_file[23034] <= 8'h00;
            reg_file[23035] <= 8'h00;
            reg_file[23036] <= 8'h00;
            reg_file[23037] <= 8'h00;
            reg_file[23038] <= 8'h00;
            reg_file[23039] <= 8'h00;
            reg_file[23040] <= 8'h00;
            reg_file[23041] <= 8'h00;
            reg_file[23042] <= 8'h00;
            reg_file[23043] <= 8'h00;
            reg_file[23044] <= 8'h00;
            reg_file[23045] <= 8'h00;
            reg_file[23046] <= 8'h00;
            reg_file[23047] <= 8'h00;
            reg_file[23048] <= 8'h00;
            reg_file[23049] <= 8'h00;
            reg_file[23050] <= 8'h00;
            reg_file[23051] <= 8'h00;
            reg_file[23052] <= 8'h00;
            reg_file[23053] <= 8'h00;
            reg_file[23054] <= 8'h00;
            reg_file[23055] <= 8'h00;
            reg_file[23056] <= 8'h00;
            reg_file[23057] <= 8'h00;
            reg_file[23058] <= 8'h00;
            reg_file[23059] <= 8'h00;
            reg_file[23060] <= 8'h00;
            reg_file[23061] <= 8'h00;
            reg_file[23062] <= 8'h00;
            reg_file[23063] <= 8'h00;
            reg_file[23064] <= 8'h00;
            reg_file[23065] <= 8'h00;
            reg_file[23066] <= 8'h00;
            reg_file[23067] <= 8'h00;
            reg_file[23068] <= 8'h00;
            reg_file[23069] <= 8'h00;
            reg_file[23070] <= 8'h00;
            reg_file[23071] <= 8'h00;
            reg_file[23072] <= 8'h00;
            reg_file[23073] <= 8'h00;
            reg_file[23074] <= 8'h00;
            reg_file[23075] <= 8'h00;
            reg_file[23076] <= 8'h00;
            reg_file[23077] <= 8'h00;
            reg_file[23078] <= 8'h00;
            reg_file[23079] <= 8'h00;
            reg_file[23080] <= 8'h00;
            reg_file[23081] <= 8'h00;
            reg_file[23082] <= 8'h00;
            reg_file[23083] <= 8'h00;
            reg_file[23084] <= 8'h00;
            reg_file[23085] <= 8'h00;
            reg_file[23086] <= 8'h00;
            reg_file[23087] <= 8'h00;
            reg_file[23088] <= 8'h00;
            reg_file[23089] <= 8'h00;
            reg_file[23090] <= 8'h00;
            reg_file[23091] <= 8'h00;
            reg_file[23092] <= 8'h00;
            reg_file[23093] <= 8'h00;
            reg_file[23094] <= 8'h00;
            reg_file[23095] <= 8'h00;
            reg_file[23096] <= 8'h00;
            reg_file[23097] <= 8'h00;
            reg_file[23098] <= 8'h00;
            reg_file[23099] <= 8'h00;
            reg_file[23100] <= 8'h00;
            reg_file[23101] <= 8'h00;
            reg_file[23102] <= 8'h00;
            reg_file[23103] <= 8'h00;
            reg_file[23104] <= 8'h00;
            reg_file[23105] <= 8'h00;
            reg_file[23106] <= 8'h00;
            reg_file[23107] <= 8'h00;
            reg_file[23108] <= 8'h00;
            reg_file[23109] <= 8'h00;
            reg_file[23110] <= 8'h00;
            reg_file[23111] <= 8'h00;
            reg_file[23112] <= 8'h00;
            reg_file[23113] <= 8'h00;
            reg_file[23114] <= 8'h00;
            reg_file[23115] <= 8'h00;
            reg_file[23116] <= 8'h00;
            reg_file[23117] <= 8'h00;
            reg_file[23118] <= 8'h00;
            reg_file[23119] <= 8'h00;
            reg_file[23120] <= 8'h00;
            reg_file[23121] <= 8'h00;
            reg_file[23122] <= 8'h00;
            reg_file[23123] <= 8'h00;
            reg_file[23124] <= 8'h00;
            reg_file[23125] <= 8'h00;
            reg_file[23126] <= 8'h00;
            reg_file[23127] <= 8'h00;
            reg_file[23128] <= 8'h00;
            reg_file[23129] <= 8'h00;
            reg_file[23130] <= 8'h00;
            reg_file[23131] <= 8'h00;
            reg_file[23132] <= 8'h00;
            reg_file[23133] <= 8'h00;
            reg_file[23134] <= 8'h00;
            reg_file[23135] <= 8'h00;
            reg_file[23136] <= 8'h00;
            reg_file[23137] <= 8'h00;
            reg_file[23138] <= 8'h00;
            reg_file[23139] <= 8'h00;
            reg_file[23140] <= 8'h00;
            reg_file[23141] <= 8'h00;
            reg_file[23142] <= 8'h00;
            reg_file[23143] <= 8'h00;
            reg_file[23144] <= 8'h00;
            reg_file[23145] <= 8'h00;
            reg_file[23146] <= 8'h00;
            reg_file[23147] <= 8'h00;
            reg_file[23148] <= 8'h00;
            reg_file[23149] <= 8'h00;
            reg_file[23150] <= 8'h00;
            reg_file[23151] <= 8'h00;
            reg_file[23152] <= 8'h00;
            reg_file[23153] <= 8'h00;
            reg_file[23154] <= 8'h00;
            reg_file[23155] <= 8'h00;
            reg_file[23156] <= 8'h00;
            reg_file[23157] <= 8'h00;
            reg_file[23158] <= 8'h00;
            reg_file[23159] <= 8'h00;
            reg_file[23160] <= 8'h00;
            reg_file[23161] <= 8'h00;
            reg_file[23162] <= 8'h00;
            reg_file[23163] <= 8'h00;
            reg_file[23164] <= 8'h00;
            reg_file[23165] <= 8'h00;
            reg_file[23166] <= 8'h00;
            reg_file[23167] <= 8'h00;
            reg_file[23168] <= 8'h00;
            reg_file[23169] <= 8'h00;
            reg_file[23170] <= 8'h00;
            reg_file[23171] <= 8'h00;
            reg_file[23172] <= 8'h00;
            reg_file[23173] <= 8'h00;
            reg_file[23174] <= 8'h00;
            reg_file[23175] <= 8'h00;
            reg_file[23176] <= 8'h00;
            reg_file[23177] <= 8'h00;
            reg_file[23178] <= 8'h00;
            reg_file[23179] <= 8'h00;
            reg_file[23180] <= 8'h00;
            reg_file[23181] <= 8'h00;
            reg_file[23182] <= 8'h00;
            reg_file[23183] <= 8'h00;
            reg_file[23184] <= 8'h00;
            reg_file[23185] <= 8'h00;
            reg_file[23186] <= 8'h00;
            reg_file[23187] <= 8'h00;
            reg_file[23188] <= 8'h00;
            reg_file[23189] <= 8'h00;
            reg_file[23190] <= 8'h00;
            reg_file[23191] <= 8'h00;
            reg_file[23192] <= 8'h00;
            reg_file[23193] <= 8'h00;
            reg_file[23194] <= 8'h00;
            reg_file[23195] <= 8'h00;
            reg_file[23196] <= 8'h00;
            reg_file[23197] <= 8'h00;
            reg_file[23198] <= 8'h00;
            reg_file[23199] <= 8'h00;
            reg_file[23200] <= 8'h00;
            reg_file[23201] <= 8'h00;
            reg_file[23202] <= 8'h00;
            reg_file[23203] <= 8'h00;
            reg_file[23204] <= 8'h00;
            reg_file[23205] <= 8'h00;
            reg_file[23206] <= 8'h00;
            reg_file[23207] <= 8'h00;
            reg_file[23208] <= 8'h00;
            reg_file[23209] <= 8'h00;
            reg_file[23210] <= 8'h00;
            reg_file[23211] <= 8'h00;
            reg_file[23212] <= 8'h00;
            reg_file[23213] <= 8'h00;
            reg_file[23214] <= 8'h00;
            reg_file[23215] <= 8'h00;
            reg_file[23216] <= 8'h00;
            reg_file[23217] <= 8'h00;
            reg_file[23218] <= 8'h00;
            reg_file[23219] <= 8'h00;
            reg_file[23220] <= 8'h00;
            reg_file[23221] <= 8'h00;
            reg_file[23222] <= 8'h00;
            reg_file[23223] <= 8'h00;
            reg_file[23224] <= 8'h00;
            reg_file[23225] <= 8'h00;
            reg_file[23226] <= 8'h00;
            reg_file[23227] <= 8'h00;
            reg_file[23228] <= 8'h00;
            reg_file[23229] <= 8'h00;
            reg_file[23230] <= 8'h00;
            reg_file[23231] <= 8'h00;
            reg_file[23232] <= 8'h00;
            reg_file[23233] <= 8'h00;
            reg_file[23234] <= 8'h00;
            reg_file[23235] <= 8'h00;
            reg_file[23236] <= 8'h00;
            reg_file[23237] <= 8'h00;
            reg_file[23238] <= 8'h00;
            reg_file[23239] <= 8'h00;
            reg_file[23240] <= 8'h00;
            reg_file[23241] <= 8'h00;
            reg_file[23242] <= 8'h00;
            reg_file[23243] <= 8'h00;
            reg_file[23244] <= 8'h00;
            reg_file[23245] <= 8'h00;
            reg_file[23246] <= 8'h00;
            reg_file[23247] <= 8'h00;
            reg_file[23248] <= 8'h00;
            reg_file[23249] <= 8'h00;
            reg_file[23250] <= 8'h00;
            reg_file[23251] <= 8'h00;
            reg_file[23252] <= 8'h00;
            reg_file[23253] <= 8'h00;
            reg_file[23254] <= 8'h00;
            reg_file[23255] <= 8'h00;
            reg_file[23256] <= 8'h00;
            reg_file[23257] <= 8'h00;
            reg_file[23258] <= 8'h00;
            reg_file[23259] <= 8'h00;
            reg_file[23260] <= 8'h00;
            reg_file[23261] <= 8'h00;
            reg_file[23262] <= 8'h00;
            reg_file[23263] <= 8'h00;
            reg_file[23264] <= 8'h00;
            reg_file[23265] <= 8'h00;
            reg_file[23266] <= 8'h00;
            reg_file[23267] <= 8'h00;
            reg_file[23268] <= 8'h00;
            reg_file[23269] <= 8'h00;
            reg_file[23270] <= 8'h00;
            reg_file[23271] <= 8'h00;
            reg_file[23272] <= 8'h00;
            reg_file[23273] <= 8'h00;
            reg_file[23274] <= 8'h00;
            reg_file[23275] <= 8'h00;
            reg_file[23276] <= 8'h00;
            reg_file[23277] <= 8'h00;
            reg_file[23278] <= 8'h00;
            reg_file[23279] <= 8'h00;
            reg_file[23280] <= 8'h00;
            reg_file[23281] <= 8'h00;
            reg_file[23282] <= 8'h00;
            reg_file[23283] <= 8'h00;
            reg_file[23284] <= 8'h00;
            reg_file[23285] <= 8'h00;
            reg_file[23286] <= 8'h00;
            reg_file[23287] <= 8'h00;
            reg_file[23288] <= 8'h00;
            reg_file[23289] <= 8'h00;
            reg_file[23290] <= 8'h00;
            reg_file[23291] <= 8'h00;
            reg_file[23292] <= 8'h00;
            reg_file[23293] <= 8'h00;
            reg_file[23294] <= 8'h00;
            reg_file[23295] <= 8'h00;
            reg_file[23296] <= 8'h00;
            reg_file[23297] <= 8'h00;
            reg_file[23298] <= 8'h00;
            reg_file[23299] <= 8'h00;
            reg_file[23300] <= 8'h00;
            reg_file[23301] <= 8'h00;
            reg_file[23302] <= 8'h00;
            reg_file[23303] <= 8'h00;
            reg_file[23304] <= 8'h00;
            reg_file[23305] <= 8'h00;
            reg_file[23306] <= 8'h00;
            reg_file[23307] <= 8'h00;
            reg_file[23308] <= 8'h00;
            reg_file[23309] <= 8'h00;
            reg_file[23310] <= 8'h00;
            reg_file[23311] <= 8'h00;
            reg_file[23312] <= 8'h00;
            reg_file[23313] <= 8'h00;
            reg_file[23314] <= 8'h00;
            reg_file[23315] <= 8'h00;
            reg_file[23316] <= 8'h00;
            reg_file[23317] <= 8'h00;
            reg_file[23318] <= 8'h00;
            reg_file[23319] <= 8'h00;
            reg_file[23320] <= 8'h00;
            reg_file[23321] <= 8'h00;
            reg_file[23322] <= 8'h00;
            reg_file[23323] <= 8'h00;
            reg_file[23324] <= 8'h00;
            reg_file[23325] <= 8'h00;
            reg_file[23326] <= 8'h00;
            reg_file[23327] <= 8'h00;
            reg_file[23328] <= 8'h00;
            reg_file[23329] <= 8'h00;
            reg_file[23330] <= 8'h00;
            reg_file[23331] <= 8'h00;
            reg_file[23332] <= 8'h00;
            reg_file[23333] <= 8'h00;
            reg_file[23334] <= 8'h00;
            reg_file[23335] <= 8'h00;
            reg_file[23336] <= 8'h00;
            reg_file[23337] <= 8'h00;
            reg_file[23338] <= 8'h00;
            reg_file[23339] <= 8'h00;
            reg_file[23340] <= 8'h00;
            reg_file[23341] <= 8'h00;
            reg_file[23342] <= 8'h00;
            reg_file[23343] <= 8'h00;
            reg_file[23344] <= 8'h00;
            reg_file[23345] <= 8'h00;
            reg_file[23346] <= 8'h00;
            reg_file[23347] <= 8'h00;
            reg_file[23348] <= 8'h00;
            reg_file[23349] <= 8'h00;
            reg_file[23350] <= 8'h00;
            reg_file[23351] <= 8'h00;
            reg_file[23352] <= 8'h00;
            reg_file[23353] <= 8'h00;
            reg_file[23354] <= 8'h00;
            reg_file[23355] <= 8'h00;
            reg_file[23356] <= 8'h00;
            reg_file[23357] <= 8'h00;
            reg_file[23358] <= 8'h00;
            reg_file[23359] <= 8'h00;
            reg_file[23360] <= 8'h00;
            reg_file[23361] <= 8'h00;
            reg_file[23362] <= 8'h00;
            reg_file[23363] <= 8'h00;
            reg_file[23364] <= 8'h00;
            reg_file[23365] <= 8'h00;
            reg_file[23366] <= 8'h00;
            reg_file[23367] <= 8'h00;
            reg_file[23368] <= 8'h00;
            reg_file[23369] <= 8'h00;
            reg_file[23370] <= 8'h00;
            reg_file[23371] <= 8'h00;
            reg_file[23372] <= 8'h00;
            reg_file[23373] <= 8'h00;
            reg_file[23374] <= 8'h00;
            reg_file[23375] <= 8'h00;
            reg_file[23376] <= 8'h00;
            reg_file[23377] <= 8'h00;
            reg_file[23378] <= 8'h00;
            reg_file[23379] <= 8'h00;
            reg_file[23380] <= 8'h00;
            reg_file[23381] <= 8'h00;
            reg_file[23382] <= 8'h00;
            reg_file[23383] <= 8'h00;
            reg_file[23384] <= 8'h00;
            reg_file[23385] <= 8'h00;
            reg_file[23386] <= 8'h00;
            reg_file[23387] <= 8'h00;
            reg_file[23388] <= 8'h00;
            reg_file[23389] <= 8'h00;
            reg_file[23390] <= 8'h00;
            reg_file[23391] <= 8'h00;
            reg_file[23392] <= 8'h00;
            reg_file[23393] <= 8'h00;
            reg_file[23394] <= 8'h00;
            reg_file[23395] <= 8'h00;
            reg_file[23396] <= 8'h00;
            reg_file[23397] <= 8'h00;
            reg_file[23398] <= 8'h00;
            reg_file[23399] <= 8'h00;
            reg_file[23400] <= 8'h00;
            reg_file[23401] <= 8'h00;
            reg_file[23402] <= 8'h00;
            reg_file[23403] <= 8'h00;
            reg_file[23404] <= 8'h00;
            reg_file[23405] <= 8'h00;
            reg_file[23406] <= 8'h00;
            reg_file[23407] <= 8'h00;
            reg_file[23408] <= 8'h00;
            reg_file[23409] <= 8'h00;
            reg_file[23410] <= 8'h00;
            reg_file[23411] <= 8'h00;
            reg_file[23412] <= 8'h00;
            reg_file[23413] <= 8'h00;
            reg_file[23414] <= 8'h00;
            reg_file[23415] <= 8'h00;
            reg_file[23416] <= 8'h00;
            reg_file[23417] <= 8'h00;
            reg_file[23418] <= 8'h00;
            reg_file[23419] <= 8'h00;
            reg_file[23420] <= 8'h00;
            reg_file[23421] <= 8'h00;
            reg_file[23422] <= 8'h00;
            reg_file[23423] <= 8'h00;
            reg_file[23424] <= 8'h00;
            reg_file[23425] <= 8'h00;
            reg_file[23426] <= 8'h00;
            reg_file[23427] <= 8'h00;
            reg_file[23428] <= 8'h00;
            reg_file[23429] <= 8'h00;
            reg_file[23430] <= 8'h00;
            reg_file[23431] <= 8'h00;
            reg_file[23432] <= 8'h00;
            reg_file[23433] <= 8'h00;
            reg_file[23434] <= 8'h00;
            reg_file[23435] <= 8'h00;
            reg_file[23436] <= 8'h00;
            reg_file[23437] <= 8'h00;
            reg_file[23438] <= 8'h00;
            reg_file[23439] <= 8'h00;
            reg_file[23440] <= 8'h00;
            reg_file[23441] <= 8'h00;
            reg_file[23442] <= 8'h00;
            reg_file[23443] <= 8'h00;
            reg_file[23444] <= 8'h00;
            reg_file[23445] <= 8'h00;
            reg_file[23446] <= 8'h00;
            reg_file[23447] <= 8'h00;
            reg_file[23448] <= 8'h00;
            reg_file[23449] <= 8'h00;
            reg_file[23450] <= 8'h00;
            reg_file[23451] <= 8'h00;
            reg_file[23452] <= 8'h00;
            reg_file[23453] <= 8'h00;
            reg_file[23454] <= 8'h00;
            reg_file[23455] <= 8'h00;
            reg_file[23456] <= 8'h00;
            reg_file[23457] <= 8'h00;
            reg_file[23458] <= 8'h00;
            reg_file[23459] <= 8'h00;
            reg_file[23460] <= 8'h00;
            reg_file[23461] <= 8'h00;
            reg_file[23462] <= 8'h00;
            reg_file[23463] <= 8'h00;
            reg_file[23464] <= 8'h00;
            reg_file[23465] <= 8'h00;
            reg_file[23466] <= 8'h00;
            reg_file[23467] <= 8'h00;
            reg_file[23468] <= 8'h00;
            reg_file[23469] <= 8'h00;
            reg_file[23470] <= 8'h00;
            reg_file[23471] <= 8'h00;
            reg_file[23472] <= 8'h00;
            reg_file[23473] <= 8'h00;
            reg_file[23474] <= 8'h00;
            reg_file[23475] <= 8'h00;
            reg_file[23476] <= 8'h00;
            reg_file[23477] <= 8'h00;
            reg_file[23478] <= 8'h00;
            reg_file[23479] <= 8'h00;
            reg_file[23480] <= 8'h00;
            reg_file[23481] <= 8'h00;
            reg_file[23482] <= 8'h00;
            reg_file[23483] <= 8'h00;
            reg_file[23484] <= 8'h00;
            reg_file[23485] <= 8'h00;
            reg_file[23486] <= 8'h00;
            reg_file[23487] <= 8'h00;
            reg_file[23488] <= 8'h00;
            reg_file[23489] <= 8'h00;
            reg_file[23490] <= 8'h00;
            reg_file[23491] <= 8'h00;
            reg_file[23492] <= 8'h00;
            reg_file[23493] <= 8'h00;
            reg_file[23494] <= 8'h00;
            reg_file[23495] <= 8'h00;
            reg_file[23496] <= 8'h00;
            reg_file[23497] <= 8'h00;
            reg_file[23498] <= 8'h00;
            reg_file[23499] <= 8'h00;
            reg_file[23500] <= 8'h00;
            reg_file[23501] <= 8'h00;
            reg_file[23502] <= 8'h00;
            reg_file[23503] <= 8'h00;
            reg_file[23504] <= 8'h00;
            reg_file[23505] <= 8'h00;
            reg_file[23506] <= 8'h00;
            reg_file[23507] <= 8'h00;
            reg_file[23508] <= 8'h00;
            reg_file[23509] <= 8'h00;
            reg_file[23510] <= 8'h00;
            reg_file[23511] <= 8'h00;
            reg_file[23512] <= 8'h00;
            reg_file[23513] <= 8'h00;
            reg_file[23514] <= 8'h00;
            reg_file[23515] <= 8'h00;
            reg_file[23516] <= 8'h00;
            reg_file[23517] <= 8'h00;
            reg_file[23518] <= 8'h00;
            reg_file[23519] <= 8'h00;
            reg_file[23520] <= 8'h00;
            reg_file[23521] <= 8'h00;
            reg_file[23522] <= 8'h00;
            reg_file[23523] <= 8'h00;
            reg_file[23524] <= 8'h00;
            reg_file[23525] <= 8'h00;
            reg_file[23526] <= 8'h00;
            reg_file[23527] <= 8'h00;
            reg_file[23528] <= 8'h00;
            reg_file[23529] <= 8'h00;
            reg_file[23530] <= 8'h00;
            reg_file[23531] <= 8'h00;
            reg_file[23532] <= 8'h00;
            reg_file[23533] <= 8'h00;
            reg_file[23534] <= 8'h00;
            reg_file[23535] <= 8'h00;
            reg_file[23536] <= 8'h00;
            reg_file[23537] <= 8'h00;
            reg_file[23538] <= 8'h00;
            reg_file[23539] <= 8'h00;
            reg_file[23540] <= 8'h00;
            reg_file[23541] <= 8'h00;
            reg_file[23542] <= 8'h00;
            reg_file[23543] <= 8'h00;
            reg_file[23544] <= 8'h00;
            reg_file[23545] <= 8'h00;
            reg_file[23546] <= 8'h00;
            reg_file[23547] <= 8'h00;
            reg_file[23548] <= 8'h00;
            reg_file[23549] <= 8'h00;
            reg_file[23550] <= 8'h00;
            reg_file[23551] <= 8'h00;
            reg_file[23552] <= 8'h00;
            reg_file[23553] <= 8'h00;
            reg_file[23554] <= 8'h00;
            reg_file[23555] <= 8'h00;
            reg_file[23556] <= 8'h00;
            reg_file[23557] <= 8'h00;
            reg_file[23558] <= 8'h00;
            reg_file[23559] <= 8'h00;
            reg_file[23560] <= 8'h00;
            reg_file[23561] <= 8'h00;
            reg_file[23562] <= 8'h00;
            reg_file[23563] <= 8'h00;
            reg_file[23564] <= 8'h00;
            reg_file[23565] <= 8'h00;
            reg_file[23566] <= 8'h00;
            reg_file[23567] <= 8'h00;
            reg_file[23568] <= 8'h00;
            reg_file[23569] <= 8'h00;
            reg_file[23570] <= 8'h00;
            reg_file[23571] <= 8'h00;
            reg_file[23572] <= 8'h00;
            reg_file[23573] <= 8'h00;
            reg_file[23574] <= 8'h00;
            reg_file[23575] <= 8'h00;
            reg_file[23576] <= 8'h00;
            reg_file[23577] <= 8'h00;
            reg_file[23578] <= 8'h00;
            reg_file[23579] <= 8'h00;
            reg_file[23580] <= 8'h00;
            reg_file[23581] <= 8'h00;
            reg_file[23582] <= 8'h00;
            reg_file[23583] <= 8'h00;
            reg_file[23584] <= 8'h00;
            reg_file[23585] <= 8'h00;
            reg_file[23586] <= 8'h00;
            reg_file[23587] <= 8'h00;
            reg_file[23588] <= 8'h00;
            reg_file[23589] <= 8'h00;
            reg_file[23590] <= 8'h00;
            reg_file[23591] <= 8'h00;
            reg_file[23592] <= 8'h00;
            reg_file[23593] <= 8'h00;
            reg_file[23594] <= 8'h00;
            reg_file[23595] <= 8'h00;
            reg_file[23596] <= 8'h00;
            reg_file[23597] <= 8'h00;
            reg_file[23598] <= 8'h00;
            reg_file[23599] <= 8'h00;
            reg_file[23600] <= 8'h00;
            reg_file[23601] <= 8'h00;
            reg_file[23602] <= 8'h00;
            reg_file[23603] <= 8'h00;
            reg_file[23604] <= 8'h00;
            reg_file[23605] <= 8'h00;
            reg_file[23606] <= 8'h00;
            reg_file[23607] <= 8'h00;
            reg_file[23608] <= 8'h00;
            reg_file[23609] <= 8'h00;
            reg_file[23610] <= 8'h00;
            reg_file[23611] <= 8'h00;
            reg_file[23612] <= 8'h00;
            reg_file[23613] <= 8'h00;
            reg_file[23614] <= 8'h00;
            reg_file[23615] <= 8'h00;
            reg_file[23616] <= 8'h00;
            reg_file[23617] <= 8'h00;
            reg_file[23618] <= 8'h00;
            reg_file[23619] <= 8'h00;
            reg_file[23620] <= 8'h00;
            reg_file[23621] <= 8'h00;
            reg_file[23622] <= 8'h00;
            reg_file[23623] <= 8'h00;
            reg_file[23624] <= 8'h00;
            reg_file[23625] <= 8'h00;
            reg_file[23626] <= 8'h00;
            reg_file[23627] <= 8'h00;
            reg_file[23628] <= 8'h00;
            reg_file[23629] <= 8'h00;
            reg_file[23630] <= 8'h00;
            reg_file[23631] <= 8'h00;
            reg_file[23632] <= 8'h00;
            reg_file[23633] <= 8'h00;
            reg_file[23634] <= 8'h00;
            reg_file[23635] <= 8'h00;
            reg_file[23636] <= 8'h00;
            reg_file[23637] <= 8'h00;
            reg_file[23638] <= 8'h00;
            reg_file[23639] <= 8'h00;
            reg_file[23640] <= 8'h00;
            reg_file[23641] <= 8'h00;
            reg_file[23642] <= 8'h00;
            reg_file[23643] <= 8'h00;
            reg_file[23644] <= 8'h00;
            reg_file[23645] <= 8'h00;
            reg_file[23646] <= 8'h00;
            reg_file[23647] <= 8'h00;
            reg_file[23648] <= 8'h00;
            reg_file[23649] <= 8'h00;
            reg_file[23650] <= 8'h00;
            reg_file[23651] <= 8'h00;
            reg_file[23652] <= 8'h00;
            reg_file[23653] <= 8'h00;
            reg_file[23654] <= 8'h00;
            reg_file[23655] <= 8'h00;
            reg_file[23656] <= 8'h00;
            reg_file[23657] <= 8'h00;
            reg_file[23658] <= 8'h00;
            reg_file[23659] <= 8'h00;
            reg_file[23660] <= 8'h00;
            reg_file[23661] <= 8'h00;
            reg_file[23662] <= 8'h00;
            reg_file[23663] <= 8'h00;
            reg_file[23664] <= 8'h00;
            reg_file[23665] <= 8'h00;
            reg_file[23666] <= 8'h00;
            reg_file[23667] <= 8'h00;
            reg_file[23668] <= 8'h00;
            reg_file[23669] <= 8'h00;
            reg_file[23670] <= 8'h00;
            reg_file[23671] <= 8'h00;
            reg_file[23672] <= 8'h00;
            reg_file[23673] <= 8'h00;
            reg_file[23674] <= 8'h00;
            reg_file[23675] <= 8'h00;
            reg_file[23676] <= 8'h00;
            reg_file[23677] <= 8'h00;
            reg_file[23678] <= 8'h00;
            reg_file[23679] <= 8'h00;
            reg_file[23680] <= 8'h00;
            reg_file[23681] <= 8'h00;
            reg_file[23682] <= 8'h00;
            reg_file[23683] <= 8'h00;
            reg_file[23684] <= 8'h00;
            reg_file[23685] <= 8'h00;
            reg_file[23686] <= 8'h00;
            reg_file[23687] <= 8'h00;
            reg_file[23688] <= 8'h00;
            reg_file[23689] <= 8'h00;
            reg_file[23690] <= 8'h00;
            reg_file[23691] <= 8'h00;
            reg_file[23692] <= 8'h00;
            reg_file[23693] <= 8'h00;
            reg_file[23694] <= 8'h00;
            reg_file[23695] <= 8'h00;
            reg_file[23696] <= 8'h00;
            reg_file[23697] <= 8'h00;
            reg_file[23698] <= 8'h00;
            reg_file[23699] <= 8'h00;
            reg_file[23700] <= 8'h00;
            reg_file[23701] <= 8'h00;
            reg_file[23702] <= 8'h00;
            reg_file[23703] <= 8'h00;
            reg_file[23704] <= 8'h00;
            reg_file[23705] <= 8'h00;
            reg_file[23706] <= 8'h00;
            reg_file[23707] <= 8'h00;
            reg_file[23708] <= 8'h00;
            reg_file[23709] <= 8'h00;
            reg_file[23710] <= 8'h00;
            reg_file[23711] <= 8'h00;
            reg_file[23712] <= 8'h00;
            reg_file[23713] <= 8'h00;
            reg_file[23714] <= 8'h00;
            reg_file[23715] <= 8'h00;
            reg_file[23716] <= 8'h00;
            reg_file[23717] <= 8'h00;
            reg_file[23718] <= 8'h00;
            reg_file[23719] <= 8'h00;
            reg_file[23720] <= 8'h00;
            reg_file[23721] <= 8'h00;
            reg_file[23722] <= 8'h00;
            reg_file[23723] <= 8'h00;
            reg_file[23724] <= 8'h00;
            reg_file[23725] <= 8'h00;
            reg_file[23726] <= 8'h00;
            reg_file[23727] <= 8'h00;
            reg_file[23728] <= 8'h00;
            reg_file[23729] <= 8'h00;
            reg_file[23730] <= 8'h00;
            reg_file[23731] <= 8'h00;
            reg_file[23732] <= 8'h00;
            reg_file[23733] <= 8'h00;
            reg_file[23734] <= 8'h00;
            reg_file[23735] <= 8'h00;
            reg_file[23736] <= 8'h00;
            reg_file[23737] <= 8'h00;
            reg_file[23738] <= 8'h00;
            reg_file[23739] <= 8'h00;
            reg_file[23740] <= 8'h00;
            reg_file[23741] <= 8'h00;
            reg_file[23742] <= 8'h00;
            reg_file[23743] <= 8'h00;
            reg_file[23744] <= 8'h00;
            reg_file[23745] <= 8'h00;
            reg_file[23746] <= 8'h00;
            reg_file[23747] <= 8'h00;
            reg_file[23748] <= 8'h00;
            reg_file[23749] <= 8'h00;
            reg_file[23750] <= 8'h00;
            reg_file[23751] <= 8'h00;
            reg_file[23752] <= 8'h00;
            reg_file[23753] <= 8'h00;
            reg_file[23754] <= 8'h00;
            reg_file[23755] <= 8'h00;
            reg_file[23756] <= 8'h00;
            reg_file[23757] <= 8'h00;
            reg_file[23758] <= 8'h00;
            reg_file[23759] <= 8'h00;
            reg_file[23760] <= 8'h00;
            reg_file[23761] <= 8'h00;
            reg_file[23762] <= 8'h00;
            reg_file[23763] <= 8'h00;
            reg_file[23764] <= 8'h00;
            reg_file[23765] <= 8'h00;
            reg_file[23766] <= 8'h00;
            reg_file[23767] <= 8'h00;
            reg_file[23768] <= 8'h00;
            reg_file[23769] <= 8'h00;
            reg_file[23770] <= 8'h00;
            reg_file[23771] <= 8'h00;
            reg_file[23772] <= 8'h00;
            reg_file[23773] <= 8'h00;
            reg_file[23774] <= 8'h00;
            reg_file[23775] <= 8'h00;
            reg_file[23776] <= 8'h00;
            reg_file[23777] <= 8'h00;
            reg_file[23778] <= 8'h00;
            reg_file[23779] <= 8'h00;
            reg_file[23780] <= 8'h00;
            reg_file[23781] <= 8'h00;
            reg_file[23782] <= 8'h00;
            reg_file[23783] <= 8'h00;
            reg_file[23784] <= 8'h00;
            reg_file[23785] <= 8'h00;
            reg_file[23786] <= 8'h00;
            reg_file[23787] <= 8'h00;
            reg_file[23788] <= 8'h00;
            reg_file[23789] <= 8'h00;
            reg_file[23790] <= 8'h00;
            reg_file[23791] <= 8'h00;
            reg_file[23792] <= 8'h00;
            reg_file[23793] <= 8'h00;
            reg_file[23794] <= 8'h00;
            reg_file[23795] <= 8'h00;
            reg_file[23796] <= 8'h00;
            reg_file[23797] <= 8'h00;
            reg_file[23798] <= 8'h00;
            reg_file[23799] <= 8'h00;
            reg_file[23800] <= 8'h00;
            reg_file[23801] <= 8'h00;
            reg_file[23802] <= 8'h00;
            reg_file[23803] <= 8'h00;
            reg_file[23804] <= 8'h00;
            reg_file[23805] <= 8'h00;
            reg_file[23806] <= 8'h00;
            reg_file[23807] <= 8'h00;
            reg_file[23808] <= 8'h00;
            reg_file[23809] <= 8'h00;
            reg_file[23810] <= 8'h00;
            reg_file[23811] <= 8'h00;
            reg_file[23812] <= 8'h00;
            reg_file[23813] <= 8'h00;
            reg_file[23814] <= 8'h00;
            reg_file[23815] <= 8'h00;
            reg_file[23816] <= 8'h00;
            reg_file[23817] <= 8'h00;
            reg_file[23818] <= 8'h00;
            reg_file[23819] <= 8'h00;
            reg_file[23820] <= 8'h00;
            reg_file[23821] <= 8'h00;
            reg_file[23822] <= 8'h00;
            reg_file[23823] <= 8'h00;
            reg_file[23824] <= 8'h00;
            reg_file[23825] <= 8'h00;
            reg_file[23826] <= 8'h00;
            reg_file[23827] <= 8'h00;
            reg_file[23828] <= 8'h00;
            reg_file[23829] <= 8'h00;
            reg_file[23830] <= 8'h00;
            reg_file[23831] <= 8'h00;
            reg_file[23832] <= 8'h00;
            reg_file[23833] <= 8'h00;
            reg_file[23834] <= 8'h00;
            reg_file[23835] <= 8'h00;
            reg_file[23836] <= 8'h00;
            reg_file[23837] <= 8'h00;
            reg_file[23838] <= 8'h00;
            reg_file[23839] <= 8'h00;
            reg_file[23840] <= 8'h00;
            reg_file[23841] <= 8'h00;
            reg_file[23842] <= 8'h00;
            reg_file[23843] <= 8'h00;
            reg_file[23844] <= 8'h00;
            reg_file[23845] <= 8'h00;
            reg_file[23846] <= 8'h00;
            reg_file[23847] <= 8'h00;
            reg_file[23848] <= 8'h00;
            reg_file[23849] <= 8'h00;
            reg_file[23850] <= 8'h00;
            reg_file[23851] <= 8'h00;
            reg_file[23852] <= 8'h00;
            reg_file[23853] <= 8'h00;
            reg_file[23854] <= 8'h00;
            reg_file[23855] <= 8'h00;
            reg_file[23856] <= 8'h00;
            reg_file[23857] <= 8'h00;
            reg_file[23858] <= 8'h00;
            reg_file[23859] <= 8'h00;
            reg_file[23860] <= 8'h00;
            reg_file[23861] <= 8'h00;
            reg_file[23862] <= 8'h00;
            reg_file[23863] <= 8'h00;
            reg_file[23864] <= 8'h00;
            reg_file[23865] <= 8'h00;
            reg_file[23866] <= 8'h00;
            reg_file[23867] <= 8'h00;
            reg_file[23868] <= 8'h00;
            reg_file[23869] <= 8'h00;
            reg_file[23870] <= 8'h00;
            reg_file[23871] <= 8'h00;
            reg_file[23872] <= 8'h00;
            reg_file[23873] <= 8'h00;
            reg_file[23874] <= 8'h00;
            reg_file[23875] <= 8'h00;
            reg_file[23876] <= 8'h00;
            reg_file[23877] <= 8'h00;
            reg_file[23878] <= 8'h00;
            reg_file[23879] <= 8'h00;
            reg_file[23880] <= 8'h00;
            reg_file[23881] <= 8'h00;
            reg_file[23882] <= 8'h00;
            reg_file[23883] <= 8'h00;
            reg_file[23884] <= 8'h00;
            reg_file[23885] <= 8'h00;
            reg_file[23886] <= 8'h00;
            reg_file[23887] <= 8'h00;
            reg_file[23888] <= 8'h00;
            reg_file[23889] <= 8'h00;
            reg_file[23890] <= 8'h00;
            reg_file[23891] <= 8'h00;
            reg_file[23892] <= 8'h00;
            reg_file[23893] <= 8'h00;
            reg_file[23894] <= 8'h00;
            reg_file[23895] <= 8'h00;
            reg_file[23896] <= 8'h00;
            reg_file[23897] <= 8'h00;
            reg_file[23898] <= 8'h00;
            reg_file[23899] <= 8'h00;
            reg_file[23900] <= 8'h00;
            reg_file[23901] <= 8'h00;
            reg_file[23902] <= 8'h00;
            reg_file[23903] <= 8'h00;
            reg_file[23904] <= 8'h00;
            reg_file[23905] <= 8'h00;
            reg_file[23906] <= 8'h00;
            reg_file[23907] <= 8'h00;
            reg_file[23908] <= 8'h00;
            reg_file[23909] <= 8'h00;
            reg_file[23910] <= 8'h00;
            reg_file[23911] <= 8'h00;
            reg_file[23912] <= 8'h00;
            reg_file[23913] <= 8'h00;
            reg_file[23914] <= 8'h00;
            reg_file[23915] <= 8'h00;
            reg_file[23916] <= 8'h00;
            reg_file[23917] <= 8'h00;
            reg_file[23918] <= 8'h00;
            reg_file[23919] <= 8'h00;
            reg_file[23920] <= 8'h00;
            reg_file[23921] <= 8'h00;
            reg_file[23922] <= 8'h00;
            reg_file[23923] <= 8'h00;
            reg_file[23924] <= 8'h00;
            reg_file[23925] <= 8'h00;
            reg_file[23926] <= 8'h00;
            reg_file[23927] <= 8'h00;
            reg_file[23928] <= 8'h00;
            reg_file[23929] <= 8'h00;
            reg_file[23930] <= 8'h00;
            reg_file[23931] <= 8'h00;
            reg_file[23932] <= 8'h00;
            reg_file[23933] <= 8'h00;
            reg_file[23934] <= 8'h00;
            reg_file[23935] <= 8'h00;
            reg_file[23936] <= 8'h00;
            reg_file[23937] <= 8'h00;
            reg_file[23938] <= 8'h00;
            reg_file[23939] <= 8'h00;
            reg_file[23940] <= 8'h00;
            reg_file[23941] <= 8'h00;
            reg_file[23942] <= 8'h00;
            reg_file[23943] <= 8'h00;
            reg_file[23944] <= 8'h00;
            reg_file[23945] <= 8'h00;
            reg_file[23946] <= 8'h00;
            reg_file[23947] <= 8'h00;
            reg_file[23948] <= 8'h00;
            reg_file[23949] <= 8'h00;
            reg_file[23950] <= 8'h00;
            reg_file[23951] <= 8'h00;
            reg_file[23952] <= 8'h00;
            reg_file[23953] <= 8'h00;
            reg_file[23954] <= 8'h00;
            reg_file[23955] <= 8'h00;
            reg_file[23956] <= 8'h00;
            reg_file[23957] <= 8'h00;
            reg_file[23958] <= 8'h00;
            reg_file[23959] <= 8'h00;
            reg_file[23960] <= 8'h00;
            reg_file[23961] <= 8'h00;
            reg_file[23962] <= 8'h00;
            reg_file[23963] <= 8'h00;
            reg_file[23964] <= 8'h00;
            reg_file[23965] <= 8'h00;
            reg_file[23966] <= 8'h00;
            reg_file[23967] <= 8'h00;
            reg_file[23968] <= 8'h00;
            reg_file[23969] <= 8'h00;
            reg_file[23970] <= 8'h00;
            reg_file[23971] <= 8'h00;
            reg_file[23972] <= 8'h00;
            reg_file[23973] <= 8'h00;
            reg_file[23974] <= 8'h00;
            reg_file[23975] <= 8'h00;
            reg_file[23976] <= 8'h00;
            reg_file[23977] <= 8'h00;
            reg_file[23978] <= 8'h00;
            reg_file[23979] <= 8'h00;
            reg_file[23980] <= 8'h00;
            reg_file[23981] <= 8'h00;
            reg_file[23982] <= 8'h00;
            reg_file[23983] <= 8'h00;
            reg_file[23984] <= 8'h00;
            reg_file[23985] <= 8'h00;
            reg_file[23986] <= 8'h00;
            reg_file[23987] <= 8'h00;
            reg_file[23988] <= 8'h00;
            reg_file[23989] <= 8'h00;
            reg_file[23990] <= 8'h00;
            reg_file[23991] <= 8'h00;
            reg_file[23992] <= 8'h00;
            reg_file[23993] <= 8'h00;
            reg_file[23994] <= 8'h00;
            reg_file[23995] <= 8'h00;
            reg_file[23996] <= 8'h00;
            reg_file[23997] <= 8'h00;
            reg_file[23998] <= 8'h00;
            reg_file[23999] <= 8'h00;
            reg_file[24000] <= 8'h00;
            reg_file[24001] <= 8'h00;
            reg_file[24002] <= 8'h00;
            reg_file[24003] <= 8'h00;
            reg_file[24004] <= 8'h00;
            reg_file[24005] <= 8'h00;
            reg_file[24006] <= 8'h00;
            reg_file[24007] <= 8'h00;
            reg_file[24008] <= 8'h00;
            reg_file[24009] <= 8'h00;
            reg_file[24010] <= 8'h00;
            reg_file[24011] <= 8'h00;
            reg_file[24012] <= 8'h00;
            reg_file[24013] <= 8'h00;
            reg_file[24014] <= 8'h00;
            reg_file[24015] <= 8'h00;
            reg_file[24016] <= 8'h00;
            reg_file[24017] <= 8'h00;
            reg_file[24018] <= 8'h00;
            reg_file[24019] <= 8'h00;
            reg_file[24020] <= 8'h00;
            reg_file[24021] <= 8'h00;
            reg_file[24022] <= 8'h00;
            reg_file[24023] <= 8'h00;
            reg_file[24024] <= 8'h00;
            reg_file[24025] <= 8'h00;
            reg_file[24026] <= 8'h00;
            reg_file[24027] <= 8'h00;
            reg_file[24028] <= 8'h00;
            reg_file[24029] <= 8'h00;
            reg_file[24030] <= 8'h00;
            reg_file[24031] <= 8'h00;
            reg_file[24032] <= 8'h00;
            reg_file[24033] <= 8'h00;
            reg_file[24034] <= 8'h00;
            reg_file[24035] <= 8'h00;
            reg_file[24036] <= 8'h00;
            reg_file[24037] <= 8'h00;
            reg_file[24038] <= 8'h00;
            reg_file[24039] <= 8'h00;
            reg_file[24040] <= 8'h00;
            reg_file[24041] <= 8'h00;
            reg_file[24042] <= 8'h00;
            reg_file[24043] <= 8'h00;
            reg_file[24044] <= 8'h00;
            reg_file[24045] <= 8'h00;
            reg_file[24046] <= 8'h00;
            reg_file[24047] <= 8'h00;
            reg_file[24048] <= 8'h00;
            reg_file[24049] <= 8'h00;
            reg_file[24050] <= 8'h00;
            reg_file[24051] <= 8'h00;
            reg_file[24052] <= 8'h00;
            reg_file[24053] <= 8'h00;
            reg_file[24054] <= 8'h00;
            reg_file[24055] <= 8'h00;
            reg_file[24056] <= 8'h00;
            reg_file[24057] <= 8'h00;
            reg_file[24058] <= 8'h00;
            reg_file[24059] <= 8'h00;
            reg_file[24060] <= 8'h00;
            reg_file[24061] <= 8'h00;
            reg_file[24062] <= 8'h00;
            reg_file[24063] <= 8'h00;
            reg_file[24064] <= 8'h00;
            reg_file[24065] <= 8'h00;
            reg_file[24066] <= 8'h00;
            reg_file[24067] <= 8'h00;
            reg_file[24068] <= 8'h00;
            reg_file[24069] <= 8'h00;
            reg_file[24070] <= 8'h00;
            reg_file[24071] <= 8'h00;
            reg_file[24072] <= 8'h00;
            reg_file[24073] <= 8'h00;
            reg_file[24074] <= 8'h00;
            reg_file[24075] <= 8'h00;
            reg_file[24076] <= 8'h00;
            reg_file[24077] <= 8'h00;
            reg_file[24078] <= 8'h00;
            reg_file[24079] <= 8'h00;
            reg_file[24080] <= 8'h00;
            reg_file[24081] <= 8'h00;
            reg_file[24082] <= 8'h00;
            reg_file[24083] <= 8'h00;
            reg_file[24084] <= 8'h00;
            reg_file[24085] <= 8'h00;
            reg_file[24086] <= 8'h00;
            reg_file[24087] <= 8'h00;
            reg_file[24088] <= 8'h00;
            reg_file[24089] <= 8'h00;
            reg_file[24090] <= 8'h00;
            reg_file[24091] <= 8'h00;
            reg_file[24092] <= 8'h00;
            reg_file[24093] <= 8'h00;
            reg_file[24094] <= 8'h00;
            reg_file[24095] <= 8'h00;
            reg_file[24096] <= 8'h00;
            reg_file[24097] <= 8'h00;
            reg_file[24098] <= 8'h00;
            reg_file[24099] <= 8'h00;
            reg_file[24100] <= 8'h00;
            reg_file[24101] <= 8'h00;
            reg_file[24102] <= 8'h00;
            reg_file[24103] <= 8'h00;
            reg_file[24104] <= 8'h00;
            reg_file[24105] <= 8'h00;
            reg_file[24106] <= 8'h00;
            reg_file[24107] <= 8'h00;
            reg_file[24108] <= 8'h00;
            reg_file[24109] <= 8'h00;
            reg_file[24110] <= 8'h00;
            reg_file[24111] <= 8'h00;
            reg_file[24112] <= 8'h00;
            reg_file[24113] <= 8'h00;
            reg_file[24114] <= 8'h00;
            reg_file[24115] <= 8'h00;
            reg_file[24116] <= 8'h00;
            reg_file[24117] <= 8'h00;
            reg_file[24118] <= 8'h00;
            reg_file[24119] <= 8'h00;
            reg_file[24120] <= 8'h00;
            reg_file[24121] <= 8'h00;
            reg_file[24122] <= 8'h00;
            reg_file[24123] <= 8'h00;
            reg_file[24124] <= 8'h00;
            reg_file[24125] <= 8'h00;
            reg_file[24126] <= 8'h00;
            reg_file[24127] <= 8'h00;
            reg_file[24128] <= 8'h00;
            reg_file[24129] <= 8'h00;
            reg_file[24130] <= 8'h00;
            reg_file[24131] <= 8'h00;
            reg_file[24132] <= 8'h00;
            reg_file[24133] <= 8'h00;
            reg_file[24134] <= 8'h00;
            reg_file[24135] <= 8'h00;
            reg_file[24136] <= 8'h00;
            reg_file[24137] <= 8'h00;
            reg_file[24138] <= 8'h00;
            reg_file[24139] <= 8'h00;
            reg_file[24140] <= 8'h00;
            reg_file[24141] <= 8'h00;
            reg_file[24142] <= 8'h00;
            reg_file[24143] <= 8'h00;
            reg_file[24144] <= 8'h00;
            reg_file[24145] <= 8'h00;
            reg_file[24146] <= 8'h00;
            reg_file[24147] <= 8'h00;
            reg_file[24148] <= 8'h00;
            reg_file[24149] <= 8'h00;
            reg_file[24150] <= 8'h00;
            reg_file[24151] <= 8'h00;
            reg_file[24152] <= 8'h00;
            reg_file[24153] <= 8'h00;
            reg_file[24154] <= 8'h00;
            reg_file[24155] <= 8'h00;
            reg_file[24156] <= 8'h00;
            reg_file[24157] <= 8'h00;
            reg_file[24158] <= 8'h00;
            reg_file[24159] <= 8'h00;
            reg_file[24160] <= 8'h00;
            reg_file[24161] <= 8'h00;
            reg_file[24162] <= 8'h00;
            reg_file[24163] <= 8'h00;
            reg_file[24164] <= 8'h00;
            reg_file[24165] <= 8'h00;
            reg_file[24166] <= 8'h00;
            reg_file[24167] <= 8'h00;
            reg_file[24168] <= 8'h00;
            reg_file[24169] <= 8'h00;
            reg_file[24170] <= 8'h00;
            reg_file[24171] <= 8'h00;
            reg_file[24172] <= 8'h00;
            reg_file[24173] <= 8'h00;
            reg_file[24174] <= 8'h00;
            reg_file[24175] <= 8'h00;
            reg_file[24176] <= 8'h00;
            reg_file[24177] <= 8'h00;
            reg_file[24178] <= 8'h00;
            reg_file[24179] <= 8'h00;
            reg_file[24180] <= 8'h00;
            reg_file[24181] <= 8'h00;
            reg_file[24182] <= 8'h00;
            reg_file[24183] <= 8'h00;
            reg_file[24184] <= 8'h00;
            reg_file[24185] <= 8'h00;
            reg_file[24186] <= 8'h00;
            reg_file[24187] <= 8'h00;
            reg_file[24188] <= 8'h00;
            reg_file[24189] <= 8'h00;
            reg_file[24190] <= 8'h00;
            reg_file[24191] <= 8'h00;
            reg_file[24192] <= 8'h00;
            reg_file[24193] <= 8'h00;
            reg_file[24194] <= 8'h00;
            reg_file[24195] <= 8'h00;
            reg_file[24196] <= 8'h00;
            reg_file[24197] <= 8'h00;
            reg_file[24198] <= 8'h00;
            reg_file[24199] <= 8'h00;
            reg_file[24200] <= 8'h00;
            reg_file[24201] <= 8'h00;
            reg_file[24202] <= 8'h00;
            reg_file[24203] <= 8'h00;
            reg_file[24204] <= 8'h00;
            reg_file[24205] <= 8'h00;
            reg_file[24206] <= 8'h00;
            reg_file[24207] <= 8'h00;
            reg_file[24208] <= 8'h00;
            reg_file[24209] <= 8'h00;
            reg_file[24210] <= 8'h00;
            reg_file[24211] <= 8'h00;
            reg_file[24212] <= 8'h00;
            reg_file[24213] <= 8'h00;
            reg_file[24214] <= 8'h00;
            reg_file[24215] <= 8'h00;
            reg_file[24216] <= 8'h00;
            reg_file[24217] <= 8'h00;
            reg_file[24218] <= 8'h00;
            reg_file[24219] <= 8'h00;
            reg_file[24220] <= 8'h00;
            reg_file[24221] <= 8'h00;
            reg_file[24222] <= 8'h00;
            reg_file[24223] <= 8'h00;
            reg_file[24224] <= 8'h00;
            reg_file[24225] <= 8'h00;
            reg_file[24226] <= 8'h00;
            reg_file[24227] <= 8'h00;
            reg_file[24228] <= 8'h00;
            reg_file[24229] <= 8'h00;
            reg_file[24230] <= 8'h00;
            reg_file[24231] <= 8'h00;
            reg_file[24232] <= 8'h00;
            reg_file[24233] <= 8'h00;
            reg_file[24234] <= 8'h00;
            reg_file[24235] <= 8'h00;
            reg_file[24236] <= 8'h00;
            reg_file[24237] <= 8'h00;
            reg_file[24238] <= 8'h00;
            reg_file[24239] <= 8'h00;
            reg_file[24240] <= 8'h00;
            reg_file[24241] <= 8'h00;
            reg_file[24242] <= 8'h00;
            reg_file[24243] <= 8'h00;
            reg_file[24244] <= 8'h00;
            reg_file[24245] <= 8'h00;
            reg_file[24246] <= 8'h00;
            reg_file[24247] <= 8'h00;
            reg_file[24248] <= 8'h00;
            reg_file[24249] <= 8'h00;
            reg_file[24250] <= 8'h00;
            reg_file[24251] <= 8'h00;
            reg_file[24252] <= 8'h00;
            reg_file[24253] <= 8'h00;
            reg_file[24254] <= 8'h00;
            reg_file[24255] <= 8'h00;
            reg_file[24256] <= 8'h00;
            reg_file[24257] <= 8'h00;
            reg_file[24258] <= 8'h00;
            reg_file[24259] <= 8'h00;
            reg_file[24260] <= 8'h00;
            reg_file[24261] <= 8'h00;
            reg_file[24262] <= 8'h00;
            reg_file[24263] <= 8'h00;
            reg_file[24264] <= 8'h00;
            reg_file[24265] <= 8'h00;
            reg_file[24266] <= 8'h00;
            reg_file[24267] <= 8'h00;
            reg_file[24268] <= 8'h00;
            reg_file[24269] <= 8'h00;
            reg_file[24270] <= 8'h00;
            reg_file[24271] <= 8'h00;
            reg_file[24272] <= 8'h00;
            reg_file[24273] <= 8'h00;
            reg_file[24274] <= 8'h00;
            reg_file[24275] <= 8'h00;
            reg_file[24276] <= 8'h00;
            reg_file[24277] <= 8'h00;
            reg_file[24278] <= 8'h00;
            reg_file[24279] <= 8'h00;
            reg_file[24280] <= 8'h00;
            reg_file[24281] <= 8'h00;
            reg_file[24282] <= 8'h00;
            reg_file[24283] <= 8'h00;
            reg_file[24284] <= 8'h00;
            reg_file[24285] <= 8'h00;
            reg_file[24286] <= 8'h00;
            reg_file[24287] <= 8'h00;
            reg_file[24288] <= 8'h00;
            reg_file[24289] <= 8'h00;
            reg_file[24290] <= 8'h00;
            reg_file[24291] <= 8'h00;
            reg_file[24292] <= 8'h00;
            reg_file[24293] <= 8'h00;
            reg_file[24294] <= 8'h00;
            reg_file[24295] <= 8'h00;
            reg_file[24296] <= 8'h00;
            reg_file[24297] <= 8'h00;
            reg_file[24298] <= 8'h00;
            reg_file[24299] <= 8'h00;
            reg_file[24300] <= 8'h00;
            reg_file[24301] <= 8'h00;
            reg_file[24302] <= 8'h00;
            reg_file[24303] <= 8'h00;
            reg_file[24304] <= 8'h00;
            reg_file[24305] <= 8'h00;
            reg_file[24306] <= 8'h00;
            reg_file[24307] <= 8'h00;
            reg_file[24308] <= 8'h00;
            reg_file[24309] <= 8'h00;
            reg_file[24310] <= 8'h00;
            reg_file[24311] <= 8'h00;
            reg_file[24312] <= 8'h00;
            reg_file[24313] <= 8'h00;
            reg_file[24314] <= 8'h00;
            reg_file[24315] <= 8'h00;
            reg_file[24316] <= 8'h00;
            reg_file[24317] <= 8'h00;
            reg_file[24318] <= 8'h00;
            reg_file[24319] <= 8'h00;
            reg_file[24320] <= 8'h00;
            reg_file[24321] <= 8'h00;
            reg_file[24322] <= 8'h00;
            reg_file[24323] <= 8'h00;
            reg_file[24324] <= 8'h00;
            reg_file[24325] <= 8'h00;
            reg_file[24326] <= 8'h00;
            reg_file[24327] <= 8'h00;
            reg_file[24328] <= 8'h00;
            reg_file[24329] <= 8'h00;
            reg_file[24330] <= 8'h00;
            reg_file[24331] <= 8'h00;
            reg_file[24332] <= 8'h00;
            reg_file[24333] <= 8'h00;
            reg_file[24334] <= 8'h00;
            reg_file[24335] <= 8'h00;
            reg_file[24336] <= 8'h00;
            reg_file[24337] <= 8'h00;
            reg_file[24338] <= 8'h00;
            reg_file[24339] <= 8'h00;
            reg_file[24340] <= 8'h00;
            reg_file[24341] <= 8'h00;
            reg_file[24342] <= 8'h00;
            reg_file[24343] <= 8'h00;
            reg_file[24344] <= 8'h00;
            reg_file[24345] <= 8'h00;
            reg_file[24346] <= 8'h00;
            reg_file[24347] <= 8'h00;
            reg_file[24348] <= 8'h00;
            reg_file[24349] <= 8'h00;
            reg_file[24350] <= 8'h00;
            reg_file[24351] <= 8'h00;
            reg_file[24352] <= 8'h00;
            reg_file[24353] <= 8'h00;
            reg_file[24354] <= 8'h00;
            reg_file[24355] <= 8'h00;
            reg_file[24356] <= 8'h00;
            reg_file[24357] <= 8'h00;
            reg_file[24358] <= 8'h00;
            reg_file[24359] <= 8'h00;
            reg_file[24360] <= 8'h00;
            reg_file[24361] <= 8'h00;
            reg_file[24362] <= 8'h00;
            reg_file[24363] <= 8'h00;
            reg_file[24364] <= 8'h00;
            reg_file[24365] <= 8'h00;
            reg_file[24366] <= 8'h00;
            reg_file[24367] <= 8'h00;
            reg_file[24368] <= 8'h00;
            reg_file[24369] <= 8'h00;
            reg_file[24370] <= 8'h00;
            reg_file[24371] <= 8'h00;
            reg_file[24372] <= 8'h00;
            reg_file[24373] <= 8'h00;
            reg_file[24374] <= 8'h00;
            reg_file[24375] <= 8'h00;
            reg_file[24376] <= 8'h00;
            reg_file[24377] <= 8'h00;
            reg_file[24378] <= 8'h00;
            reg_file[24379] <= 8'h00;
            reg_file[24380] <= 8'h00;
            reg_file[24381] <= 8'h00;
            reg_file[24382] <= 8'h00;
            reg_file[24383] <= 8'h00;
            reg_file[24384] <= 8'h00;
            reg_file[24385] <= 8'h00;
            reg_file[24386] <= 8'h00;
            reg_file[24387] <= 8'h00;
            reg_file[24388] <= 8'h00;
            reg_file[24389] <= 8'h00;
            reg_file[24390] <= 8'h00;
            reg_file[24391] <= 8'h00;
            reg_file[24392] <= 8'h00;
            reg_file[24393] <= 8'h00;
            reg_file[24394] <= 8'h00;
            reg_file[24395] <= 8'h00;
            reg_file[24396] <= 8'h00;
            reg_file[24397] <= 8'h00;
            reg_file[24398] <= 8'h00;
            reg_file[24399] <= 8'h00;
            reg_file[24400] <= 8'h00;
            reg_file[24401] <= 8'h00;
            reg_file[24402] <= 8'h00;
            reg_file[24403] <= 8'h00;
            reg_file[24404] <= 8'h00;
            reg_file[24405] <= 8'h00;
            reg_file[24406] <= 8'h00;
            reg_file[24407] <= 8'h00;
            reg_file[24408] <= 8'h00;
            reg_file[24409] <= 8'h00;
            reg_file[24410] <= 8'h00;
            reg_file[24411] <= 8'h00;
            reg_file[24412] <= 8'h00;
            reg_file[24413] <= 8'h00;
            reg_file[24414] <= 8'h00;
            reg_file[24415] <= 8'h00;
            reg_file[24416] <= 8'h00;
            reg_file[24417] <= 8'h00;
            reg_file[24418] <= 8'h00;
            reg_file[24419] <= 8'h00;
            reg_file[24420] <= 8'h00;
            reg_file[24421] <= 8'h00;
            reg_file[24422] <= 8'h00;
            reg_file[24423] <= 8'h00;
            reg_file[24424] <= 8'h00;
            reg_file[24425] <= 8'h00;
            reg_file[24426] <= 8'h00;
            reg_file[24427] <= 8'h00;
            reg_file[24428] <= 8'h00;
            reg_file[24429] <= 8'h00;
            reg_file[24430] <= 8'h00;
            reg_file[24431] <= 8'h00;
            reg_file[24432] <= 8'h00;
            reg_file[24433] <= 8'h00;
            reg_file[24434] <= 8'h00;
            reg_file[24435] <= 8'h00;
            reg_file[24436] <= 8'h00;
            reg_file[24437] <= 8'h00;
            reg_file[24438] <= 8'h00;
            reg_file[24439] <= 8'h00;
            reg_file[24440] <= 8'h00;
            reg_file[24441] <= 8'h00;
            reg_file[24442] <= 8'h00;
            reg_file[24443] <= 8'h00;
            reg_file[24444] <= 8'h00;
            reg_file[24445] <= 8'h00;
            reg_file[24446] <= 8'h00;
            reg_file[24447] <= 8'h00;
            reg_file[24448] <= 8'h00;
            reg_file[24449] <= 8'h00;
            reg_file[24450] <= 8'h00;
            reg_file[24451] <= 8'h00;
            reg_file[24452] <= 8'h00;
            reg_file[24453] <= 8'h00;
            reg_file[24454] <= 8'h00;
            reg_file[24455] <= 8'h00;
            reg_file[24456] <= 8'h00;
            reg_file[24457] <= 8'h00;
            reg_file[24458] <= 8'h00;
            reg_file[24459] <= 8'h00;
            reg_file[24460] <= 8'h00;
            reg_file[24461] <= 8'h00;
            reg_file[24462] <= 8'h00;
            reg_file[24463] <= 8'h00;
            reg_file[24464] <= 8'h00;
            reg_file[24465] <= 8'h00;
            reg_file[24466] <= 8'h00;
            reg_file[24467] <= 8'h00;
            reg_file[24468] <= 8'h00;
            reg_file[24469] <= 8'h00;
            reg_file[24470] <= 8'h00;
            reg_file[24471] <= 8'h00;
            reg_file[24472] <= 8'h00;
            reg_file[24473] <= 8'h00;
            reg_file[24474] <= 8'h00;
            reg_file[24475] <= 8'h00;
            reg_file[24476] <= 8'h00;
            reg_file[24477] <= 8'h00;
            reg_file[24478] <= 8'h00;
            reg_file[24479] <= 8'h00;
            reg_file[24480] <= 8'h00;
            reg_file[24481] <= 8'h00;
            reg_file[24482] <= 8'h00;
            reg_file[24483] <= 8'h00;
            reg_file[24484] <= 8'h00;
            reg_file[24485] <= 8'h00;
            reg_file[24486] <= 8'h00;
            reg_file[24487] <= 8'h00;
            reg_file[24488] <= 8'h00;
            reg_file[24489] <= 8'h00;
            reg_file[24490] <= 8'h00;
            reg_file[24491] <= 8'h00;
            reg_file[24492] <= 8'h00;
            reg_file[24493] <= 8'h00;
            reg_file[24494] <= 8'h00;
            reg_file[24495] <= 8'h00;
            reg_file[24496] <= 8'h00;
            reg_file[24497] <= 8'h00;
            reg_file[24498] <= 8'h00;
            reg_file[24499] <= 8'h00;
            reg_file[24500] <= 8'h00;
            reg_file[24501] <= 8'h00;
            reg_file[24502] <= 8'h00;
            reg_file[24503] <= 8'h00;
            reg_file[24504] <= 8'h00;
            reg_file[24505] <= 8'h00;
            reg_file[24506] <= 8'h00;
            reg_file[24507] <= 8'h00;
            reg_file[24508] <= 8'h00;
            reg_file[24509] <= 8'h00;
            reg_file[24510] <= 8'h00;
            reg_file[24511] <= 8'h00;
            reg_file[24512] <= 8'h00;
            reg_file[24513] <= 8'h00;
            reg_file[24514] <= 8'h00;
            reg_file[24515] <= 8'h00;
            reg_file[24516] <= 8'h00;
            reg_file[24517] <= 8'h00;
            reg_file[24518] <= 8'h00;
            reg_file[24519] <= 8'h00;
            reg_file[24520] <= 8'h00;
            reg_file[24521] <= 8'h00;
            reg_file[24522] <= 8'h00;
            reg_file[24523] <= 8'h00;
            reg_file[24524] <= 8'h00;
            reg_file[24525] <= 8'h00;
            reg_file[24526] <= 8'h00;
            reg_file[24527] <= 8'h00;
            reg_file[24528] <= 8'h00;
            reg_file[24529] <= 8'h00;
            reg_file[24530] <= 8'h00;
            reg_file[24531] <= 8'h00;
            reg_file[24532] <= 8'h00;
            reg_file[24533] <= 8'h00;
            reg_file[24534] <= 8'h00;
            reg_file[24535] <= 8'h00;
            reg_file[24536] <= 8'h00;
            reg_file[24537] <= 8'h00;
            reg_file[24538] <= 8'h00;
            reg_file[24539] <= 8'h00;
            reg_file[24540] <= 8'h00;
            reg_file[24541] <= 8'h00;
            reg_file[24542] <= 8'h00;
            reg_file[24543] <= 8'h00;
            reg_file[24544] <= 8'h00;
            reg_file[24545] <= 8'h00;
            reg_file[24546] <= 8'h00;
            reg_file[24547] <= 8'h00;
            reg_file[24548] <= 8'h00;
            reg_file[24549] <= 8'h00;
            reg_file[24550] <= 8'h00;
            reg_file[24551] <= 8'h00;
            reg_file[24552] <= 8'h00;
            reg_file[24553] <= 8'h00;
            reg_file[24554] <= 8'h00;
            reg_file[24555] <= 8'h00;
            reg_file[24556] <= 8'h00;
            reg_file[24557] <= 8'h00;
            reg_file[24558] <= 8'h00;
            reg_file[24559] <= 8'h00;
            reg_file[24560] <= 8'h00;
            reg_file[24561] <= 8'h00;
            reg_file[24562] <= 8'h00;
            reg_file[24563] <= 8'h00;
            reg_file[24564] <= 8'h00;
            reg_file[24565] <= 8'h00;
            reg_file[24566] <= 8'h00;
            reg_file[24567] <= 8'h00;
            reg_file[24568] <= 8'h00;
            reg_file[24569] <= 8'h00;
            reg_file[24570] <= 8'h00;
            reg_file[24571] <= 8'h00;
            reg_file[24572] <= 8'h00;
            reg_file[24573] <= 8'h00;
            reg_file[24574] <= 8'h00;
            reg_file[24575] <= 8'h00;
            reg_file[24576] <= 8'h00;
            reg_file[24577] <= 8'h00;
            reg_file[24578] <= 8'h00;
            reg_file[24579] <= 8'h00;
            reg_file[24580] <= 8'h00;
            reg_file[24581] <= 8'h00;
            reg_file[24582] <= 8'h00;
            reg_file[24583] <= 8'h00;
            reg_file[24584] <= 8'h00;
            reg_file[24585] <= 8'h00;
            reg_file[24586] <= 8'h00;
            reg_file[24587] <= 8'h00;
            reg_file[24588] <= 8'h00;
            reg_file[24589] <= 8'h00;
            reg_file[24590] <= 8'h00;
            reg_file[24591] <= 8'h00;
            reg_file[24592] <= 8'h00;
            reg_file[24593] <= 8'h00;
            reg_file[24594] <= 8'h00;
            reg_file[24595] <= 8'h00;
            reg_file[24596] <= 8'h00;
            reg_file[24597] <= 8'h00;
            reg_file[24598] <= 8'h00;
            reg_file[24599] <= 8'h00;
            reg_file[24600] <= 8'h00;
            reg_file[24601] <= 8'h00;
            reg_file[24602] <= 8'h00;
            reg_file[24603] <= 8'h00;
            reg_file[24604] <= 8'h00;
            reg_file[24605] <= 8'h00;
            reg_file[24606] <= 8'h00;
            reg_file[24607] <= 8'h00;
            reg_file[24608] <= 8'h00;
            reg_file[24609] <= 8'h00;
            reg_file[24610] <= 8'h00;
            reg_file[24611] <= 8'h00;
            reg_file[24612] <= 8'h00;
            reg_file[24613] <= 8'h00;
            reg_file[24614] <= 8'h00;
            reg_file[24615] <= 8'h00;
            reg_file[24616] <= 8'h00;
            reg_file[24617] <= 8'h00;
            reg_file[24618] <= 8'h00;
            reg_file[24619] <= 8'h00;
            reg_file[24620] <= 8'h00;
            reg_file[24621] <= 8'h00;
            reg_file[24622] <= 8'h00;
            reg_file[24623] <= 8'h00;
            reg_file[24624] <= 8'h00;
            reg_file[24625] <= 8'h00;
            reg_file[24626] <= 8'h00;
            reg_file[24627] <= 8'h00;
            reg_file[24628] <= 8'h00;
            reg_file[24629] <= 8'h00;
            reg_file[24630] <= 8'h00;
            reg_file[24631] <= 8'h00;
            reg_file[24632] <= 8'h00;
            reg_file[24633] <= 8'h00;
            reg_file[24634] <= 8'h00;
            reg_file[24635] <= 8'h00;
            reg_file[24636] <= 8'h00;
            reg_file[24637] <= 8'h00;
            reg_file[24638] <= 8'h00;
            reg_file[24639] <= 8'h00;
            reg_file[24640] <= 8'h00;
            reg_file[24641] <= 8'h00;
            reg_file[24642] <= 8'h00;
            reg_file[24643] <= 8'h00;
            reg_file[24644] <= 8'h00;
            reg_file[24645] <= 8'h00;
            reg_file[24646] <= 8'h00;
            reg_file[24647] <= 8'h00;
            reg_file[24648] <= 8'h00;
            reg_file[24649] <= 8'h00;
            reg_file[24650] <= 8'h00;
            reg_file[24651] <= 8'h00;
            reg_file[24652] <= 8'h00;
            reg_file[24653] <= 8'h00;
            reg_file[24654] <= 8'h00;
            reg_file[24655] <= 8'h00;
            reg_file[24656] <= 8'h00;
            reg_file[24657] <= 8'h00;
            reg_file[24658] <= 8'h00;
            reg_file[24659] <= 8'h00;
            reg_file[24660] <= 8'h00;
            reg_file[24661] <= 8'h00;
            reg_file[24662] <= 8'h00;
            reg_file[24663] <= 8'h00;
            reg_file[24664] <= 8'h00;
            reg_file[24665] <= 8'h00;
            reg_file[24666] <= 8'h00;
            reg_file[24667] <= 8'h00;
            reg_file[24668] <= 8'h00;
            reg_file[24669] <= 8'h00;
            reg_file[24670] <= 8'h00;
            reg_file[24671] <= 8'h00;
            reg_file[24672] <= 8'h00;
            reg_file[24673] <= 8'h00;
            reg_file[24674] <= 8'h00;
            reg_file[24675] <= 8'h00;
            reg_file[24676] <= 8'h00;
            reg_file[24677] <= 8'h00;
            reg_file[24678] <= 8'h00;
            reg_file[24679] <= 8'h00;
            reg_file[24680] <= 8'h00;
            reg_file[24681] <= 8'h00;
            reg_file[24682] <= 8'h00;
            reg_file[24683] <= 8'h00;
            reg_file[24684] <= 8'h00;
            reg_file[24685] <= 8'h00;
            reg_file[24686] <= 8'h00;
            reg_file[24687] <= 8'h00;
            reg_file[24688] <= 8'h00;
            reg_file[24689] <= 8'h00;
            reg_file[24690] <= 8'h00;
            reg_file[24691] <= 8'h00;
            reg_file[24692] <= 8'h00;
            reg_file[24693] <= 8'h00;
            reg_file[24694] <= 8'h00;
            reg_file[24695] <= 8'h00;
            reg_file[24696] <= 8'h00;
            reg_file[24697] <= 8'h00;
            reg_file[24698] <= 8'h00;
            reg_file[24699] <= 8'h00;
            reg_file[24700] <= 8'h00;
            reg_file[24701] <= 8'h00;
            reg_file[24702] <= 8'h00;
            reg_file[24703] <= 8'h00;
            reg_file[24704] <= 8'h00;
            reg_file[24705] <= 8'h00;
            reg_file[24706] <= 8'h00;
            reg_file[24707] <= 8'h00;
            reg_file[24708] <= 8'h00;
            reg_file[24709] <= 8'h00;
            reg_file[24710] <= 8'h00;
            reg_file[24711] <= 8'h00;
            reg_file[24712] <= 8'h00;
            reg_file[24713] <= 8'h00;
            reg_file[24714] <= 8'h00;
            reg_file[24715] <= 8'h00;
            reg_file[24716] <= 8'h00;
            reg_file[24717] <= 8'h00;
            reg_file[24718] <= 8'h00;
            reg_file[24719] <= 8'h00;
            reg_file[24720] <= 8'h00;
            reg_file[24721] <= 8'h00;
            reg_file[24722] <= 8'h00;
            reg_file[24723] <= 8'h00;
            reg_file[24724] <= 8'h00;
            reg_file[24725] <= 8'h00;
            reg_file[24726] <= 8'h00;
            reg_file[24727] <= 8'h00;
            reg_file[24728] <= 8'h00;
            reg_file[24729] <= 8'h00;
            reg_file[24730] <= 8'h00;
            reg_file[24731] <= 8'h00;
            reg_file[24732] <= 8'h00;
            reg_file[24733] <= 8'h00;
            reg_file[24734] <= 8'h00;
            reg_file[24735] <= 8'h00;
            reg_file[24736] <= 8'h00;
            reg_file[24737] <= 8'h00;
            reg_file[24738] <= 8'h00;
            reg_file[24739] <= 8'h00;
            reg_file[24740] <= 8'h00;
            reg_file[24741] <= 8'h00;
            reg_file[24742] <= 8'h00;
            reg_file[24743] <= 8'h00;
            reg_file[24744] <= 8'h00;
            reg_file[24745] <= 8'h00;
            reg_file[24746] <= 8'h00;
            reg_file[24747] <= 8'h00;
            reg_file[24748] <= 8'h00;
            reg_file[24749] <= 8'h00;
            reg_file[24750] <= 8'h00;
            reg_file[24751] <= 8'h00;
            reg_file[24752] <= 8'h00;
            reg_file[24753] <= 8'h00;
            reg_file[24754] <= 8'h00;
            reg_file[24755] <= 8'h00;
            reg_file[24756] <= 8'h00;
            reg_file[24757] <= 8'h00;
            reg_file[24758] <= 8'h00;
            reg_file[24759] <= 8'h00;
            reg_file[24760] <= 8'h00;
            reg_file[24761] <= 8'h00;
            reg_file[24762] <= 8'h00;
            reg_file[24763] <= 8'h00;
            reg_file[24764] <= 8'h00;
            reg_file[24765] <= 8'h00;
            reg_file[24766] <= 8'h00;
            reg_file[24767] <= 8'h00;
            reg_file[24768] <= 8'h00;
            reg_file[24769] <= 8'h00;
            reg_file[24770] <= 8'h00;
            reg_file[24771] <= 8'h00;
            reg_file[24772] <= 8'h00;
            reg_file[24773] <= 8'h00;
            reg_file[24774] <= 8'h00;
            reg_file[24775] <= 8'h00;
            reg_file[24776] <= 8'h00;
            reg_file[24777] <= 8'h00;
            reg_file[24778] <= 8'h00;
            reg_file[24779] <= 8'h00;
            reg_file[24780] <= 8'h00;
            reg_file[24781] <= 8'h00;
            reg_file[24782] <= 8'h00;
            reg_file[24783] <= 8'h00;
            reg_file[24784] <= 8'h00;
            reg_file[24785] <= 8'h00;
            reg_file[24786] <= 8'h00;
            reg_file[24787] <= 8'h00;
            reg_file[24788] <= 8'h00;
            reg_file[24789] <= 8'h00;
            reg_file[24790] <= 8'h00;
            reg_file[24791] <= 8'h00;
            reg_file[24792] <= 8'h00;
            reg_file[24793] <= 8'h00;
            reg_file[24794] <= 8'h00;
            reg_file[24795] <= 8'h00;
            reg_file[24796] <= 8'h00;
            reg_file[24797] <= 8'h00;
            reg_file[24798] <= 8'h00;
            reg_file[24799] <= 8'h00;
            reg_file[24800] <= 8'h00;
            reg_file[24801] <= 8'h00;
            reg_file[24802] <= 8'h00;
            reg_file[24803] <= 8'h00;
            reg_file[24804] <= 8'h00;
            reg_file[24805] <= 8'h00;
            reg_file[24806] <= 8'h00;
            reg_file[24807] <= 8'h00;
            reg_file[24808] <= 8'h00;
            reg_file[24809] <= 8'h00;
            reg_file[24810] <= 8'h00;
            reg_file[24811] <= 8'h00;
            reg_file[24812] <= 8'h00;
            reg_file[24813] <= 8'h00;
            reg_file[24814] <= 8'h00;
            reg_file[24815] <= 8'h00;
            reg_file[24816] <= 8'h00;
            reg_file[24817] <= 8'h00;
            reg_file[24818] <= 8'h00;
            reg_file[24819] <= 8'h00;
            reg_file[24820] <= 8'h00;
            reg_file[24821] <= 8'h00;
            reg_file[24822] <= 8'h00;
            reg_file[24823] <= 8'h00;
            reg_file[24824] <= 8'h00;
            reg_file[24825] <= 8'h00;
            reg_file[24826] <= 8'h00;
            reg_file[24827] <= 8'h00;
            reg_file[24828] <= 8'h00;
            reg_file[24829] <= 8'h00;
            reg_file[24830] <= 8'h00;
            reg_file[24831] <= 8'h00;
            reg_file[24832] <= 8'h00;
            reg_file[24833] <= 8'h00;
            reg_file[24834] <= 8'h00;
            reg_file[24835] <= 8'h00;
            reg_file[24836] <= 8'h00;
            reg_file[24837] <= 8'h00;
            reg_file[24838] <= 8'h00;
            reg_file[24839] <= 8'h00;
            reg_file[24840] <= 8'h00;
            reg_file[24841] <= 8'h00;
            reg_file[24842] <= 8'h00;
            reg_file[24843] <= 8'h00;
            reg_file[24844] <= 8'h00;
            reg_file[24845] <= 8'h00;
            reg_file[24846] <= 8'h00;
            reg_file[24847] <= 8'h00;
            reg_file[24848] <= 8'h00;
            reg_file[24849] <= 8'h00;
            reg_file[24850] <= 8'h00;
            reg_file[24851] <= 8'h00;
            reg_file[24852] <= 8'h00;
            reg_file[24853] <= 8'h00;
            reg_file[24854] <= 8'h00;
            reg_file[24855] <= 8'h00;
            reg_file[24856] <= 8'h00;
            reg_file[24857] <= 8'h00;
            reg_file[24858] <= 8'h00;
            reg_file[24859] <= 8'h00;
            reg_file[24860] <= 8'h00;
            reg_file[24861] <= 8'h00;
            reg_file[24862] <= 8'h00;
            reg_file[24863] <= 8'h00;
            reg_file[24864] <= 8'h00;
            reg_file[24865] <= 8'h00;
            reg_file[24866] <= 8'h00;
            reg_file[24867] <= 8'h00;
            reg_file[24868] <= 8'h00;
            reg_file[24869] <= 8'h00;
            reg_file[24870] <= 8'h00;
            reg_file[24871] <= 8'h00;
            reg_file[24872] <= 8'h00;
            reg_file[24873] <= 8'h00;
            reg_file[24874] <= 8'h00;
            reg_file[24875] <= 8'h00;
            reg_file[24876] <= 8'h00;
            reg_file[24877] <= 8'h00;
            reg_file[24878] <= 8'h00;
            reg_file[24879] <= 8'h00;
            reg_file[24880] <= 8'h00;
            reg_file[24881] <= 8'h00;
            reg_file[24882] <= 8'h00;
            reg_file[24883] <= 8'h00;
            reg_file[24884] <= 8'h00;
            reg_file[24885] <= 8'h00;
            reg_file[24886] <= 8'h00;
            reg_file[24887] <= 8'h00;
            reg_file[24888] <= 8'h00;
            reg_file[24889] <= 8'h00;
            reg_file[24890] <= 8'h00;
            reg_file[24891] <= 8'h00;
            reg_file[24892] <= 8'h00;
            reg_file[24893] <= 8'h00;
            reg_file[24894] <= 8'h00;
            reg_file[24895] <= 8'h00;
            reg_file[24896] <= 8'h00;
            reg_file[24897] <= 8'h00;
            reg_file[24898] <= 8'h00;
            reg_file[24899] <= 8'h00;
            reg_file[24900] <= 8'h00;
            reg_file[24901] <= 8'h00;
            reg_file[24902] <= 8'h00;
            reg_file[24903] <= 8'h00;
            reg_file[24904] <= 8'h00;
            reg_file[24905] <= 8'h00;
            reg_file[24906] <= 8'h00;
            reg_file[24907] <= 8'h00;
            reg_file[24908] <= 8'h00;
            reg_file[24909] <= 8'h00;
            reg_file[24910] <= 8'h00;
            reg_file[24911] <= 8'h00;
            reg_file[24912] <= 8'h00;
            reg_file[24913] <= 8'h00;
            reg_file[24914] <= 8'h00;
            reg_file[24915] <= 8'h00;
            reg_file[24916] <= 8'h00;
            reg_file[24917] <= 8'h00;
            reg_file[24918] <= 8'h00;
            reg_file[24919] <= 8'h00;
            reg_file[24920] <= 8'h00;
            reg_file[24921] <= 8'h00;
            reg_file[24922] <= 8'h00;
            reg_file[24923] <= 8'h00;
            reg_file[24924] <= 8'h00;
            reg_file[24925] <= 8'h00;
            reg_file[24926] <= 8'h00;
            reg_file[24927] <= 8'h00;
            reg_file[24928] <= 8'h00;
            reg_file[24929] <= 8'h00;
            reg_file[24930] <= 8'h00;
            reg_file[24931] <= 8'h00;
            reg_file[24932] <= 8'h00;
            reg_file[24933] <= 8'h00;
            reg_file[24934] <= 8'h00;
            reg_file[24935] <= 8'h00;
            reg_file[24936] <= 8'h00;
            reg_file[24937] <= 8'h00;
            reg_file[24938] <= 8'h00;
            reg_file[24939] <= 8'h00;
            reg_file[24940] <= 8'h00;
            reg_file[24941] <= 8'h00;
            reg_file[24942] <= 8'h00;
            reg_file[24943] <= 8'h00;
            reg_file[24944] <= 8'h00;
            reg_file[24945] <= 8'h00;
            reg_file[24946] <= 8'h00;
            reg_file[24947] <= 8'h00;
            reg_file[24948] <= 8'h00;
            reg_file[24949] <= 8'h00;
            reg_file[24950] <= 8'h00;
            reg_file[24951] <= 8'h00;
            reg_file[24952] <= 8'h00;
            reg_file[24953] <= 8'h00;
            reg_file[24954] <= 8'h00;
            reg_file[24955] <= 8'h00;
            reg_file[24956] <= 8'h00;
            reg_file[24957] <= 8'h00;
            reg_file[24958] <= 8'h00;
            reg_file[24959] <= 8'h00;
            reg_file[24960] <= 8'h00;
            reg_file[24961] <= 8'h00;
            reg_file[24962] <= 8'h00;
            reg_file[24963] <= 8'h00;
            reg_file[24964] <= 8'h00;
            reg_file[24965] <= 8'h00;
            reg_file[24966] <= 8'h00;
            reg_file[24967] <= 8'h00;
            reg_file[24968] <= 8'h00;
            reg_file[24969] <= 8'h00;
            reg_file[24970] <= 8'h00;
            reg_file[24971] <= 8'h00;
            reg_file[24972] <= 8'h00;
            reg_file[24973] <= 8'h00;
            reg_file[24974] <= 8'h00;
            reg_file[24975] <= 8'h00;
            reg_file[24976] <= 8'h00;
            reg_file[24977] <= 8'h00;
            reg_file[24978] <= 8'h00;
            reg_file[24979] <= 8'h00;
            reg_file[24980] <= 8'h00;
            reg_file[24981] <= 8'h00;
            reg_file[24982] <= 8'h00;
            reg_file[24983] <= 8'h00;
            reg_file[24984] <= 8'h00;
            reg_file[24985] <= 8'h00;
            reg_file[24986] <= 8'h00;
            reg_file[24987] <= 8'h00;
            reg_file[24988] <= 8'h00;
            reg_file[24989] <= 8'h00;
            reg_file[24990] <= 8'h00;
            reg_file[24991] <= 8'h00;
            reg_file[24992] <= 8'h00;
            reg_file[24993] <= 8'h00;
            reg_file[24994] <= 8'h00;
            reg_file[24995] <= 8'h00;
            reg_file[24996] <= 8'h00;
            reg_file[24997] <= 8'h00;
            reg_file[24998] <= 8'h00;
            reg_file[24999] <= 8'h00;
            reg_file[25000] <= 8'h00;
            reg_file[25001] <= 8'h00;
            reg_file[25002] <= 8'h00;
            reg_file[25003] <= 8'h00;
            reg_file[25004] <= 8'h00;
            reg_file[25005] <= 8'h00;
            reg_file[25006] <= 8'h00;
            reg_file[25007] <= 8'h00;
            reg_file[25008] <= 8'h00;
            reg_file[25009] <= 8'h00;
            reg_file[25010] <= 8'h00;
            reg_file[25011] <= 8'h00;
            reg_file[25012] <= 8'h00;
            reg_file[25013] <= 8'h00;
            reg_file[25014] <= 8'h00;
            reg_file[25015] <= 8'h00;
            reg_file[25016] <= 8'h00;
            reg_file[25017] <= 8'h00;
            reg_file[25018] <= 8'h00;
            reg_file[25019] <= 8'h00;
            reg_file[25020] <= 8'h00;
            reg_file[25021] <= 8'h00;
            reg_file[25022] <= 8'h00;
            reg_file[25023] <= 8'h00;
            reg_file[25024] <= 8'h00;
            reg_file[25025] <= 8'h00;
            reg_file[25026] <= 8'h00;
            reg_file[25027] <= 8'h00;
            reg_file[25028] <= 8'h00;
            reg_file[25029] <= 8'h00;
            reg_file[25030] <= 8'h00;
            reg_file[25031] <= 8'h00;
            reg_file[25032] <= 8'h00;
            reg_file[25033] <= 8'h00;
            reg_file[25034] <= 8'h00;
            reg_file[25035] <= 8'h00;
            reg_file[25036] <= 8'h00;
            reg_file[25037] <= 8'h00;
            reg_file[25038] <= 8'h00;
            reg_file[25039] <= 8'h00;
            reg_file[25040] <= 8'h00;
            reg_file[25041] <= 8'h00;
            reg_file[25042] <= 8'h00;
            reg_file[25043] <= 8'h00;
            reg_file[25044] <= 8'h00;
            reg_file[25045] <= 8'h00;
            reg_file[25046] <= 8'h00;
            reg_file[25047] <= 8'h00;
            reg_file[25048] <= 8'h00;
            reg_file[25049] <= 8'h00;
            reg_file[25050] <= 8'h00;
            reg_file[25051] <= 8'h00;
            reg_file[25052] <= 8'h00;
            reg_file[25053] <= 8'h00;
            reg_file[25054] <= 8'h00;
            reg_file[25055] <= 8'h00;
            reg_file[25056] <= 8'h00;
            reg_file[25057] <= 8'h00;
            reg_file[25058] <= 8'h00;
            reg_file[25059] <= 8'h00;
            reg_file[25060] <= 8'h00;
            reg_file[25061] <= 8'h00;
            reg_file[25062] <= 8'h00;
            reg_file[25063] <= 8'h00;
            reg_file[25064] <= 8'h00;
            reg_file[25065] <= 8'h00;
            reg_file[25066] <= 8'h00;
            reg_file[25067] <= 8'h00;
            reg_file[25068] <= 8'h00;
            reg_file[25069] <= 8'h00;
            reg_file[25070] <= 8'h00;
            reg_file[25071] <= 8'h00;
            reg_file[25072] <= 8'h00;
            reg_file[25073] <= 8'h00;
            reg_file[25074] <= 8'h00;
            reg_file[25075] <= 8'h00;
            reg_file[25076] <= 8'h00;
            reg_file[25077] <= 8'h00;
            reg_file[25078] <= 8'h00;
            reg_file[25079] <= 8'h00;
            reg_file[25080] <= 8'h00;
            reg_file[25081] <= 8'h00;
            reg_file[25082] <= 8'h00;
            reg_file[25083] <= 8'h00;
            reg_file[25084] <= 8'h00;
            reg_file[25085] <= 8'h00;
            reg_file[25086] <= 8'h00;
            reg_file[25087] <= 8'h00;
            reg_file[25088] <= 8'h00;
            reg_file[25089] <= 8'h00;
            reg_file[25090] <= 8'h00;
            reg_file[25091] <= 8'h00;
            reg_file[25092] <= 8'h00;
            reg_file[25093] <= 8'h00;
            reg_file[25094] <= 8'h00;
            reg_file[25095] <= 8'h00;
            reg_file[25096] <= 8'h00;
            reg_file[25097] <= 8'h00;
            reg_file[25098] <= 8'h00;
            reg_file[25099] <= 8'h00;
            reg_file[25100] <= 8'h00;
            reg_file[25101] <= 8'h00;
            reg_file[25102] <= 8'h00;
            reg_file[25103] <= 8'h00;
            reg_file[25104] <= 8'h00;
            reg_file[25105] <= 8'h00;
            reg_file[25106] <= 8'h00;
            reg_file[25107] <= 8'h00;
            reg_file[25108] <= 8'h00;
            reg_file[25109] <= 8'h00;
            reg_file[25110] <= 8'h00;
            reg_file[25111] <= 8'h00;
            reg_file[25112] <= 8'h00;
            reg_file[25113] <= 8'h00;
            reg_file[25114] <= 8'h00;
            reg_file[25115] <= 8'h00;
            reg_file[25116] <= 8'h00;
            reg_file[25117] <= 8'h00;
            reg_file[25118] <= 8'h00;
            reg_file[25119] <= 8'h00;
            reg_file[25120] <= 8'h00;
            reg_file[25121] <= 8'h00;
            reg_file[25122] <= 8'h00;
            reg_file[25123] <= 8'h00;
            reg_file[25124] <= 8'h00;
            reg_file[25125] <= 8'h00;
            reg_file[25126] <= 8'h00;
            reg_file[25127] <= 8'h00;
            reg_file[25128] <= 8'h00;
            reg_file[25129] <= 8'h00;
            reg_file[25130] <= 8'h00;
            reg_file[25131] <= 8'h00;
            reg_file[25132] <= 8'h00;
            reg_file[25133] <= 8'h00;
            reg_file[25134] <= 8'h00;
            reg_file[25135] <= 8'h00;
            reg_file[25136] <= 8'h00;
            reg_file[25137] <= 8'h00;
            reg_file[25138] <= 8'h00;
            reg_file[25139] <= 8'h00;
            reg_file[25140] <= 8'h00;
            reg_file[25141] <= 8'h00;
            reg_file[25142] <= 8'h00;
            reg_file[25143] <= 8'h00;
            reg_file[25144] <= 8'h00;
            reg_file[25145] <= 8'h00;
            reg_file[25146] <= 8'h00;
            reg_file[25147] <= 8'h00;
            reg_file[25148] <= 8'h00;
            reg_file[25149] <= 8'h00;
            reg_file[25150] <= 8'h00;
            reg_file[25151] <= 8'h00;
            reg_file[25152] <= 8'h00;
            reg_file[25153] <= 8'h00;
            reg_file[25154] <= 8'h00;
            reg_file[25155] <= 8'h00;
            reg_file[25156] <= 8'h00;
            reg_file[25157] <= 8'h00;
            reg_file[25158] <= 8'h00;
            reg_file[25159] <= 8'h00;
            reg_file[25160] <= 8'h00;
            reg_file[25161] <= 8'h00;
            reg_file[25162] <= 8'h00;
            reg_file[25163] <= 8'h00;
            reg_file[25164] <= 8'h00;
            reg_file[25165] <= 8'h00;
            reg_file[25166] <= 8'h00;
            reg_file[25167] <= 8'h00;
            reg_file[25168] <= 8'h00;
            reg_file[25169] <= 8'h00;
            reg_file[25170] <= 8'h00;
            reg_file[25171] <= 8'h00;
            reg_file[25172] <= 8'h00;
            reg_file[25173] <= 8'h00;
            reg_file[25174] <= 8'h00;
            reg_file[25175] <= 8'h00;
            reg_file[25176] <= 8'h00;
            reg_file[25177] <= 8'h00;
            reg_file[25178] <= 8'h00;
            reg_file[25179] <= 8'h00;
            reg_file[25180] <= 8'h00;
            reg_file[25181] <= 8'h00;
            reg_file[25182] <= 8'h00;
            reg_file[25183] <= 8'h00;
            reg_file[25184] <= 8'h00;
            reg_file[25185] <= 8'h00;
            reg_file[25186] <= 8'h00;
            reg_file[25187] <= 8'h00;
            reg_file[25188] <= 8'h00;
            reg_file[25189] <= 8'h00;
            reg_file[25190] <= 8'h00;
            reg_file[25191] <= 8'h00;
            reg_file[25192] <= 8'h00;
            reg_file[25193] <= 8'h00;
            reg_file[25194] <= 8'h00;
            reg_file[25195] <= 8'h00;
            reg_file[25196] <= 8'h00;
            reg_file[25197] <= 8'h00;
            reg_file[25198] <= 8'h00;
            reg_file[25199] <= 8'h00;
            reg_file[25200] <= 8'h00;
            reg_file[25201] <= 8'h00;
            reg_file[25202] <= 8'h00;
            reg_file[25203] <= 8'h00;
            reg_file[25204] <= 8'h00;
            reg_file[25205] <= 8'h00;
            reg_file[25206] <= 8'h00;
            reg_file[25207] <= 8'h00;
            reg_file[25208] <= 8'h00;
            reg_file[25209] <= 8'h00;
            reg_file[25210] <= 8'h00;
            reg_file[25211] <= 8'h00;
            reg_file[25212] <= 8'h00;
            reg_file[25213] <= 8'h00;
            reg_file[25214] <= 8'h00;
            reg_file[25215] <= 8'h00;
            reg_file[25216] <= 8'h00;
            reg_file[25217] <= 8'h00;
            reg_file[25218] <= 8'h00;
            reg_file[25219] <= 8'h00;
            reg_file[25220] <= 8'h00;
            reg_file[25221] <= 8'h00;
            reg_file[25222] <= 8'h00;
            reg_file[25223] <= 8'h00;
            reg_file[25224] <= 8'h00;
            reg_file[25225] <= 8'h00;
            reg_file[25226] <= 8'h00;
            reg_file[25227] <= 8'h00;
            reg_file[25228] <= 8'h00;
            reg_file[25229] <= 8'h00;
            reg_file[25230] <= 8'h00;
            reg_file[25231] <= 8'h00;
            reg_file[25232] <= 8'h00;
            reg_file[25233] <= 8'h00;
            reg_file[25234] <= 8'h00;
            reg_file[25235] <= 8'h00;
            reg_file[25236] <= 8'h00;
            reg_file[25237] <= 8'h00;
            reg_file[25238] <= 8'h00;
            reg_file[25239] <= 8'h00;
            reg_file[25240] <= 8'h00;
            reg_file[25241] <= 8'h00;
            reg_file[25242] <= 8'h00;
            reg_file[25243] <= 8'h00;
            reg_file[25244] <= 8'h00;
            reg_file[25245] <= 8'h00;
            reg_file[25246] <= 8'h00;
            reg_file[25247] <= 8'h00;
            reg_file[25248] <= 8'h00;
            reg_file[25249] <= 8'h00;
            reg_file[25250] <= 8'h00;
            reg_file[25251] <= 8'h00;
            reg_file[25252] <= 8'h00;
            reg_file[25253] <= 8'h00;
            reg_file[25254] <= 8'h00;
            reg_file[25255] <= 8'h00;
            reg_file[25256] <= 8'h00;
            reg_file[25257] <= 8'h00;
            reg_file[25258] <= 8'h00;
            reg_file[25259] <= 8'h00;
            reg_file[25260] <= 8'h00;
            reg_file[25261] <= 8'h00;
            reg_file[25262] <= 8'h00;
            reg_file[25263] <= 8'h00;
            reg_file[25264] <= 8'h00;
            reg_file[25265] <= 8'h00;
            reg_file[25266] <= 8'h00;
            reg_file[25267] <= 8'h00;
            reg_file[25268] <= 8'h00;
            reg_file[25269] <= 8'h00;
            reg_file[25270] <= 8'h00;
            reg_file[25271] <= 8'h00;
            reg_file[25272] <= 8'h00;
            reg_file[25273] <= 8'h00;
            reg_file[25274] <= 8'h00;
            reg_file[25275] <= 8'h00;
            reg_file[25276] <= 8'h00;
            reg_file[25277] <= 8'h00;
            reg_file[25278] <= 8'h00;
            reg_file[25279] <= 8'h00;
            reg_file[25280] <= 8'h00;
            reg_file[25281] <= 8'h00;
            reg_file[25282] <= 8'h00;
            reg_file[25283] <= 8'h00;
            reg_file[25284] <= 8'h00;
            reg_file[25285] <= 8'h00;
            reg_file[25286] <= 8'h00;
            reg_file[25287] <= 8'h00;
            reg_file[25288] <= 8'h00;
            reg_file[25289] <= 8'h00;
            reg_file[25290] <= 8'h00;
            reg_file[25291] <= 8'h00;
            reg_file[25292] <= 8'h00;
            reg_file[25293] <= 8'h00;
            reg_file[25294] <= 8'h00;
            reg_file[25295] <= 8'h00;
            reg_file[25296] <= 8'h00;
            reg_file[25297] <= 8'h00;
            reg_file[25298] <= 8'h00;
            reg_file[25299] <= 8'h00;
            reg_file[25300] <= 8'h00;
            reg_file[25301] <= 8'h00;
            reg_file[25302] <= 8'h00;
            reg_file[25303] <= 8'h00;
            reg_file[25304] <= 8'h00;
            reg_file[25305] <= 8'h00;
            reg_file[25306] <= 8'h00;
            reg_file[25307] <= 8'h00;
            reg_file[25308] <= 8'h00;
            reg_file[25309] <= 8'h00;
            reg_file[25310] <= 8'h00;
            reg_file[25311] <= 8'h00;
            reg_file[25312] <= 8'h00;
            reg_file[25313] <= 8'h00;
            reg_file[25314] <= 8'h00;
            reg_file[25315] <= 8'h00;
            reg_file[25316] <= 8'h00;
            reg_file[25317] <= 8'h00;
            reg_file[25318] <= 8'h00;
            reg_file[25319] <= 8'h00;
            reg_file[25320] <= 8'h00;
            reg_file[25321] <= 8'h00;
            reg_file[25322] <= 8'h00;
            reg_file[25323] <= 8'h00;
            reg_file[25324] <= 8'h00;
            reg_file[25325] <= 8'h00;
            reg_file[25326] <= 8'h00;
            reg_file[25327] <= 8'h00;
            reg_file[25328] <= 8'h00;
            reg_file[25329] <= 8'h00;
            reg_file[25330] <= 8'h00;
            reg_file[25331] <= 8'h00;
            reg_file[25332] <= 8'h00;
            reg_file[25333] <= 8'h00;
            reg_file[25334] <= 8'h00;
            reg_file[25335] <= 8'h00;
            reg_file[25336] <= 8'h00;
            reg_file[25337] <= 8'h00;
            reg_file[25338] <= 8'h00;
            reg_file[25339] <= 8'h00;
            reg_file[25340] <= 8'h00;
            reg_file[25341] <= 8'h00;
            reg_file[25342] <= 8'h00;
            reg_file[25343] <= 8'h00;
            reg_file[25344] <= 8'h00;
            reg_file[25345] <= 8'h00;
            reg_file[25346] <= 8'h00;
            reg_file[25347] <= 8'h00;
            reg_file[25348] <= 8'h00;
            reg_file[25349] <= 8'h00;
            reg_file[25350] <= 8'h00;
            reg_file[25351] <= 8'h00;
            reg_file[25352] <= 8'h00;
            reg_file[25353] <= 8'h00;
            reg_file[25354] <= 8'h00;
            reg_file[25355] <= 8'h00;
            reg_file[25356] <= 8'h00;
            reg_file[25357] <= 8'h00;
            reg_file[25358] <= 8'h00;
            reg_file[25359] <= 8'h00;
            reg_file[25360] <= 8'h00;
            reg_file[25361] <= 8'h00;
            reg_file[25362] <= 8'h00;
            reg_file[25363] <= 8'h00;
            reg_file[25364] <= 8'h00;
            reg_file[25365] <= 8'h00;
            reg_file[25366] <= 8'h00;
            reg_file[25367] <= 8'h00;
            reg_file[25368] <= 8'h00;
            reg_file[25369] <= 8'h00;
            reg_file[25370] <= 8'h00;
            reg_file[25371] <= 8'h00;
            reg_file[25372] <= 8'h00;
            reg_file[25373] <= 8'h00;
            reg_file[25374] <= 8'h00;
            reg_file[25375] <= 8'h00;
            reg_file[25376] <= 8'h00;
            reg_file[25377] <= 8'h00;
            reg_file[25378] <= 8'h00;
            reg_file[25379] <= 8'h00;
            reg_file[25380] <= 8'h00;
            reg_file[25381] <= 8'h00;
            reg_file[25382] <= 8'h00;
            reg_file[25383] <= 8'h00;
            reg_file[25384] <= 8'h00;
            reg_file[25385] <= 8'h00;
            reg_file[25386] <= 8'h00;
            reg_file[25387] <= 8'h00;
            reg_file[25388] <= 8'h00;
            reg_file[25389] <= 8'h00;
            reg_file[25390] <= 8'h00;
            reg_file[25391] <= 8'h00;
            reg_file[25392] <= 8'h00;
            reg_file[25393] <= 8'h00;
            reg_file[25394] <= 8'h00;
            reg_file[25395] <= 8'h00;
            reg_file[25396] <= 8'h00;
            reg_file[25397] <= 8'h00;
            reg_file[25398] <= 8'h00;
            reg_file[25399] <= 8'h00;
            reg_file[25400] <= 8'h00;
            reg_file[25401] <= 8'h00;
            reg_file[25402] <= 8'h00;
            reg_file[25403] <= 8'h00;
            reg_file[25404] <= 8'h00;
            reg_file[25405] <= 8'h00;
            reg_file[25406] <= 8'h00;
            reg_file[25407] <= 8'h00;
            reg_file[25408] <= 8'h00;
            reg_file[25409] <= 8'h00;
            reg_file[25410] <= 8'h00;
            reg_file[25411] <= 8'h00;
            reg_file[25412] <= 8'h00;
            reg_file[25413] <= 8'h00;
            reg_file[25414] <= 8'h00;
            reg_file[25415] <= 8'h00;
            reg_file[25416] <= 8'h00;
            reg_file[25417] <= 8'h00;
            reg_file[25418] <= 8'h00;
            reg_file[25419] <= 8'h00;
            reg_file[25420] <= 8'h00;
            reg_file[25421] <= 8'h00;
            reg_file[25422] <= 8'h00;
            reg_file[25423] <= 8'h00;
            reg_file[25424] <= 8'h00;
            reg_file[25425] <= 8'h00;
            reg_file[25426] <= 8'h00;
            reg_file[25427] <= 8'h00;
            reg_file[25428] <= 8'h00;
            reg_file[25429] <= 8'h00;
            reg_file[25430] <= 8'h00;
            reg_file[25431] <= 8'h00;
            reg_file[25432] <= 8'h00;
            reg_file[25433] <= 8'h00;
            reg_file[25434] <= 8'h00;
            reg_file[25435] <= 8'h00;
            reg_file[25436] <= 8'h00;
            reg_file[25437] <= 8'h00;
            reg_file[25438] <= 8'h00;
            reg_file[25439] <= 8'h00;
            reg_file[25440] <= 8'h00;
            reg_file[25441] <= 8'h00;
            reg_file[25442] <= 8'h00;
            reg_file[25443] <= 8'h00;
            reg_file[25444] <= 8'h00;
            reg_file[25445] <= 8'h00;
            reg_file[25446] <= 8'h00;
            reg_file[25447] <= 8'h00;
            reg_file[25448] <= 8'h00;
            reg_file[25449] <= 8'h00;
            reg_file[25450] <= 8'h00;
            reg_file[25451] <= 8'h00;
            reg_file[25452] <= 8'h00;
            reg_file[25453] <= 8'h00;
            reg_file[25454] <= 8'h00;
            reg_file[25455] <= 8'h00;
            reg_file[25456] <= 8'h00;
            reg_file[25457] <= 8'h00;
            reg_file[25458] <= 8'h00;
            reg_file[25459] <= 8'h00;
            reg_file[25460] <= 8'h00;
            reg_file[25461] <= 8'h00;
            reg_file[25462] <= 8'h00;
            reg_file[25463] <= 8'h00;
            reg_file[25464] <= 8'h00;
            reg_file[25465] <= 8'h00;
            reg_file[25466] <= 8'h00;
            reg_file[25467] <= 8'h00;
            reg_file[25468] <= 8'h00;
            reg_file[25469] <= 8'h00;
            reg_file[25470] <= 8'h00;
            reg_file[25471] <= 8'h00;
            reg_file[25472] <= 8'h00;
            reg_file[25473] <= 8'h00;
            reg_file[25474] <= 8'h00;
            reg_file[25475] <= 8'h00;
            reg_file[25476] <= 8'h00;
            reg_file[25477] <= 8'h00;
            reg_file[25478] <= 8'h00;
            reg_file[25479] <= 8'h00;
            reg_file[25480] <= 8'h00;
            reg_file[25481] <= 8'h00;
            reg_file[25482] <= 8'h00;
            reg_file[25483] <= 8'h00;
            reg_file[25484] <= 8'h00;
            reg_file[25485] <= 8'h00;
            reg_file[25486] <= 8'h00;
            reg_file[25487] <= 8'h00;
            reg_file[25488] <= 8'h00;
            reg_file[25489] <= 8'h00;
            reg_file[25490] <= 8'h00;
            reg_file[25491] <= 8'h00;
            reg_file[25492] <= 8'h00;
            reg_file[25493] <= 8'h00;
            reg_file[25494] <= 8'h00;
            reg_file[25495] <= 8'h00;
            reg_file[25496] <= 8'h00;
            reg_file[25497] <= 8'h00;
            reg_file[25498] <= 8'h00;
            reg_file[25499] <= 8'h00;
            reg_file[25500] <= 8'h00;
            reg_file[25501] <= 8'h00;
            reg_file[25502] <= 8'h00;
            reg_file[25503] <= 8'h00;
            reg_file[25504] <= 8'h00;
            reg_file[25505] <= 8'h00;
            reg_file[25506] <= 8'h00;
            reg_file[25507] <= 8'h00;
            reg_file[25508] <= 8'h00;
            reg_file[25509] <= 8'h00;
            reg_file[25510] <= 8'h00;
            reg_file[25511] <= 8'h00;
            reg_file[25512] <= 8'h00;
            reg_file[25513] <= 8'h00;
            reg_file[25514] <= 8'h00;
            reg_file[25515] <= 8'h00;
            reg_file[25516] <= 8'h00;
            reg_file[25517] <= 8'h00;
            reg_file[25518] <= 8'h00;
            reg_file[25519] <= 8'h00;
            reg_file[25520] <= 8'h00;
            reg_file[25521] <= 8'h00;
            reg_file[25522] <= 8'h00;
            reg_file[25523] <= 8'h00;
            reg_file[25524] <= 8'h00;
            reg_file[25525] <= 8'h00;
            reg_file[25526] <= 8'h00;
            reg_file[25527] <= 8'h00;
            reg_file[25528] <= 8'h00;
            reg_file[25529] <= 8'h00;
            reg_file[25530] <= 8'h00;
            reg_file[25531] <= 8'h00;
            reg_file[25532] <= 8'h00;
            reg_file[25533] <= 8'h00;
            reg_file[25534] <= 8'h00;
            reg_file[25535] <= 8'h00;
            reg_file[25536] <= 8'h00;
            reg_file[25537] <= 8'h00;
            reg_file[25538] <= 8'h00;
            reg_file[25539] <= 8'h00;
            reg_file[25540] <= 8'h00;
            reg_file[25541] <= 8'h00;
            reg_file[25542] <= 8'h00;
            reg_file[25543] <= 8'h00;
            reg_file[25544] <= 8'h00;
            reg_file[25545] <= 8'h00;
            reg_file[25546] <= 8'h00;
            reg_file[25547] <= 8'h00;
            reg_file[25548] <= 8'h00;
            reg_file[25549] <= 8'h00;
            reg_file[25550] <= 8'h00;
            reg_file[25551] <= 8'h00;
            reg_file[25552] <= 8'h00;
            reg_file[25553] <= 8'h00;
            reg_file[25554] <= 8'h00;
            reg_file[25555] <= 8'h00;
            reg_file[25556] <= 8'h00;
            reg_file[25557] <= 8'h00;
            reg_file[25558] <= 8'h00;
            reg_file[25559] <= 8'h00;
            reg_file[25560] <= 8'h00;
            reg_file[25561] <= 8'h00;
            reg_file[25562] <= 8'h00;
            reg_file[25563] <= 8'h00;
            reg_file[25564] <= 8'h00;
            reg_file[25565] <= 8'h00;
            reg_file[25566] <= 8'h00;
            reg_file[25567] <= 8'h00;
            reg_file[25568] <= 8'h00;
            reg_file[25569] <= 8'h00;
            reg_file[25570] <= 8'h00;
            reg_file[25571] <= 8'h00;
            reg_file[25572] <= 8'h00;
            reg_file[25573] <= 8'h00;
            reg_file[25574] <= 8'h00;
            reg_file[25575] <= 8'h00;
            reg_file[25576] <= 8'h00;
            reg_file[25577] <= 8'h00;
            reg_file[25578] <= 8'h00;
            reg_file[25579] <= 8'h00;
            reg_file[25580] <= 8'h00;
            reg_file[25581] <= 8'h00;
            reg_file[25582] <= 8'h00;
            reg_file[25583] <= 8'h00;
            reg_file[25584] <= 8'h00;
            reg_file[25585] <= 8'h00;
            reg_file[25586] <= 8'h00;
            reg_file[25587] <= 8'h00;
            reg_file[25588] <= 8'h00;
            reg_file[25589] <= 8'h00;
            reg_file[25590] <= 8'h00;
            reg_file[25591] <= 8'h00;
            reg_file[25592] <= 8'h00;
            reg_file[25593] <= 8'h00;
            reg_file[25594] <= 8'h00;
            reg_file[25595] <= 8'h00;
            reg_file[25596] <= 8'h00;
            reg_file[25597] <= 8'h00;
            reg_file[25598] <= 8'h00;
            reg_file[25599] <= 8'h00;
            reg_file[25600] <= 8'h00;
            reg_file[25601] <= 8'h00;
            reg_file[25602] <= 8'h00;
            reg_file[25603] <= 8'h00;
            reg_file[25604] <= 8'h00;
            reg_file[25605] <= 8'h00;
            reg_file[25606] <= 8'h00;
            reg_file[25607] <= 8'h00;
            reg_file[25608] <= 8'h00;
            reg_file[25609] <= 8'h00;
            reg_file[25610] <= 8'h00;
            reg_file[25611] <= 8'h00;
            reg_file[25612] <= 8'h00;
            reg_file[25613] <= 8'h00;
            reg_file[25614] <= 8'h00;
            reg_file[25615] <= 8'h00;
            reg_file[25616] <= 8'h00;
            reg_file[25617] <= 8'h00;
            reg_file[25618] <= 8'h00;
            reg_file[25619] <= 8'h00;
            reg_file[25620] <= 8'h00;
            reg_file[25621] <= 8'h00;
            reg_file[25622] <= 8'h00;
            reg_file[25623] <= 8'h00;
            reg_file[25624] <= 8'h00;
            reg_file[25625] <= 8'h00;
            reg_file[25626] <= 8'h00;
            reg_file[25627] <= 8'h00;
            reg_file[25628] <= 8'h00;
            reg_file[25629] <= 8'h00;
            reg_file[25630] <= 8'h00;
            reg_file[25631] <= 8'h00;
            reg_file[25632] <= 8'h00;
            reg_file[25633] <= 8'h00;
            reg_file[25634] <= 8'h00;
            reg_file[25635] <= 8'h00;
            reg_file[25636] <= 8'h00;
            reg_file[25637] <= 8'h00;
            reg_file[25638] <= 8'h00;
            reg_file[25639] <= 8'h00;
            reg_file[25640] <= 8'h00;
            reg_file[25641] <= 8'h00;
            reg_file[25642] <= 8'h00;
            reg_file[25643] <= 8'h00;
            reg_file[25644] <= 8'h00;
            reg_file[25645] <= 8'h00;
            reg_file[25646] <= 8'h00;
            reg_file[25647] <= 8'h00;
            reg_file[25648] <= 8'h00;
            reg_file[25649] <= 8'h00;
            reg_file[25650] <= 8'h00;
            reg_file[25651] <= 8'h00;
            reg_file[25652] <= 8'h00;
            reg_file[25653] <= 8'h00;
            reg_file[25654] <= 8'h00;
            reg_file[25655] <= 8'h00;
            reg_file[25656] <= 8'h00;
            reg_file[25657] <= 8'h00;
            reg_file[25658] <= 8'h00;
            reg_file[25659] <= 8'h00;
            reg_file[25660] <= 8'h00;
            reg_file[25661] <= 8'h00;
            reg_file[25662] <= 8'h00;
            reg_file[25663] <= 8'h00;
            reg_file[25664] <= 8'h00;
            reg_file[25665] <= 8'h00;
            reg_file[25666] <= 8'h00;
            reg_file[25667] <= 8'h00;
            reg_file[25668] <= 8'h00;
            reg_file[25669] <= 8'h00;
            reg_file[25670] <= 8'h00;
            reg_file[25671] <= 8'h00;
            reg_file[25672] <= 8'h00;
            reg_file[25673] <= 8'h00;
            reg_file[25674] <= 8'h00;
            reg_file[25675] <= 8'h00;
            reg_file[25676] <= 8'h00;
            reg_file[25677] <= 8'h00;
            reg_file[25678] <= 8'h00;
            reg_file[25679] <= 8'h00;
            reg_file[25680] <= 8'h00;
            reg_file[25681] <= 8'h00;
            reg_file[25682] <= 8'h00;
            reg_file[25683] <= 8'h00;
            reg_file[25684] <= 8'h00;
            reg_file[25685] <= 8'h00;
            reg_file[25686] <= 8'h00;
            reg_file[25687] <= 8'h00;
            reg_file[25688] <= 8'h00;
            reg_file[25689] <= 8'h00;
            reg_file[25690] <= 8'h00;
            reg_file[25691] <= 8'h00;
            reg_file[25692] <= 8'h00;
            reg_file[25693] <= 8'h00;
            reg_file[25694] <= 8'h00;
            reg_file[25695] <= 8'h00;
            reg_file[25696] <= 8'h00;
            reg_file[25697] <= 8'h00;
            reg_file[25698] <= 8'h00;
            reg_file[25699] <= 8'h00;
            reg_file[25700] <= 8'h00;
            reg_file[25701] <= 8'h00;
            reg_file[25702] <= 8'h00;
            reg_file[25703] <= 8'h00;
            reg_file[25704] <= 8'h00;
            reg_file[25705] <= 8'h00;
            reg_file[25706] <= 8'h00;
            reg_file[25707] <= 8'h00;
            reg_file[25708] <= 8'h00;
            reg_file[25709] <= 8'h00;
            reg_file[25710] <= 8'h00;
            reg_file[25711] <= 8'h00;
            reg_file[25712] <= 8'h00;
            reg_file[25713] <= 8'h00;
            reg_file[25714] <= 8'h00;
            reg_file[25715] <= 8'h00;
            reg_file[25716] <= 8'h00;
            reg_file[25717] <= 8'h00;
            reg_file[25718] <= 8'h00;
            reg_file[25719] <= 8'h00;
            reg_file[25720] <= 8'h00;
            reg_file[25721] <= 8'h00;
            reg_file[25722] <= 8'h00;
            reg_file[25723] <= 8'h00;
            reg_file[25724] <= 8'h00;
            reg_file[25725] <= 8'h00;
            reg_file[25726] <= 8'h00;
            reg_file[25727] <= 8'h00;
            reg_file[25728] <= 8'h00;
            reg_file[25729] <= 8'h00;
            reg_file[25730] <= 8'h00;
            reg_file[25731] <= 8'h00;
            reg_file[25732] <= 8'h00;
            reg_file[25733] <= 8'h00;
            reg_file[25734] <= 8'h00;
            reg_file[25735] <= 8'h00;
            reg_file[25736] <= 8'h00;
            reg_file[25737] <= 8'h00;
            reg_file[25738] <= 8'h00;
            reg_file[25739] <= 8'h00;
            reg_file[25740] <= 8'h00;
            reg_file[25741] <= 8'h00;
            reg_file[25742] <= 8'h00;
            reg_file[25743] <= 8'h00;
            reg_file[25744] <= 8'h00;
            reg_file[25745] <= 8'h00;
            reg_file[25746] <= 8'h00;
            reg_file[25747] <= 8'h00;
            reg_file[25748] <= 8'h00;
            reg_file[25749] <= 8'h00;
            reg_file[25750] <= 8'h00;
            reg_file[25751] <= 8'h00;
            reg_file[25752] <= 8'h00;
            reg_file[25753] <= 8'h00;
            reg_file[25754] <= 8'h00;
            reg_file[25755] <= 8'h00;
            reg_file[25756] <= 8'h00;
            reg_file[25757] <= 8'h00;
            reg_file[25758] <= 8'h00;
            reg_file[25759] <= 8'h00;
            reg_file[25760] <= 8'h00;
            reg_file[25761] <= 8'h00;
            reg_file[25762] <= 8'h00;
            reg_file[25763] <= 8'h00;
            reg_file[25764] <= 8'h00;
            reg_file[25765] <= 8'h00;
            reg_file[25766] <= 8'h00;
            reg_file[25767] <= 8'h00;
            reg_file[25768] <= 8'h00;
            reg_file[25769] <= 8'h00;
            reg_file[25770] <= 8'h00;
            reg_file[25771] <= 8'h00;
            reg_file[25772] <= 8'h00;
            reg_file[25773] <= 8'h00;
            reg_file[25774] <= 8'h00;
            reg_file[25775] <= 8'h00;
            reg_file[25776] <= 8'h00;
            reg_file[25777] <= 8'h00;
            reg_file[25778] <= 8'h00;
            reg_file[25779] <= 8'h00;
            reg_file[25780] <= 8'h00;
            reg_file[25781] <= 8'h00;
            reg_file[25782] <= 8'h00;
            reg_file[25783] <= 8'h00;
            reg_file[25784] <= 8'h00;
            reg_file[25785] <= 8'h00;
            reg_file[25786] <= 8'h00;
            reg_file[25787] <= 8'h00;
            reg_file[25788] <= 8'h00;
            reg_file[25789] <= 8'h00;
            reg_file[25790] <= 8'h00;
            reg_file[25791] <= 8'h00;
            reg_file[25792] <= 8'h00;
            reg_file[25793] <= 8'h00;
            reg_file[25794] <= 8'h00;
            reg_file[25795] <= 8'h00;
            reg_file[25796] <= 8'h00;
            reg_file[25797] <= 8'h00;
            reg_file[25798] <= 8'h00;
            reg_file[25799] <= 8'h00;
            reg_file[25800] <= 8'h00;
            reg_file[25801] <= 8'h00;
            reg_file[25802] <= 8'h00;
            reg_file[25803] <= 8'h00;
            reg_file[25804] <= 8'h00;
            reg_file[25805] <= 8'h00;
            reg_file[25806] <= 8'h00;
            reg_file[25807] <= 8'h00;
            reg_file[25808] <= 8'h00;
            reg_file[25809] <= 8'h00;
            reg_file[25810] <= 8'h00;
            reg_file[25811] <= 8'h00;
            reg_file[25812] <= 8'h00;
            reg_file[25813] <= 8'h00;
            reg_file[25814] <= 8'h00;
            reg_file[25815] <= 8'h00;
            reg_file[25816] <= 8'h00;
            reg_file[25817] <= 8'h00;
            reg_file[25818] <= 8'h00;
            reg_file[25819] <= 8'h00;
            reg_file[25820] <= 8'h00;
            reg_file[25821] <= 8'h00;
            reg_file[25822] <= 8'h00;
            reg_file[25823] <= 8'h00;
            reg_file[25824] <= 8'h00;
            reg_file[25825] <= 8'h00;
            reg_file[25826] <= 8'h00;
            reg_file[25827] <= 8'h00;
            reg_file[25828] <= 8'h00;
            reg_file[25829] <= 8'h00;
            reg_file[25830] <= 8'h00;
            reg_file[25831] <= 8'h00;
            reg_file[25832] <= 8'h00;
            reg_file[25833] <= 8'h00;
            reg_file[25834] <= 8'h00;
            reg_file[25835] <= 8'h00;
            reg_file[25836] <= 8'h00;
            reg_file[25837] <= 8'h00;
            reg_file[25838] <= 8'h00;
            reg_file[25839] <= 8'h00;
            reg_file[25840] <= 8'h00;
            reg_file[25841] <= 8'h00;
            reg_file[25842] <= 8'h00;
            reg_file[25843] <= 8'h00;
            reg_file[25844] <= 8'h00;
            reg_file[25845] <= 8'h00;
            reg_file[25846] <= 8'h00;
            reg_file[25847] <= 8'h00;
            reg_file[25848] <= 8'h00;
            reg_file[25849] <= 8'h00;
            reg_file[25850] <= 8'h00;
            reg_file[25851] <= 8'h00;
            reg_file[25852] <= 8'h00;
            reg_file[25853] <= 8'h00;
            reg_file[25854] <= 8'h00;
            reg_file[25855] <= 8'h00;
            reg_file[25856] <= 8'h00;
            reg_file[25857] <= 8'h00;
            reg_file[25858] <= 8'h00;
            reg_file[25859] <= 8'h00;
            reg_file[25860] <= 8'h00;
            reg_file[25861] <= 8'h00;
            reg_file[25862] <= 8'h00;
            reg_file[25863] <= 8'h00;
            reg_file[25864] <= 8'h00;
            reg_file[25865] <= 8'h00;
            reg_file[25866] <= 8'h00;
            reg_file[25867] <= 8'h00;
            reg_file[25868] <= 8'h00;
            reg_file[25869] <= 8'h00;
            reg_file[25870] <= 8'h00;
            reg_file[25871] <= 8'h00;
            reg_file[25872] <= 8'h00;
            reg_file[25873] <= 8'h00;
            reg_file[25874] <= 8'h00;
            reg_file[25875] <= 8'h00;
            reg_file[25876] <= 8'h00;
            reg_file[25877] <= 8'h00;
            reg_file[25878] <= 8'h00;
            reg_file[25879] <= 8'h00;
            reg_file[25880] <= 8'h00;
            reg_file[25881] <= 8'h00;
            reg_file[25882] <= 8'h00;
            reg_file[25883] <= 8'h00;
            reg_file[25884] <= 8'h00;
            reg_file[25885] <= 8'h00;
            reg_file[25886] <= 8'h00;
            reg_file[25887] <= 8'h00;
            reg_file[25888] <= 8'h00;
            reg_file[25889] <= 8'h00;
            reg_file[25890] <= 8'h00;
            reg_file[25891] <= 8'h00;
            reg_file[25892] <= 8'h00;
            reg_file[25893] <= 8'h00;
            reg_file[25894] <= 8'h00;
            reg_file[25895] <= 8'h00;
            reg_file[25896] <= 8'h00;
            reg_file[25897] <= 8'h00;
            reg_file[25898] <= 8'h00;
            reg_file[25899] <= 8'h00;
            reg_file[25900] <= 8'h00;
            reg_file[25901] <= 8'h00;
            reg_file[25902] <= 8'h00;
            reg_file[25903] <= 8'h00;
            reg_file[25904] <= 8'h00;
            reg_file[25905] <= 8'h00;
            reg_file[25906] <= 8'h00;
            reg_file[25907] <= 8'h00;
            reg_file[25908] <= 8'h00;
            reg_file[25909] <= 8'h00;
            reg_file[25910] <= 8'h00;
            reg_file[25911] <= 8'h00;
            reg_file[25912] <= 8'h00;
            reg_file[25913] <= 8'h00;
            reg_file[25914] <= 8'h00;
            reg_file[25915] <= 8'h00;
            reg_file[25916] <= 8'h00;
            reg_file[25917] <= 8'h00;
            reg_file[25918] <= 8'h00;
            reg_file[25919] <= 8'h00;
            reg_file[25920] <= 8'h00;
            reg_file[25921] <= 8'h00;
            reg_file[25922] <= 8'h00;
            reg_file[25923] <= 8'h00;
            reg_file[25924] <= 8'h00;
            reg_file[25925] <= 8'h00;
            reg_file[25926] <= 8'h00;
            reg_file[25927] <= 8'h00;
            reg_file[25928] <= 8'h00;
            reg_file[25929] <= 8'h00;
            reg_file[25930] <= 8'h00;
            reg_file[25931] <= 8'h00;
            reg_file[25932] <= 8'h00;
            reg_file[25933] <= 8'h00;
            reg_file[25934] <= 8'h00;
            reg_file[25935] <= 8'h00;
            reg_file[25936] <= 8'h00;
            reg_file[25937] <= 8'h00;
            reg_file[25938] <= 8'h00;
            reg_file[25939] <= 8'h00;
            reg_file[25940] <= 8'h00;
            reg_file[25941] <= 8'h00;
            reg_file[25942] <= 8'h00;
            reg_file[25943] <= 8'h00;
            reg_file[25944] <= 8'h00;
            reg_file[25945] <= 8'h00;
            reg_file[25946] <= 8'h00;
            reg_file[25947] <= 8'h00;
            reg_file[25948] <= 8'h00;
            reg_file[25949] <= 8'h00;
            reg_file[25950] <= 8'h00;
            reg_file[25951] <= 8'h00;
            reg_file[25952] <= 8'h00;
            reg_file[25953] <= 8'h00;
            reg_file[25954] <= 8'h00;
            reg_file[25955] <= 8'h00;
            reg_file[25956] <= 8'h00;
            reg_file[25957] <= 8'h00;
            reg_file[25958] <= 8'h00;
            reg_file[25959] <= 8'h00;
            reg_file[25960] <= 8'h00;
            reg_file[25961] <= 8'h00;
            reg_file[25962] <= 8'h00;
            reg_file[25963] <= 8'h00;
            reg_file[25964] <= 8'h00;
            reg_file[25965] <= 8'h00;
            reg_file[25966] <= 8'h00;
            reg_file[25967] <= 8'h00;
            reg_file[25968] <= 8'h00;
            reg_file[25969] <= 8'h00;
            reg_file[25970] <= 8'h00;
            reg_file[25971] <= 8'h00;
            reg_file[25972] <= 8'h00;
            reg_file[25973] <= 8'h00;
            reg_file[25974] <= 8'h00;
            reg_file[25975] <= 8'h00;
            reg_file[25976] <= 8'h00;
            reg_file[25977] <= 8'h00;
            reg_file[25978] <= 8'h00;
            reg_file[25979] <= 8'h00;
            reg_file[25980] <= 8'h00;
            reg_file[25981] <= 8'h00;
            reg_file[25982] <= 8'h00;
            reg_file[25983] <= 8'h00;
            reg_file[25984] <= 8'h00;
            reg_file[25985] <= 8'h00;
            reg_file[25986] <= 8'h00;
            reg_file[25987] <= 8'h00;
            reg_file[25988] <= 8'h00;
            reg_file[25989] <= 8'h00;
            reg_file[25990] <= 8'h00;
            reg_file[25991] <= 8'h00;
            reg_file[25992] <= 8'h00;
            reg_file[25993] <= 8'h00;
            reg_file[25994] <= 8'h00;
            reg_file[25995] <= 8'h00;
            reg_file[25996] <= 8'h00;
            reg_file[25997] <= 8'h00;
            reg_file[25998] <= 8'h00;
            reg_file[25999] <= 8'h00;
            reg_file[26000] <= 8'h00;
            reg_file[26001] <= 8'h00;
            reg_file[26002] <= 8'h00;
            reg_file[26003] <= 8'h00;
            reg_file[26004] <= 8'h00;
            reg_file[26005] <= 8'h00;
            reg_file[26006] <= 8'h00;
            reg_file[26007] <= 8'h00;
            reg_file[26008] <= 8'h00;
            reg_file[26009] <= 8'h00;
            reg_file[26010] <= 8'h00;
            reg_file[26011] <= 8'h00;
            reg_file[26012] <= 8'h00;
            reg_file[26013] <= 8'h00;
            reg_file[26014] <= 8'h00;
            reg_file[26015] <= 8'h00;
            reg_file[26016] <= 8'h00;
            reg_file[26017] <= 8'h00;
            reg_file[26018] <= 8'h00;
            reg_file[26019] <= 8'h00;
            reg_file[26020] <= 8'h00;
            reg_file[26021] <= 8'h00;
            reg_file[26022] <= 8'h00;
            reg_file[26023] <= 8'h00;
            reg_file[26024] <= 8'h00;
            reg_file[26025] <= 8'h00;
            reg_file[26026] <= 8'h00;
            reg_file[26027] <= 8'h00;
            reg_file[26028] <= 8'h00;
            reg_file[26029] <= 8'h00;
            reg_file[26030] <= 8'h00;
            reg_file[26031] <= 8'h00;
            reg_file[26032] <= 8'h00;
            reg_file[26033] <= 8'h00;
            reg_file[26034] <= 8'h00;
            reg_file[26035] <= 8'h00;
            reg_file[26036] <= 8'h00;
            reg_file[26037] <= 8'h00;
            reg_file[26038] <= 8'h00;
            reg_file[26039] <= 8'h00;
            reg_file[26040] <= 8'h00;
            reg_file[26041] <= 8'h00;
            reg_file[26042] <= 8'h00;
            reg_file[26043] <= 8'h00;
            reg_file[26044] <= 8'h00;
            reg_file[26045] <= 8'h00;
            reg_file[26046] <= 8'h00;
            reg_file[26047] <= 8'h00;
            reg_file[26048] <= 8'h00;
            reg_file[26049] <= 8'h00;
            reg_file[26050] <= 8'h00;
            reg_file[26051] <= 8'h00;
            reg_file[26052] <= 8'h00;
            reg_file[26053] <= 8'h00;
            reg_file[26054] <= 8'h00;
            reg_file[26055] <= 8'h00;
            reg_file[26056] <= 8'h00;
            reg_file[26057] <= 8'h00;
            reg_file[26058] <= 8'h00;
            reg_file[26059] <= 8'h00;
            reg_file[26060] <= 8'h00;
            reg_file[26061] <= 8'h00;
            reg_file[26062] <= 8'h00;
            reg_file[26063] <= 8'h00;
            reg_file[26064] <= 8'h00;
            reg_file[26065] <= 8'h00;
            reg_file[26066] <= 8'h00;
            reg_file[26067] <= 8'h00;
            reg_file[26068] <= 8'h00;
            reg_file[26069] <= 8'h00;
            reg_file[26070] <= 8'h00;
            reg_file[26071] <= 8'h00;
            reg_file[26072] <= 8'h00;
            reg_file[26073] <= 8'h00;
            reg_file[26074] <= 8'h00;
            reg_file[26075] <= 8'h00;
            reg_file[26076] <= 8'h00;
            reg_file[26077] <= 8'h00;
            reg_file[26078] <= 8'h00;
            reg_file[26079] <= 8'h00;
            reg_file[26080] <= 8'h00;
            reg_file[26081] <= 8'h00;
            reg_file[26082] <= 8'h00;
            reg_file[26083] <= 8'h00;
            reg_file[26084] <= 8'h00;
            reg_file[26085] <= 8'h00;
            reg_file[26086] <= 8'h00;
            reg_file[26087] <= 8'h00;
            reg_file[26088] <= 8'h00;
            reg_file[26089] <= 8'h00;
            reg_file[26090] <= 8'h00;
            reg_file[26091] <= 8'h00;
            reg_file[26092] <= 8'h00;
            reg_file[26093] <= 8'h00;
            reg_file[26094] <= 8'h00;
            reg_file[26095] <= 8'h00;
            reg_file[26096] <= 8'h00;
            reg_file[26097] <= 8'h00;
            reg_file[26098] <= 8'h00;
            reg_file[26099] <= 8'h00;
            reg_file[26100] <= 8'h00;
            reg_file[26101] <= 8'h00;
            reg_file[26102] <= 8'h00;
            reg_file[26103] <= 8'h00;
            reg_file[26104] <= 8'h00;
            reg_file[26105] <= 8'h00;
            reg_file[26106] <= 8'h00;
            reg_file[26107] <= 8'h00;
            reg_file[26108] <= 8'h00;
            reg_file[26109] <= 8'h00;
            reg_file[26110] <= 8'h00;
            reg_file[26111] <= 8'h00;
            reg_file[26112] <= 8'h00;
            reg_file[26113] <= 8'h00;
            reg_file[26114] <= 8'h00;
            reg_file[26115] <= 8'h00;
            reg_file[26116] <= 8'h00;
            reg_file[26117] <= 8'h00;
            reg_file[26118] <= 8'h00;
            reg_file[26119] <= 8'h00;
            reg_file[26120] <= 8'h00;
            reg_file[26121] <= 8'h00;
            reg_file[26122] <= 8'h00;
            reg_file[26123] <= 8'h00;
            reg_file[26124] <= 8'h00;
            reg_file[26125] <= 8'h00;
            reg_file[26126] <= 8'h00;
            reg_file[26127] <= 8'h00;
            reg_file[26128] <= 8'h00;
            reg_file[26129] <= 8'h00;
            reg_file[26130] <= 8'h00;
            reg_file[26131] <= 8'h00;
            reg_file[26132] <= 8'h00;
            reg_file[26133] <= 8'h00;
            reg_file[26134] <= 8'h00;
            reg_file[26135] <= 8'h00;
            reg_file[26136] <= 8'h00;
            reg_file[26137] <= 8'h00;
            reg_file[26138] <= 8'h00;
            reg_file[26139] <= 8'h00;
            reg_file[26140] <= 8'h00;
            reg_file[26141] <= 8'h00;
            reg_file[26142] <= 8'h00;
            reg_file[26143] <= 8'h00;
            reg_file[26144] <= 8'h00;
            reg_file[26145] <= 8'h00;
            reg_file[26146] <= 8'h00;
            reg_file[26147] <= 8'h00;
            reg_file[26148] <= 8'h00;
            reg_file[26149] <= 8'h00;
            reg_file[26150] <= 8'h00;
            reg_file[26151] <= 8'h00;
            reg_file[26152] <= 8'h00;
            reg_file[26153] <= 8'h00;
            reg_file[26154] <= 8'h00;
            reg_file[26155] <= 8'h00;
            reg_file[26156] <= 8'h00;
            reg_file[26157] <= 8'h00;
            reg_file[26158] <= 8'h00;
            reg_file[26159] <= 8'h00;
            reg_file[26160] <= 8'h00;
            reg_file[26161] <= 8'h00;
            reg_file[26162] <= 8'h00;
            reg_file[26163] <= 8'h00;
            reg_file[26164] <= 8'h00;
            reg_file[26165] <= 8'h00;
            reg_file[26166] <= 8'h00;
            reg_file[26167] <= 8'h00;
            reg_file[26168] <= 8'h00;
            reg_file[26169] <= 8'h00;
            reg_file[26170] <= 8'h00;
            reg_file[26171] <= 8'h00;
            reg_file[26172] <= 8'h00;
            reg_file[26173] <= 8'h00;
            reg_file[26174] <= 8'h00;
            reg_file[26175] <= 8'h00;
            reg_file[26176] <= 8'h00;
            reg_file[26177] <= 8'h00;
            reg_file[26178] <= 8'h00;
            reg_file[26179] <= 8'h00;
            reg_file[26180] <= 8'h00;
            reg_file[26181] <= 8'h00;
            reg_file[26182] <= 8'h00;
            reg_file[26183] <= 8'h00;
            reg_file[26184] <= 8'h00;
            reg_file[26185] <= 8'h00;
            reg_file[26186] <= 8'h00;
            reg_file[26187] <= 8'h00;
            reg_file[26188] <= 8'h00;
            reg_file[26189] <= 8'h00;
            reg_file[26190] <= 8'h00;
            reg_file[26191] <= 8'h00;
            reg_file[26192] <= 8'h00;
            reg_file[26193] <= 8'h00;
            reg_file[26194] <= 8'h00;
            reg_file[26195] <= 8'h00;
            reg_file[26196] <= 8'h00;
            reg_file[26197] <= 8'h00;
            reg_file[26198] <= 8'h00;
            reg_file[26199] <= 8'h00;
            reg_file[26200] <= 8'h00;
            reg_file[26201] <= 8'h00;
            reg_file[26202] <= 8'h00;
            reg_file[26203] <= 8'h00;
            reg_file[26204] <= 8'h00;
            reg_file[26205] <= 8'h00;
            reg_file[26206] <= 8'h00;
            reg_file[26207] <= 8'h00;
            reg_file[26208] <= 8'h00;
            reg_file[26209] <= 8'h00;
            reg_file[26210] <= 8'h00;
            reg_file[26211] <= 8'h00;
            reg_file[26212] <= 8'h00;
            reg_file[26213] <= 8'h00;
            reg_file[26214] <= 8'h00;
            reg_file[26215] <= 8'h00;
            reg_file[26216] <= 8'h00;
            reg_file[26217] <= 8'h00;
            reg_file[26218] <= 8'h00;
            reg_file[26219] <= 8'h00;
            reg_file[26220] <= 8'h00;
            reg_file[26221] <= 8'h00;
            reg_file[26222] <= 8'h00;
            reg_file[26223] <= 8'h00;
            reg_file[26224] <= 8'h00;
            reg_file[26225] <= 8'h00;
            reg_file[26226] <= 8'h00;
            reg_file[26227] <= 8'h00;
            reg_file[26228] <= 8'h00;
            reg_file[26229] <= 8'h00;
            reg_file[26230] <= 8'h00;
            reg_file[26231] <= 8'h00;
            reg_file[26232] <= 8'h00;
            reg_file[26233] <= 8'h00;
            reg_file[26234] <= 8'h00;
            reg_file[26235] <= 8'h00;
            reg_file[26236] <= 8'h00;
            reg_file[26237] <= 8'h00;
            reg_file[26238] <= 8'h00;
            reg_file[26239] <= 8'h00;
            reg_file[26240] <= 8'h00;
            reg_file[26241] <= 8'h00;
            reg_file[26242] <= 8'h00;
            reg_file[26243] <= 8'h00;
            reg_file[26244] <= 8'h00;
            reg_file[26245] <= 8'h00;
            reg_file[26246] <= 8'h00;
            reg_file[26247] <= 8'h00;
            reg_file[26248] <= 8'h00;
            reg_file[26249] <= 8'h00;
            reg_file[26250] <= 8'h00;
            reg_file[26251] <= 8'h00;
            reg_file[26252] <= 8'h00;
            reg_file[26253] <= 8'h00;
            reg_file[26254] <= 8'h00;
            reg_file[26255] <= 8'h00;
            reg_file[26256] <= 8'h00;
            reg_file[26257] <= 8'h00;
            reg_file[26258] <= 8'h00;
            reg_file[26259] <= 8'h00;
            reg_file[26260] <= 8'h00;
            reg_file[26261] <= 8'h00;
            reg_file[26262] <= 8'h00;
            reg_file[26263] <= 8'h00;
            reg_file[26264] <= 8'h00;
            reg_file[26265] <= 8'h00;
            reg_file[26266] <= 8'h00;
            reg_file[26267] <= 8'h00;
            reg_file[26268] <= 8'h00;
            reg_file[26269] <= 8'h00;
            reg_file[26270] <= 8'h00;
            reg_file[26271] <= 8'h00;
            reg_file[26272] <= 8'h00;
            reg_file[26273] <= 8'h00;
            reg_file[26274] <= 8'h00;
            reg_file[26275] <= 8'h00;
            reg_file[26276] <= 8'h00;
            reg_file[26277] <= 8'h00;
            reg_file[26278] <= 8'h00;
            reg_file[26279] <= 8'h00;
            reg_file[26280] <= 8'h00;
            reg_file[26281] <= 8'h00;
            reg_file[26282] <= 8'h00;
            reg_file[26283] <= 8'h00;
            reg_file[26284] <= 8'h00;
            reg_file[26285] <= 8'h00;
            reg_file[26286] <= 8'h00;
            reg_file[26287] <= 8'h00;
            reg_file[26288] <= 8'h00;
            reg_file[26289] <= 8'h00;
            reg_file[26290] <= 8'h00;
            reg_file[26291] <= 8'h00;
            reg_file[26292] <= 8'h00;
            reg_file[26293] <= 8'h00;
            reg_file[26294] <= 8'h00;
            reg_file[26295] <= 8'h00;
            reg_file[26296] <= 8'h00;
            reg_file[26297] <= 8'h00;
            reg_file[26298] <= 8'h00;
            reg_file[26299] <= 8'h00;
            reg_file[26300] <= 8'h00;
            reg_file[26301] <= 8'h00;
            reg_file[26302] <= 8'h00;
            reg_file[26303] <= 8'h00;
            reg_file[26304] <= 8'h00;
            reg_file[26305] <= 8'h00;
            reg_file[26306] <= 8'h00;
            reg_file[26307] <= 8'h00;
            reg_file[26308] <= 8'h00;
            reg_file[26309] <= 8'h00;
            reg_file[26310] <= 8'h00;
            reg_file[26311] <= 8'h00;
            reg_file[26312] <= 8'h00;
            reg_file[26313] <= 8'h00;
            reg_file[26314] <= 8'h00;
            reg_file[26315] <= 8'h00;
            reg_file[26316] <= 8'h00;
            reg_file[26317] <= 8'h00;
            reg_file[26318] <= 8'h00;
            reg_file[26319] <= 8'h00;
            reg_file[26320] <= 8'h00;
            reg_file[26321] <= 8'h00;
            reg_file[26322] <= 8'h00;
            reg_file[26323] <= 8'h00;
            reg_file[26324] <= 8'h00;
            reg_file[26325] <= 8'h00;
            reg_file[26326] <= 8'h00;
            reg_file[26327] <= 8'h00;
            reg_file[26328] <= 8'h00;
            reg_file[26329] <= 8'h00;
            reg_file[26330] <= 8'h00;
            reg_file[26331] <= 8'h00;
            reg_file[26332] <= 8'h00;
            reg_file[26333] <= 8'h00;
            reg_file[26334] <= 8'h00;
            reg_file[26335] <= 8'h00;
            reg_file[26336] <= 8'h00;
            reg_file[26337] <= 8'h00;
            reg_file[26338] <= 8'h00;
            reg_file[26339] <= 8'h00;
            reg_file[26340] <= 8'h00;
            reg_file[26341] <= 8'h00;
            reg_file[26342] <= 8'h00;
            reg_file[26343] <= 8'h00;
            reg_file[26344] <= 8'h00;
            reg_file[26345] <= 8'h00;
            reg_file[26346] <= 8'h00;
            reg_file[26347] <= 8'h00;
            reg_file[26348] <= 8'h00;
            reg_file[26349] <= 8'h00;
            reg_file[26350] <= 8'h00;
            reg_file[26351] <= 8'h00;
            reg_file[26352] <= 8'h00;
            reg_file[26353] <= 8'h00;
            reg_file[26354] <= 8'h00;
            reg_file[26355] <= 8'h00;
            reg_file[26356] <= 8'h00;
            reg_file[26357] <= 8'h00;
            reg_file[26358] <= 8'h00;
            reg_file[26359] <= 8'h00;
            reg_file[26360] <= 8'h00;
            reg_file[26361] <= 8'h00;
            reg_file[26362] <= 8'h00;
            reg_file[26363] <= 8'h00;
            reg_file[26364] <= 8'h00;
            reg_file[26365] <= 8'h00;
            reg_file[26366] <= 8'h00;
            reg_file[26367] <= 8'h00;
            reg_file[26368] <= 8'h00;
            reg_file[26369] <= 8'h00;
            reg_file[26370] <= 8'h00;
            reg_file[26371] <= 8'h00;
            reg_file[26372] <= 8'h00;
            reg_file[26373] <= 8'h00;
            reg_file[26374] <= 8'h00;
            reg_file[26375] <= 8'h00;
            reg_file[26376] <= 8'h00;
            reg_file[26377] <= 8'h00;
            reg_file[26378] <= 8'h00;
            reg_file[26379] <= 8'h00;
            reg_file[26380] <= 8'h00;
            reg_file[26381] <= 8'h00;
            reg_file[26382] <= 8'h00;
            reg_file[26383] <= 8'h00;
            reg_file[26384] <= 8'h00;
            reg_file[26385] <= 8'h00;
            reg_file[26386] <= 8'h00;
            reg_file[26387] <= 8'h00;
            reg_file[26388] <= 8'h00;
            reg_file[26389] <= 8'h00;
            reg_file[26390] <= 8'h00;
            reg_file[26391] <= 8'h00;
            reg_file[26392] <= 8'h00;
            reg_file[26393] <= 8'h00;
            reg_file[26394] <= 8'h00;
            reg_file[26395] <= 8'h00;
            reg_file[26396] <= 8'h00;
            reg_file[26397] <= 8'h00;
            reg_file[26398] <= 8'h00;
            reg_file[26399] <= 8'h00;
            reg_file[26400] <= 8'h00;
            reg_file[26401] <= 8'h00;
            reg_file[26402] <= 8'h00;
            reg_file[26403] <= 8'h00;
            reg_file[26404] <= 8'h00;
            reg_file[26405] <= 8'h00;
            reg_file[26406] <= 8'h00;
            reg_file[26407] <= 8'h00;
            reg_file[26408] <= 8'h00;
            reg_file[26409] <= 8'h00;
            reg_file[26410] <= 8'h00;
            reg_file[26411] <= 8'h00;
            reg_file[26412] <= 8'h00;
            reg_file[26413] <= 8'h00;
            reg_file[26414] <= 8'h00;
            reg_file[26415] <= 8'h00;
            reg_file[26416] <= 8'h00;
            reg_file[26417] <= 8'h00;
            reg_file[26418] <= 8'h00;
            reg_file[26419] <= 8'h00;
            reg_file[26420] <= 8'h00;
            reg_file[26421] <= 8'h00;
            reg_file[26422] <= 8'h00;
            reg_file[26423] <= 8'h00;
            reg_file[26424] <= 8'h00;
            reg_file[26425] <= 8'h00;
            reg_file[26426] <= 8'h00;
            reg_file[26427] <= 8'h00;
            reg_file[26428] <= 8'h00;
            reg_file[26429] <= 8'h00;
            reg_file[26430] <= 8'h00;
            reg_file[26431] <= 8'h00;
            reg_file[26432] <= 8'h00;
            reg_file[26433] <= 8'h00;
            reg_file[26434] <= 8'h00;
            reg_file[26435] <= 8'h00;
            reg_file[26436] <= 8'h00;
            reg_file[26437] <= 8'h00;
            reg_file[26438] <= 8'h00;
            reg_file[26439] <= 8'h00;
            reg_file[26440] <= 8'h00;
            reg_file[26441] <= 8'h00;
            reg_file[26442] <= 8'h00;
            reg_file[26443] <= 8'h00;
            reg_file[26444] <= 8'h00;
            reg_file[26445] <= 8'h00;
            reg_file[26446] <= 8'h00;
            reg_file[26447] <= 8'h00;
            reg_file[26448] <= 8'h00;
            reg_file[26449] <= 8'h00;
            reg_file[26450] <= 8'h00;
            reg_file[26451] <= 8'h00;
            reg_file[26452] <= 8'h00;
            reg_file[26453] <= 8'h00;
            reg_file[26454] <= 8'h00;
            reg_file[26455] <= 8'h00;
            reg_file[26456] <= 8'h00;
            reg_file[26457] <= 8'h00;
            reg_file[26458] <= 8'h00;
            reg_file[26459] <= 8'h00;
            reg_file[26460] <= 8'h00;
            reg_file[26461] <= 8'h00;
            reg_file[26462] <= 8'h00;
            reg_file[26463] <= 8'h00;
            reg_file[26464] <= 8'h00;
            reg_file[26465] <= 8'h00;
            reg_file[26466] <= 8'h00;
            reg_file[26467] <= 8'h00;
            reg_file[26468] <= 8'h00;
            reg_file[26469] <= 8'h00;
            reg_file[26470] <= 8'h00;
            reg_file[26471] <= 8'h00;
            reg_file[26472] <= 8'h00;
            reg_file[26473] <= 8'h00;
            reg_file[26474] <= 8'h00;
            reg_file[26475] <= 8'h00;
            reg_file[26476] <= 8'h00;
            reg_file[26477] <= 8'h00;
            reg_file[26478] <= 8'h00;
            reg_file[26479] <= 8'h00;
            reg_file[26480] <= 8'h00;
            reg_file[26481] <= 8'h00;
            reg_file[26482] <= 8'h00;
            reg_file[26483] <= 8'h00;
            reg_file[26484] <= 8'h00;
            reg_file[26485] <= 8'h00;
            reg_file[26486] <= 8'h00;
            reg_file[26487] <= 8'h00;
            reg_file[26488] <= 8'h00;
            reg_file[26489] <= 8'h00;
            reg_file[26490] <= 8'h00;
            reg_file[26491] <= 8'h00;
            reg_file[26492] <= 8'h00;
            reg_file[26493] <= 8'h00;
            reg_file[26494] <= 8'h00;
            reg_file[26495] <= 8'h00;
            reg_file[26496] <= 8'h00;
            reg_file[26497] <= 8'h00;
            reg_file[26498] <= 8'h00;
            reg_file[26499] <= 8'h00;
            reg_file[26500] <= 8'h00;
            reg_file[26501] <= 8'h00;
            reg_file[26502] <= 8'h00;
            reg_file[26503] <= 8'h00;
            reg_file[26504] <= 8'h00;
            reg_file[26505] <= 8'h00;
            reg_file[26506] <= 8'h00;
            reg_file[26507] <= 8'h00;
            reg_file[26508] <= 8'h00;
            reg_file[26509] <= 8'h00;
            reg_file[26510] <= 8'h00;
            reg_file[26511] <= 8'h00;
            reg_file[26512] <= 8'h00;
            reg_file[26513] <= 8'h00;
            reg_file[26514] <= 8'h00;
            reg_file[26515] <= 8'h00;
            reg_file[26516] <= 8'h00;
            reg_file[26517] <= 8'h00;
            reg_file[26518] <= 8'h00;
            reg_file[26519] <= 8'h00;
            reg_file[26520] <= 8'h00;
            reg_file[26521] <= 8'h00;
            reg_file[26522] <= 8'h00;
            reg_file[26523] <= 8'h00;
            reg_file[26524] <= 8'h00;
            reg_file[26525] <= 8'h00;
            reg_file[26526] <= 8'h00;
            reg_file[26527] <= 8'h00;
            reg_file[26528] <= 8'h00;
            reg_file[26529] <= 8'h00;
            reg_file[26530] <= 8'h00;
            reg_file[26531] <= 8'h00;
            reg_file[26532] <= 8'h00;
            reg_file[26533] <= 8'h00;
            reg_file[26534] <= 8'h00;
            reg_file[26535] <= 8'h00;
            reg_file[26536] <= 8'h00;
            reg_file[26537] <= 8'h00;
            reg_file[26538] <= 8'h00;
            reg_file[26539] <= 8'h00;
            reg_file[26540] <= 8'h00;
            reg_file[26541] <= 8'h00;
            reg_file[26542] <= 8'h00;
            reg_file[26543] <= 8'h00;
            reg_file[26544] <= 8'h00;
            reg_file[26545] <= 8'h00;
            reg_file[26546] <= 8'h00;
            reg_file[26547] <= 8'h00;
            reg_file[26548] <= 8'h00;
            reg_file[26549] <= 8'h00;
            reg_file[26550] <= 8'h00;
            reg_file[26551] <= 8'h00;
            reg_file[26552] <= 8'h00;
            reg_file[26553] <= 8'h00;
            reg_file[26554] <= 8'h00;
            reg_file[26555] <= 8'h00;
            reg_file[26556] <= 8'h00;
            reg_file[26557] <= 8'h00;
            reg_file[26558] <= 8'h00;
            reg_file[26559] <= 8'h00;
            reg_file[26560] <= 8'h00;
            reg_file[26561] <= 8'h00;
            reg_file[26562] <= 8'h00;
            reg_file[26563] <= 8'h00;
            reg_file[26564] <= 8'h00;
            reg_file[26565] <= 8'h00;
            reg_file[26566] <= 8'h00;
            reg_file[26567] <= 8'h00;
            reg_file[26568] <= 8'h00;
            reg_file[26569] <= 8'h00;
            reg_file[26570] <= 8'h00;
            reg_file[26571] <= 8'h00;
            reg_file[26572] <= 8'h00;
            reg_file[26573] <= 8'h00;
            reg_file[26574] <= 8'h00;
            reg_file[26575] <= 8'h00;
            reg_file[26576] <= 8'h00;
            reg_file[26577] <= 8'h00;
            reg_file[26578] <= 8'h00;
            reg_file[26579] <= 8'h00;
            reg_file[26580] <= 8'h00;
            reg_file[26581] <= 8'h00;
            reg_file[26582] <= 8'h00;
            reg_file[26583] <= 8'h00;
            reg_file[26584] <= 8'h00;
            reg_file[26585] <= 8'h00;
            reg_file[26586] <= 8'h00;
            reg_file[26587] <= 8'h00;
            reg_file[26588] <= 8'h00;
            reg_file[26589] <= 8'h00;
            reg_file[26590] <= 8'h00;
            reg_file[26591] <= 8'h00;
            reg_file[26592] <= 8'h00;
            reg_file[26593] <= 8'h00;
            reg_file[26594] <= 8'h00;
            reg_file[26595] <= 8'h00;
            reg_file[26596] <= 8'h00;
            reg_file[26597] <= 8'h00;
            reg_file[26598] <= 8'h00;
            reg_file[26599] <= 8'h00;
            reg_file[26600] <= 8'h00;
            reg_file[26601] <= 8'h00;
            reg_file[26602] <= 8'h00;
            reg_file[26603] <= 8'h00;
            reg_file[26604] <= 8'h00;
            reg_file[26605] <= 8'h00;
            reg_file[26606] <= 8'h00;
            reg_file[26607] <= 8'h00;
            reg_file[26608] <= 8'h00;
            reg_file[26609] <= 8'h00;
            reg_file[26610] <= 8'h00;
            reg_file[26611] <= 8'h00;
            reg_file[26612] <= 8'h00;
            reg_file[26613] <= 8'h00;
            reg_file[26614] <= 8'h00;
            reg_file[26615] <= 8'h00;
            reg_file[26616] <= 8'h00;
            reg_file[26617] <= 8'h00;
            reg_file[26618] <= 8'h00;
            reg_file[26619] <= 8'h00;
            reg_file[26620] <= 8'h00;
            reg_file[26621] <= 8'h00;
            reg_file[26622] <= 8'h00;
            reg_file[26623] <= 8'h00;
            reg_file[26624] <= 8'h00;
            reg_file[26625] <= 8'h00;
            reg_file[26626] <= 8'h00;
            reg_file[26627] <= 8'h00;
            reg_file[26628] <= 8'h00;
            reg_file[26629] <= 8'h00;
            reg_file[26630] <= 8'h00;
            reg_file[26631] <= 8'h00;
            reg_file[26632] <= 8'h00;
            reg_file[26633] <= 8'h00;
            reg_file[26634] <= 8'h00;
            reg_file[26635] <= 8'h00;
            reg_file[26636] <= 8'h00;
            reg_file[26637] <= 8'h00;
            reg_file[26638] <= 8'h00;
            reg_file[26639] <= 8'h00;
            reg_file[26640] <= 8'h00;
            reg_file[26641] <= 8'h00;
            reg_file[26642] <= 8'h00;
            reg_file[26643] <= 8'h00;
            reg_file[26644] <= 8'h00;
            reg_file[26645] <= 8'h00;
            reg_file[26646] <= 8'h00;
            reg_file[26647] <= 8'h00;
            reg_file[26648] <= 8'h00;
            reg_file[26649] <= 8'h00;
            reg_file[26650] <= 8'h00;
            reg_file[26651] <= 8'h00;
            reg_file[26652] <= 8'h00;
            reg_file[26653] <= 8'h00;
            reg_file[26654] <= 8'h00;
            reg_file[26655] <= 8'h00;
            reg_file[26656] <= 8'h00;
            reg_file[26657] <= 8'h00;
            reg_file[26658] <= 8'h00;
            reg_file[26659] <= 8'h00;
            reg_file[26660] <= 8'h00;
            reg_file[26661] <= 8'h00;
            reg_file[26662] <= 8'h00;
            reg_file[26663] <= 8'h00;
            reg_file[26664] <= 8'h00;
            reg_file[26665] <= 8'h00;
            reg_file[26666] <= 8'h00;
            reg_file[26667] <= 8'h00;
            reg_file[26668] <= 8'h00;
            reg_file[26669] <= 8'h00;
            reg_file[26670] <= 8'h00;
            reg_file[26671] <= 8'h00;
            reg_file[26672] <= 8'h00;
            reg_file[26673] <= 8'h00;
            reg_file[26674] <= 8'h00;
            reg_file[26675] <= 8'h00;
            reg_file[26676] <= 8'h00;
            reg_file[26677] <= 8'h00;
            reg_file[26678] <= 8'h00;
            reg_file[26679] <= 8'h00;
            reg_file[26680] <= 8'h00;
            reg_file[26681] <= 8'h00;
            reg_file[26682] <= 8'h00;
            reg_file[26683] <= 8'h00;
            reg_file[26684] <= 8'h00;
            reg_file[26685] <= 8'h00;
            reg_file[26686] <= 8'h00;
            reg_file[26687] <= 8'h00;
            reg_file[26688] <= 8'h00;
            reg_file[26689] <= 8'h00;
            reg_file[26690] <= 8'h00;
            reg_file[26691] <= 8'h00;
            reg_file[26692] <= 8'h00;
            reg_file[26693] <= 8'h00;
            reg_file[26694] <= 8'h00;
            reg_file[26695] <= 8'h00;
            reg_file[26696] <= 8'h00;
            reg_file[26697] <= 8'h00;
            reg_file[26698] <= 8'h00;
            reg_file[26699] <= 8'h00;
            reg_file[26700] <= 8'h00;
            reg_file[26701] <= 8'h00;
            reg_file[26702] <= 8'h00;
            reg_file[26703] <= 8'h00;
            reg_file[26704] <= 8'h00;
            reg_file[26705] <= 8'h00;
            reg_file[26706] <= 8'h00;
            reg_file[26707] <= 8'h00;
            reg_file[26708] <= 8'h00;
            reg_file[26709] <= 8'h00;
            reg_file[26710] <= 8'h00;
            reg_file[26711] <= 8'h00;
            reg_file[26712] <= 8'h00;
            reg_file[26713] <= 8'h00;
            reg_file[26714] <= 8'h00;
            reg_file[26715] <= 8'h00;
            reg_file[26716] <= 8'h00;
            reg_file[26717] <= 8'h00;
            reg_file[26718] <= 8'h00;
            reg_file[26719] <= 8'h00;
            reg_file[26720] <= 8'h00;
            reg_file[26721] <= 8'h00;
            reg_file[26722] <= 8'h00;
            reg_file[26723] <= 8'h00;
            reg_file[26724] <= 8'h00;
            reg_file[26725] <= 8'h00;
            reg_file[26726] <= 8'h00;
            reg_file[26727] <= 8'h00;
            reg_file[26728] <= 8'h00;
            reg_file[26729] <= 8'h00;
            reg_file[26730] <= 8'h00;
            reg_file[26731] <= 8'h00;
            reg_file[26732] <= 8'h00;
            reg_file[26733] <= 8'h00;
            reg_file[26734] <= 8'h00;
            reg_file[26735] <= 8'h00;
            reg_file[26736] <= 8'h00;
            reg_file[26737] <= 8'h00;
            reg_file[26738] <= 8'h00;
            reg_file[26739] <= 8'h00;
            reg_file[26740] <= 8'h00;
            reg_file[26741] <= 8'h00;
            reg_file[26742] <= 8'h00;
            reg_file[26743] <= 8'h00;
            reg_file[26744] <= 8'h00;
            reg_file[26745] <= 8'h00;
            reg_file[26746] <= 8'h00;
            reg_file[26747] <= 8'h00;
            reg_file[26748] <= 8'h00;
            reg_file[26749] <= 8'h00;
            reg_file[26750] <= 8'h00;
            reg_file[26751] <= 8'h00;
            reg_file[26752] <= 8'h00;
            reg_file[26753] <= 8'h00;
            reg_file[26754] <= 8'h00;
            reg_file[26755] <= 8'h00;
            reg_file[26756] <= 8'h00;
            reg_file[26757] <= 8'h00;
            reg_file[26758] <= 8'h00;
            reg_file[26759] <= 8'h00;
            reg_file[26760] <= 8'h00;
            reg_file[26761] <= 8'h00;
            reg_file[26762] <= 8'h00;
            reg_file[26763] <= 8'h00;
            reg_file[26764] <= 8'h00;
            reg_file[26765] <= 8'h00;
            reg_file[26766] <= 8'h00;
            reg_file[26767] <= 8'h00;
            reg_file[26768] <= 8'h00;
            reg_file[26769] <= 8'h00;
            reg_file[26770] <= 8'h00;
            reg_file[26771] <= 8'h00;
            reg_file[26772] <= 8'h00;
            reg_file[26773] <= 8'h00;
            reg_file[26774] <= 8'h00;
            reg_file[26775] <= 8'h00;
            reg_file[26776] <= 8'h00;
            reg_file[26777] <= 8'h00;
            reg_file[26778] <= 8'h00;
            reg_file[26779] <= 8'h00;
            reg_file[26780] <= 8'h00;
            reg_file[26781] <= 8'h00;
            reg_file[26782] <= 8'h00;
            reg_file[26783] <= 8'h00;
            reg_file[26784] <= 8'h00;
            reg_file[26785] <= 8'h00;
            reg_file[26786] <= 8'h00;
            reg_file[26787] <= 8'h00;
            reg_file[26788] <= 8'h00;
            reg_file[26789] <= 8'h00;
            reg_file[26790] <= 8'h00;
            reg_file[26791] <= 8'h00;
            reg_file[26792] <= 8'h00;
            reg_file[26793] <= 8'h00;
            reg_file[26794] <= 8'h00;
            reg_file[26795] <= 8'h00;
            reg_file[26796] <= 8'h00;
            reg_file[26797] <= 8'h00;
            reg_file[26798] <= 8'h00;
            reg_file[26799] <= 8'h00;
            reg_file[26800] <= 8'h00;
            reg_file[26801] <= 8'h00;
            reg_file[26802] <= 8'h00;
            reg_file[26803] <= 8'h00;
            reg_file[26804] <= 8'h00;
            reg_file[26805] <= 8'h00;
            reg_file[26806] <= 8'h00;
            reg_file[26807] <= 8'h00;
            reg_file[26808] <= 8'h00;
            reg_file[26809] <= 8'h00;
            reg_file[26810] <= 8'h00;
            reg_file[26811] <= 8'h00;
            reg_file[26812] <= 8'h00;
            reg_file[26813] <= 8'h00;
            reg_file[26814] <= 8'h00;
            reg_file[26815] <= 8'h00;
            reg_file[26816] <= 8'h00;
            reg_file[26817] <= 8'h00;
            reg_file[26818] <= 8'h00;
            reg_file[26819] <= 8'h00;
            reg_file[26820] <= 8'h00;
            reg_file[26821] <= 8'h00;
            reg_file[26822] <= 8'h00;
            reg_file[26823] <= 8'h00;
            reg_file[26824] <= 8'h00;
            reg_file[26825] <= 8'h00;
            reg_file[26826] <= 8'h00;
            reg_file[26827] <= 8'h00;
            reg_file[26828] <= 8'h00;
            reg_file[26829] <= 8'h00;
            reg_file[26830] <= 8'h00;
            reg_file[26831] <= 8'h00;
            reg_file[26832] <= 8'h00;
            reg_file[26833] <= 8'h00;
            reg_file[26834] <= 8'h00;
            reg_file[26835] <= 8'h00;
            reg_file[26836] <= 8'h00;
            reg_file[26837] <= 8'h00;
            reg_file[26838] <= 8'h00;
            reg_file[26839] <= 8'h00;
            reg_file[26840] <= 8'h00;
            reg_file[26841] <= 8'h00;
            reg_file[26842] <= 8'h00;
            reg_file[26843] <= 8'h00;
            reg_file[26844] <= 8'h00;
            reg_file[26845] <= 8'h00;
            reg_file[26846] <= 8'h00;
            reg_file[26847] <= 8'h00;
            reg_file[26848] <= 8'h00;
            reg_file[26849] <= 8'h00;
            reg_file[26850] <= 8'h00;
            reg_file[26851] <= 8'h00;
            reg_file[26852] <= 8'h00;
            reg_file[26853] <= 8'h00;
            reg_file[26854] <= 8'h00;
            reg_file[26855] <= 8'h00;
            reg_file[26856] <= 8'h00;
            reg_file[26857] <= 8'h00;
            reg_file[26858] <= 8'h00;
            reg_file[26859] <= 8'h00;
            reg_file[26860] <= 8'h00;
            reg_file[26861] <= 8'h00;
            reg_file[26862] <= 8'h00;
            reg_file[26863] <= 8'h00;
            reg_file[26864] <= 8'h00;
            reg_file[26865] <= 8'h00;
            reg_file[26866] <= 8'h00;
            reg_file[26867] <= 8'h00;
            reg_file[26868] <= 8'h00;
            reg_file[26869] <= 8'h00;
            reg_file[26870] <= 8'h00;
            reg_file[26871] <= 8'h00;
            reg_file[26872] <= 8'h00;
            reg_file[26873] <= 8'h00;
            reg_file[26874] <= 8'h00;
            reg_file[26875] <= 8'h00;
            reg_file[26876] <= 8'h00;
            reg_file[26877] <= 8'h00;
            reg_file[26878] <= 8'h00;
            reg_file[26879] <= 8'h00;
            reg_file[26880] <= 8'h00;
            reg_file[26881] <= 8'h00;
            reg_file[26882] <= 8'h00;
            reg_file[26883] <= 8'h00;
            reg_file[26884] <= 8'h00;
            reg_file[26885] <= 8'h00;
            reg_file[26886] <= 8'h00;
            reg_file[26887] <= 8'h00;
            reg_file[26888] <= 8'h00;
            reg_file[26889] <= 8'h00;
            reg_file[26890] <= 8'h00;
            reg_file[26891] <= 8'h00;
            reg_file[26892] <= 8'h00;
            reg_file[26893] <= 8'h00;
            reg_file[26894] <= 8'h00;
            reg_file[26895] <= 8'h00;
            reg_file[26896] <= 8'h00;
            reg_file[26897] <= 8'h00;
            reg_file[26898] <= 8'h00;
            reg_file[26899] <= 8'h00;
            reg_file[26900] <= 8'h00;
            reg_file[26901] <= 8'h00;
            reg_file[26902] <= 8'h00;
            reg_file[26903] <= 8'h00;
            reg_file[26904] <= 8'h00;
            reg_file[26905] <= 8'h00;
            reg_file[26906] <= 8'h00;
            reg_file[26907] <= 8'h00;
            reg_file[26908] <= 8'h00;
            reg_file[26909] <= 8'h00;
            reg_file[26910] <= 8'h00;
            reg_file[26911] <= 8'h00;
            reg_file[26912] <= 8'h00;
            reg_file[26913] <= 8'h00;
            reg_file[26914] <= 8'h00;
            reg_file[26915] <= 8'h00;
            reg_file[26916] <= 8'h00;
            reg_file[26917] <= 8'h00;
            reg_file[26918] <= 8'h00;
            reg_file[26919] <= 8'h00;
            reg_file[26920] <= 8'h00;
            reg_file[26921] <= 8'h00;
            reg_file[26922] <= 8'h00;
            reg_file[26923] <= 8'h00;
            reg_file[26924] <= 8'h00;
            reg_file[26925] <= 8'h00;
            reg_file[26926] <= 8'h00;
            reg_file[26927] <= 8'h00;
            reg_file[26928] <= 8'h00;
            reg_file[26929] <= 8'h00;
            reg_file[26930] <= 8'h00;
            reg_file[26931] <= 8'h00;
            reg_file[26932] <= 8'h00;
            reg_file[26933] <= 8'h00;
            reg_file[26934] <= 8'h00;
            reg_file[26935] <= 8'h00;
            reg_file[26936] <= 8'h00;
            reg_file[26937] <= 8'h00;
            reg_file[26938] <= 8'h00;
            reg_file[26939] <= 8'h00;
            reg_file[26940] <= 8'h00;
            reg_file[26941] <= 8'h00;
            reg_file[26942] <= 8'h00;
            reg_file[26943] <= 8'h00;
            reg_file[26944] <= 8'h00;
            reg_file[26945] <= 8'h00;
            reg_file[26946] <= 8'h00;
            reg_file[26947] <= 8'h00;
            reg_file[26948] <= 8'h00;
            reg_file[26949] <= 8'h00;
            reg_file[26950] <= 8'h00;
            reg_file[26951] <= 8'h00;
            reg_file[26952] <= 8'h00;
            reg_file[26953] <= 8'h00;
            reg_file[26954] <= 8'h00;
            reg_file[26955] <= 8'h00;
            reg_file[26956] <= 8'h00;
            reg_file[26957] <= 8'h00;
            reg_file[26958] <= 8'h00;
            reg_file[26959] <= 8'h00;
            reg_file[26960] <= 8'h00;
            reg_file[26961] <= 8'h00;
            reg_file[26962] <= 8'h00;
            reg_file[26963] <= 8'h00;
            reg_file[26964] <= 8'h00;
            reg_file[26965] <= 8'h00;
            reg_file[26966] <= 8'h00;
            reg_file[26967] <= 8'h00;
            reg_file[26968] <= 8'h00;
            reg_file[26969] <= 8'h00;
            reg_file[26970] <= 8'h00;
            reg_file[26971] <= 8'h00;
            reg_file[26972] <= 8'h00;
            reg_file[26973] <= 8'h00;
            reg_file[26974] <= 8'h00;
            reg_file[26975] <= 8'h00;
            reg_file[26976] <= 8'h00;
            reg_file[26977] <= 8'h00;
            reg_file[26978] <= 8'h00;
            reg_file[26979] <= 8'h00;
            reg_file[26980] <= 8'h00;
            reg_file[26981] <= 8'h00;
            reg_file[26982] <= 8'h00;
            reg_file[26983] <= 8'h00;
            reg_file[26984] <= 8'h00;
            reg_file[26985] <= 8'h00;
            reg_file[26986] <= 8'h00;
            reg_file[26987] <= 8'h00;
            reg_file[26988] <= 8'h00;
            reg_file[26989] <= 8'h00;
            reg_file[26990] <= 8'h00;
            reg_file[26991] <= 8'h00;
            reg_file[26992] <= 8'h00;
            reg_file[26993] <= 8'h00;
            reg_file[26994] <= 8'h00;
            reg_file[26995] <= 8'h00;
            reg_file[26996] <= 8'h00;
            reg_file[26997] <= 8'h00;
            reg_file[26998] <= 8'h00;
            reg_file[26999] <= 8'h00;
            reg_file[27000] <= 8'h00;
            reg_file[27001] <= 8'h00;
            reg_file[27002] <= 8'h00;
            reg_file[27003] <= 8'h00;
            reg_file[27004] <= 8'h00;
            reg_file[27005] <= 8'h00;
            reg_file[27006] <= 8'h00;
            reg_file[27007] <= 8'h00;
            reg_file[27008] <= 8'h00;
            reg_file[27009] <= 8'h00;
            reg_file[27010] <= 8'h00;
            reg_file[27011] <= 8'h00;
            reg_file[27012] <= 8'h00;
            reg_file[27013] <= 8'h00;
            reg_file[27014] <= 8'h00;
            reg_file[27015] <= 8'h00;
            reg_file[27016] <= 8'h00;
            reg_file[27017] <= 8'h00;
            reg_file[27018] <= 8'h00;
            reg_file[27019] <= 8'h00;
            reg_file[27020] <= 8'h00;
            reg_file[27021] <= 8'h00;
            reg_file[27022] <= 8'h00;
            reg_file[27023] <= 8'h00;
            reg_file[27024] <= 8'h00;
            reg_file[27025] <= 8'h00;
            reg_file[27026] <= 8'h00;
            reg_file[27027] <= 8'h00;
            reg_file[27028] <= 8'h00;
            reg_file[27029] <= 8'h00;
            reg_file[27030] <= 8'h00;
            reg_file[27031] <= 8'h00;
            reg_file[27032] <= 8'h00;
            reg_file[27033] <= 8'h00;
            reg_file[27034] <= 8'h00;
            reg_file[27035] <= 8'h00;
            reg_file[27036] <= 8'h00;
            reg_file[27037] <= 8'h00;
            reg_file[27038] <= 8'h00;
            reg_file[27039] <= 8'h00;
            reg_file[27040] <= 8'h00;
            reg_file[27041] <= 8'h00;
            reg_file[27042] <= 8'h00;
            reg_file[27043] <= 8'h00;
            reg_file[27044] <= 8'h00;
            reg_file[27045] <= 8'h00;
            reg_file[27046] <= 8'h00;
            reg_file[27047] <= 8'h00;
            reg_file[27048] <= 8'h00;
            reg_file[27049] <= 8'h00;
            reg_file[27050] <= 8'h00;
            reg_file[27051] <= 8'h00;
            reg_file[27052] <= 8'h00;
            reg_file[27053] <= 8'h00;
            reg_file[27054] <= 8'h00;
            reg_file[27055] <= 8'h00;
            reg_file[27056] <= 8'h00;
            reg_file[27057] <= 8'h00;
            reg_file[27058] <= 8'h00;
            reg_file[27059] <= 8'h00;
            reg_file[27060] <= 8'h00;
            reg_file[27061] <= 8'h00;
            reg_file[27062] <= 8'h00;
            reg_file[27063] <= 8'h00;
            reg_file[27064] <= 8'h00;
            reg_file[27065] <= 8'h00;
            reg_file[27066] <= 8'h00;
            reg_file[27067] <= 8'h00;
            reg_file[27068] <= 8'h00;
            reg_file[27069] <= 8'h00;
            reg_file[27070] <= 8'h00;
            reg_file[27071] <= 8'h00;
            reg_file[27072] <= 8'h00;
            reg_file[27073] <= 8'h00;
            reg_file[27074] <= 8'h00;
            reg_file[27075] <= 8'h00;
            reg_file[27076] <= 8'h00;
            reg_file[27077] <= 8'h00;
            reg_file[27078] <= 8'h00;
            reg_file[27079] <= 8'h00;
            reg_file[27080] <= 8'h00;
            reg_file[27081] <= 8'h00;
            reg_file[27082] <= 8'h00;
            reg_file[27083] <= 8'h00;
            reg_file[27084] <= 8'h00;
            reg_file[27085] <= 8'h00;
            reg_file[27086] <= 8'h00;
            reg_file[27087] <= 8'h00;
            reg_file[27088] <= 8'h00;
            reg_file[27089] <= 8'h00;
            reg_file[27090] <= 8'h00;
            reg_file[27091] <= 8'h00;
            reg_file[27092] <= 8'h00;
            reg_file[27093] <= 8'h00;
            reg_file[27094] <= 8'h00;
            reg_file[27095] <= 8'h00;
            reg_file[27096] <= 8'h00;
            reg_file[27097] <= 8'h00;
            reg_file[27098] <= 8'h00;
            reg_file[27099] <= 8'h00;
            reg_file[27100] <= 8'h00;
            reg_file[27101] <= 8'h00;
            reg_file[27102] <= 8'h00;
            reg_file[27103] <= 8'h00;
            reg_file[27104] <= 8'h00;
            reg_file[27105] <= 8'h00;
            reg_file[27106] <= 8'h00;
            reg_file[27107] <= 8'h00;
            reg_file[27108] <= 8'h00;
            reg_file[27109] <= 8'h00;
            reg_file[27110] <= 8'h00;
            reg_file[27111] <= 8'h00;
            reg_file[27112] <= 8'h00;
            reg_file[27113] <= 8'h00;
            reg_file[27114] <= 8'h00;
            reg_file[27115] <= 8'h00;
            reg_file[27116] <= 8'h00;
            reg_file[27117] <= 8'h00;
            reg_file[27118] <= 8'h00;
            reg_file[27119] <= 8'h00;
            reg_file[27120] <= 8'h00;
            reg_file[27121] <= 8'h00;
            reg_file[27122] <= 8'h00;
            reg_file[27123] <= 8'h00;
            reg_file[27124] <= 8'h00;
            reg_file[27125] <= 8'h00;
            reg_file[27126] <= 8'h00;
            reg_file[27127] <= 8'h00;
            reg_file[27128] <= 8'h00;
            reg_file[27129] <= 8'h00;
            reg_file[27130] <= 8'h00;
            reg_file[27131] <= 8'h00;
            reg_file[27132] <= 8'h00;
            reg_file[27133] <= 8'h00;
            reg_file[27134] <= 8'h00;
            reg_file[27135] <= 8'h00;
            reg_file[27136] <= 8'h00;
            reg_file[27137] <= 8'h00;
            reg_file[27138] <= 8'h00;
            reg_file[27139] <= 8'h00;
            reg_file[27140] <= 8'h00;
            reg_file[27141] <= 8'h00;
            reg_file[27142] <= 8'h00;
            reg_file[27143] <= 8'h00;
            reg_file[27144] <= 8'h00;
            reg_file[27145] <= 8'h00;
            reg_file[27146] <= 8'h00;
            reg_file[27147] <= 8'h00;
            reg_file[27148] <= 8'h00;
            reg_file[27149] <= 8'h00;
            reg_file[27150] <= 8'h00;
            reg_file[27151] <= 8'h00;
            reg_file[27152] <= 8'h00;
            reg_file[27153] <= 8'h00;
            reg_file[27154] <= 8'h00;
            reg_file[27155] <= 8'h00;
            reg_file[27156] <= 8'h00;
            reg_file[27157] <= 8'h00;
            reg_file[27158] <= 8'h00;
            reg_file[27159] <= 8'h00;
            reg_file[27160] <= 8'h00;
            reg_file[27161] <= 8'h00;
            reg_file[27162] <= 8'h00;
            reg_file[27163] <= 8'h00;
            reg_file[27164] <= 8'h00;
            reg_file[27165] <= 8'h00;
            reg_file[27166] <= 8'h00;
            reg_file[27167] <= 8'h00;
            reg_file[27168] <= 8'h00;
            reg_file[27169] <= 8'h00;
            reg_file[27170] <= 8'h00;
            reg_file[27171] <= 8'h00;
            reg_file[27172] <= 8'h00;
            reg_file[27173] <= 8'h00;
            reg_file[27174] <= 8'h00;
            reg_file[27175] <= 8'h00;
            reg_file[27176] <= 8'h00;
            reg_file[27177] <= 8'h00;
            reg_file[27178] <= 8'h00;
            reg_file[27179] <= 8'h00;
            reg_file[27180] <= 8'h00;
            reg_file[27181] <= 8'h00;
            reg_file[27182] <= 8'h00;
            reg_file[27183] <= 8'h00;
            reg_file[27184] <= 8'h00;
            reg_file[27185] <= 8'h00;
            reg_file[27186] <= 8'h00;
            reg_file[27187] <= 8'h00;
            reg_file[27188] <= 8'h00;
            reg_file[27189] <= 8'h00;
            reg_file[27190] <= 8'h00;
            reg_file[27191] <= 8'h00;
            reg_file[27192] <= 8'h00;
            reg_file[27193] <= 8'h00;
            reg_file[27194] <= 8'h00;
            reg_file[27195] <= 8'h00;
            reg_file[27196] <= 8'h00;
            reg_file[27197] <= 8'h00;
            reg_file[27198] <= 8'h00;
            reg_file[27199] <= 8'h00;
            reg_file[27200] <= 8'h00;
            reg_file[27201] <= 8'h00;
            reg_file[27202] <= 8'h00;
            reg_file[27203] <= 8'h00;
            reg_file[27204] <= 8'h00;
            reg_file[27205] <= 8'h00;
            reg_file[27206] <= 8'h00;
            reg_file[27207] <= 8'h00;
            reg_file[27208] <= 8'h00;
            reg_file[27209] <= 8'h00;
            reg_file[27210] <= 8'h00;
            reg_file[27211] <= 8'h00;
            reg_file[27212] <= 8'h00;
            reg_file[27213] <= 8'h00;
            reg_file[27214] <= 8'h00;
            reg_file[27215] <= 8'h00;
            reg_file[27216] <= 8'h00;
            reg_file[27217] <= 8'h00;
            reg_file[27218] <= 8'h00;
            reg_file[27219] <= 8'h00;
            reg_file[27220] <= 8'h00;
            reg_file[27221] <= 8'h00;
            reg_file[27222] <= 8'h00;
            reg_file[27223] <= 8'h00;
            reg_file[27224] <= 8'h00;
            reg_file[27225] <= 8'h00;
            reg_file[27226] <= 8'h00;
            reg_file[27227] <= 8'h00;
            reg_file[27228] <= 8'h00;
            reg_file[27229] <= 8'h00;
            reg_file[27230] <= 8'h00;
            reg_file[27231] <= 8'h00;
            reg_file[27232] <= 8'h00;
            reg_file[27233] <= 8'h00;
            reg_file[27234] <= 8'h00;
            reg_file[27235] <= 8'h00;
            reg_file[27236] <= 8'h00;
            reg_file[27237] <= 8'h00;
            reg_file[27238] <= 8'h00;
            reg_file[27239] <= 8'h00;
            reg_file[27240] <= 8'h00;
            reg_file[27241] <= 8'h00;
            reg_file[27242] <= 8'h00;
            reg_file[27243] <= 8'h00;
            reg_file[27244] <= 8'h00;
            reg_file[27245] <= 8'h00;
            reg_file[27246] <= 8'h00;
            reg_file[27247] <= 8'h00;
            reg_file[27248] <= 8'h00;
            reg_file[27249] <= 8'h00;
            reg_file[27250] <= 8'h00;
            reg_file[27251] <= 8'h00;
            reg_file[27252] <= 8'h00;
            reg_file[27253] <= 8'h00;
            reg_file[27254] <= 8'h00;
            reg_file[27255] <= 8'h00;
            reg_file[27256] <= 8'h00;
            reg_file[27257] <= 8'h00;
            reg_file[27258] <= 8'h00;
            reg_file[27259] <= 8'h00;
            reg_file[27260] <= 8'h00;
            reg_file[27261] <= 8'h00;
            reg_file[27262] <= 8'h00;
            reg_file[27263] <= 8'h00;
            reg_file[27264] <= 8'h00;
            reg_file[27265] <= 8'h00;
            reg_file[27266] <= 8'h00;
            reg_file[27267] <= 8'h00;
            reg_file[27268] <= 8'h00;
            reg_file[27269] <= 8'h00;
            reg_file[27270] <= 8'h00;
            reg_file[27271] <= 8'h00;
            reg_file[27272] <= 8'h00;
            reg_file[27273] <= 8'h00;
            reg_file[27274] <= 8'h00;
            reg_file[27275] <= 8'h00;
            reg_file[27276] <= 8'h00;
            reg_file[27277] <= 8'h00;
            reg_file[27278] <= 8'h00;
            reg_file[27279] <= 8'h00;
            reg_file[27280] <= 8'h00;
            reg_file[27281] <= 8'h00;
            reg_file[27282] <= 8'h00;
            reg_file[27283] <= 8'h00;
            reg_file[27284] <= 8'h00;
            reg_file[27285] <= 8'h00;
            reg_file[27286] <= 8'h00;
            reg_file[27287] <= 8'h00;
            reg_file[27288] <= 8'h00;
            reg_file[27289] <= 8'h00;
            reg_file[27290] <= 8'h00;
            reg_file[27291] <= 8'h00;
            reg_file[27292] <= 8'h00;
            reg_file[27293] <= 8'h00;
            reg_file[27294] <= 8'h00;
            reg_file[27295] <= 8'h00;
            reg_file[27296] <= 8'h00;
            reg_file[27297] <= 8'h00;
            reg_file[27298] <= 8'h00;
            reg_file[27299] <= 8'h00;
            reg_file[27300] <= 8'h00;
            reg_file[27301] <= 8'h00;
            reg_file[27302] <= 8'h00;
            reg_file[27303] <= 8'h00;
            reg_file[27304] <= 8'h00;
            reg_file[27305] <= 8'h00;
            reg_file[27306] <= 8'h00;
            reg_file[27307] <= 8'h00;
            reg_file[27308] <= 8'h00;
            reg_file[27309] <= 8'h00;
            reg_file[27310] <= 8'h00;
            reg_file[27311] <= 8'h00;
            reg_file[27312] <= 8'h00;
            reg_file[27313] <= 8'h00;
            reg_file[27314] <= 8'h00;
            reg_file[27315] <= 8'h00;
            reg_file[27316] <= 8'h00;
            reg_file[27317] <= 8'h00;
            reg_file[27318] <= 8'h00;
            reg_file[27319] <= 8'h00;
            reg_file[27320] <= 8'h00;
            reg_file[27321] <= 8'h00;
            reg_file[27322] <= 8'h00;
            reg_file[27323] <= 8'h00;
            reg_file[27324] <= 8'h00;
            reg_file[27325] <= 8'h00;
            reg_file[27326] <= 8'h00;
            reg_file[27327] <= 8'h00;
            reg_file[27328] <= 8'h00;
            reg_file[27329] <= 8'h00;
            reg_file[27330] <= 8'h00;
            reg_file[27331] <= 8'h00;
            reg_file[27332] <= 8'h00;
            reg_file[27333] <= 8'h00;
            reg_file[27334] <= 8'h00;
            reg_file[27335] <= 8'h00;
            reg_file[27336] <= 8'h00;
            reg_file[27337] <= 8'h00;
            reg_file[27338] <= 8'h00;
            reg_file[27339] <= 8'h00;
            reg_file[27340] <= 8'h00;
            reg_file[27341] <= 8'h00;
            reg_file[27342] <= 8'h00;
            reg_file[27343] <= 8'h00;
            reg_file[27344] <= 8'h00;
            reg_file[27345] <= 8'h00;
            reg_file[27346] <= 8'h00;
            reg_file[27347] <= 8'h00;
            reg_file[27348] <= 8'h00;
            reg_file[27349] <= 8'h00;
            reg_file[27350] <= 8'h00;
            reg_file[27351] <= 8'h00;
            reg_file[27352] <= 8'h00;
            reg_file[27353] <= 8'h00;
            reg_file[27354] <= 8'h00;
            reg_file[27355] <= 8'h00;
            reg_file[27356] <= 8'h00;
            reg_file[27357] <= 8'h00;
            reg_file[27358] <= 8'h00;
            reg_file[27359] <= 8'h00;
            reg_file[27360] <= 8'h00;
            reg_file[27361] <= 8'h00;
            reg_file[27362] <= 8'h00;
            reg_file[27363] <= 8'h00;
            reg_file[27364] <= 8'h00;
            reg_file[27365] <= 8'h00;
            reg_file[27366] <= 8'h00;
            reg_file[27367] <= 8'h00;
            reg_file[27368] <= 8'h00;
            reg_file[27369] <= 8'h00;
            reg_file[27370] <= 8'h00;
            reg_file[27371] <= 8'h00;
            reg_file[27372] <= 8'h00;
            reg_file[27373] <= 8'h00;
            reg_file[27374] <= 8'h00;
            reg_file[27375] <= 8'h00;
            reg_file[27376] <= 8'h00;
            reg_file[27377] <= 8'h00;
            reg_file[27378] <= 8'h00;
            reg_file[27379] <= 8'h00;
            reg_file[27380] <= 8'h00;
            reg_file[27381] <= 8'h00;
            reg_file[27382] <= 8'h00;
            reg_file[27383] <= 8'h00;
            reg_file[27384] <= 8'h00;
            reg_file[27385] <= 8'h00;
            reg_file[27386] <= 8'h00;
            reg_file[27387] <= 8'h00;
            reg_file[27388] <= 8'h00;
            reg_file[27389] <= 8'h00;
            reg_file[27390] <= 8'h00;
            reg_file[27391] <= 8'h00;
            reg_file[27392] <= 8'h00;
            reg_file[27393] <= 8'h00;
            reg_file[27394] <= 8'h00;
            reg_file[27395] <= 8'h00;
            reg_file[27396] <= 8'h00;
            reg_file[27397] <= 8'h00;
            reg_file[27398] <= 8'h00;
            reg_file[27399] <= 8'h00;
            reg_file[27400] <= 8'h00;
            reg_file[27401] <= 8'h00;
            reg_file[27402] <= 8'h00;
            reg_file[27403] <= 8'h00;
            reg_file[27404] <= 8'h00;
            reg_file[27405] <= 8'h00;
            reg_file[27406] <= 8'h00;
            reg_file[27407] <= 8'h00;
            reg_file[27408] <= 8'h00;
            reg_file[27409] <= 8'h00;
            reg_file[27410] <= 8'h00;
            reg_file[27411] <= 8'h00;
            reg_file[27412] <= 8'h00;
            reg_file[27413] <= 8'h00;
            reg_file[27414] <= 8'h00;
            reg_file[27415] <= 8'h00;
            reg_file[27416] <= 8'h00;
            reg_file[27417] <= 8'h00;
            reg_file[27418] <= 8'h00;
            reg_file[27419] <= 8'h00;
            reg_file[27420] <= 8'h00;
            reg_file[27421] <= 8'h00;
            reg_file[27422] <= 8'h00;
            reg_file[27423] <= 8'h00;
            reg_file[27424] <= 8'h00;
            reg_file[27425] <= 8'h00;
            reg_file[27426] <= 8'h00;
            reg_file[27427] <= 8'h00;
            reg_file[27428] <= 8'h00;
            reg_file[27429] <= 8'h00;
            reg_file[27430] <= 8'h00;
            reg_file[27431] <= 8'h00;
            reg_file[27432] <= 8'h00;
            reg_file[27433] <= 8'h00;
            reg_file[27434] <= 8'h00;
            reg_file[27435] <= 8'h00;
            reg_file[27436] <= 8'h00;
            reg_file[27437] <= 8'h00;
            reg_file[27438] <= 8'h00;
            reg_file[27439] <= 8'h00;
            reg_file[27440] <= 8'h00;
            reg_file[27441] <= 8'h00;
            reg_file[27442] <= 8'h00;
            reg_file[27443] <= 8'h00;
            reg_file[27444] <= 8'h00;
            reg_file[27445] <= 8'h00;
            reg_file[27446] <= 8'h00;
            reg_file[27447] <= 8'h00;
            reg_file[27448] <= 8'h00;
            reg_file[27449] <= 8'h00;
            reg_file[27450] <= 8'h00;
            reg_file[27451] <= 8'h00;
            reg_file[27452] <= 8'h00;
            reg_file[27453] <= 8'h00;
            reg_file[27454] <= 8'h00;
            reg_file[27455] <= 8'h00;
            reg_file[27456] <= 8'h00;
            reg_file[27457] <= 8'h00;
            reg_file[27458] <= 8'h00;
            reg_file[27459] <= 8'h00;
            reg_file[27460] <= 8'h00;
            reg_file[27461] <= 8'h00;
            reg_file[27462] <= 8'h00;
            reg_file[27463] <= 8'h00;
            reg_file[27464] <= 8'h00;
            reg_file[27465] <= 8'h00;
            reg_file[27466] <= 8'h00;
            reg_file[27467] <= 8'h00;
            reg_file[27468] <= 8'h00;
            reg_file[27469] <= 8'h00;
            reg_file[27470] <= 8'h00;
            reg_file[27471] <= 8'h00;
            reg_file[27472] <= 8'h00;
            reg_file[27473] <= 8'h00;
            reg_file[27474] <= 8'h00;
            reg_file[27475] <= 8'h00;
            reg_file[27476] <= 8'h00;
            reg_file[27477] <= 8'h00;
            reg_file[27478] <= 8'h00;
            reg_file[27479] <= 8'h00;
            reg_file[27480] <= 8'h00;
            reg_file[27481] <= 8'h00;
            reg_file[27482] <= 8'h00;
            reg_file[27483] <= 8'h00;
            reg_file[27484] <= 8'h00;
            reg_file[27485] <= 8'h00;
            reg_file[27486] <= 8'h00;
            reg_file[27487] <= 8'h00;
            reg_file[27488] <= 8'h00;
            reg_file[27489] <= 8'h00;
            reg_file[27490] <= 8'h00;
            reg_file[27491] <= 8'h00;
            reg_file[27492] <= 8'h00;
            reg_file[27493] <= 8'h00;
            reg_file[27494] <= 8'h00;
            reg_file[27495] <= 8'h00;
            reg_file[27496] <= 8'h00;
            reg_file[27497] <= 8'h00;
            reg_file[27498] <= 8'h00;
            reg_file[27499] <= 8'h00;
            reg_file[27500] <= 8'h00;
            reg_file[27501] <= 8'h00;
            reg_file[27502] <= 8'h00;
            reg_file[27503] <= 8'h00;
            reg_file[27504] <= 8'h00;
            reg_file[27505] <= 8'h00;
            reg_file[27506] <= 8'h00;
            reg_file[27507] <= 8'h00;
            reg_file[27508] <= 8'h00;
            reg_file[27509] <= 8'h00;
            reg_file[27510] <= 8'h00;
            reg_file[27511] <= 8'h00;
            reg_file[27512] <= 8'h00;
            reg_file[27513] <= 8'h00;
            reg_file[27514] <= 8'h00;
            reg_file[27515] <= 8'h00;
            reg_file[27516] <= 8'h00;
            reg_file[27517] <= 8'h00;
            reg_file[27518] <= 8'h00;
            reg_file[27519] <= 8'h00;
            reg_file[27520] <= 8'h00;
            reg_file[27521] <= 8'h00;
            reg_file[27522] <= 8'h00;
            reg_file[27523] <= 8'h00;
            reg_file[27524] <= 8'h00;
            reg_file[27525] <= 8'h00;
            reg_file[27526] <= 8'h00;
            reg_file[27527] <= 8'h00;
            reg_file[27528] <= 8'h00;
            reg_file[27529] <= 8'h00;
            reg_file[27530] <= 8'h00;
            reg_file[27531] <= 8'h00;
            reg_file[27532] <= 8'h00;
            reg_file[27533] <= 8'h00;
            reg_file[27534] <= 8'h00;
            reg_file[27535] <= 8'h00;
            reg_file[27536] <= 8'h00;
            reg_file[27537] <= 8'h00;
            reg_file[27538] <= 8'h00;
            reg_file[27539] <= 8'h00;
            reg_file[27540] <= 8'h00;
            reg_file[27541] <= 8'h00;
            reg_file[27542] <= 8'h00;
            reg_file[27543] <= 8'h00;
            reg_file[27544] <= 8'h00;
            reg_file[27545] <= 8'h00;
            reg_file[27546] <= 8'h00;
            reg_file[27547] <= 8'h00;
            reg_file[27548] <= 8'h00;
            reg_file[27549] <= 8'h00;
            reg_file[27550] <= 8'h00;
            reg_file[27551] <= 8'h00;
            reg_file[27552] <= 8'h00;
            reg_file[27553] <= 8'h00;
            reg_file[27554] <= 8'h00;
            reg_file[27555] <= 8'h00;
            reg_file[27556] <= 8'h00;
            reg_file[27557] <= 8'h00;
            reg_file[27558] <= 8'h00;
            reg_file[27559] <= 8'h00;
            reg_file[27560] <= 8'h00;
            reg_file[27561] <= 8'h00;
            reg_file[27562] <= 8'h00;
            reg_file[27563] <= 8'h00;
            reg_file[27564] <= 8'h00;
            reg_file[27565] <= 8'h00;
            reg_file[27566] <= 8'h00;
            reg_file[27567] <= 8'h00;
            reg_file[27568] <= 8'h00;
            reg_file[27569] <= 8'h00;
            reg_file[27570] <= 8'h00;
            reg_file[27571] <= 8'h00;
            reg_file[27572] <= 8'h00;
            reg_file[27573] <= 8'h00;
            reg_file[27574] <= 8'h00;
            reg_file[27575] <= 8'h00;
            reg_file[27576] <= 8'h00;
            reg_file[27577] <= 8'h00;
            reg_file[27578] <= 8'h00;
            reg_file[27579] <= 8'h00;
            reg_file[27580] <= 8'h00;
            reg_file[27581] <= 8'h00;
            reg_file[27582] <= 8'h00;
            reg_file[27583] <= 8'h00;
            reg_file[27584] <= 8'h00;
            reg_file[27585] <= 8'h00;
            reg_file[27586] <= 8'h00;
            reg_file[27587] <= 8'h00;
            reg_file[27588] <= 8'h00;
            reg_file[27589] <= 8'h00;
            reg_file[27590] <= 8'h00;
            reg_file[27591] <= 8'h00;
            reg_file[27592] <= 8'h00;
            reg_file[27593] <= 8'h00;
            reg_file[27594] <= 8'h00;
            reg_file[27595] <= 8'h00;
            reg_file[27596] <= 8'h00;
            reg_file[27597] <= 8'h00;
            reg_file[27598] <= 8'h00;
            reg_file[27599] <= 8'h00;
            reg_file[27600] <= 8'h00;
            reg_file[27601] <= 8'h00;
            reg_file[27602] <= 8'h00;
            reg_file[27603] <= 8'h00;
            reg_file[27604] <= 8'h00;
            reg_file[27605] <= 8'h00;
            reg_file[27606] <= 8'h00;
            reg_file[27607] <= 8'h00;
            reg_file[27608] <= 8'h00;
            reg_file[27609] <= 8'h00;
            reg_file[27610] <= 8'h00;
            reg_file[27611] <= 8'h00;
            reg_file[27612] <= 8'h00;
            reg_file[27613] <= 8'h00;
            reg_file[27614] <= 8'h00;
            reg_file[27615] <= 8'h00;
            reg_file[27616] <= 8'h00;
            reg_file[27617] <= 8'h00;
            reg_file[27618] <= 8'h00;
            reg_file[27619] <= 8'h00;
            reg_file[27620] <= 8'h00;
            reg_file[27621] <= 8'h00;
            reg_file[27622] <= 8'h00;
            reg_file[27623] <= 8'h00;
            reg_file[27624] <= 8'h00;
            reg_file[27625] <= 8'h00;
            reg_file[27626] <= 8'h00;
            reg_file[27627] <= 8'h00;
            reg_file[27628] <= 8'h00;
            reg_file[27629] <= 8'h00;
            reg_file[27630] <= 8'h00;
            reg_file[27631] <= 8'h00;
            reg_file[27632] <= 8'h00;
            reg_file[27633] <= 8'h00;
            reg_file[27634] <= 8'h00;
            reg_file[27635] <= 8'h00;
            reg_file[27636] <= 8'h00;
            reg_file[27637] <= 8'h00;
            reg_file[27638] <= 8'h00;
            reg_file[27639] <= 8'h00;
            reg_file[27640] <= 8'h00;
            reg_file[27641] <= 8'h00;
            reg_file[27642] <= 8'h00;
            reg_file[27643] <= 8'h00;
            reg_file[27644] <= 8'h00;
            reg_file[27645] <= 8'h00;
            reg_file[27646] <= 8'h00;
            reg_file[27647] <= 8'h00;
            reg_file[27648] <= 8'h00;
            reg_file[27649] <= 8'h00;
            reg_file[27650] <= 8'h00;
            reg_file[27651] <= 8'h00;
            reg_file[27652] <= 8'h00;
            reg_file[27653] <= 8'h00;
            reg_file[27654] <= 8'h00;
            reg_file[27655] <= 8'h00;
            reg_file[27656] <= 8'h00;
            reg_file[27657] <= 8'h00;
            reg_file[27658] <= 8'h00;
            reg_file[27659] <= 8'h00;
            reg_file[27660] <= 8'h00;
            reg_file[27661] <= 8'h00;
            reg_file[27662] <= 8'h00;
            reg_file[27663] <= 8'h00;
            reg_file[27664] <= 8'h00;
            reg_file[27665] <= 8'h00;
            reg_file[27666] <= 8'h00;
            reg_file[27667] <= 8'h00;
            reg_file[27668] <= 8'h00;
            reg_file[27669] <= 8'h00;
            reg_file[27670] <= 8'h00;
            reg_file[27671] <= 8'h00;
            reg_file[27672] <= 8'h00;
            reg_file[27673] <= 8'h00;
            reg_file[27674] <= 8'h00;
            reg_file[27675] <= 8'h00;
            reg_file[27676] <= 8'h00;
            reg_file[27677] <= 8'h00;
            reg_file[27678] <= 8'h00;
            reg_file[27679] <= 8'h00;
            reg_file[27680] <= 8'h00;
            reg_file[27681] <= 8'h00;
            reg_file[27682] <= 8'h00;
            reg_file[27683] <= 8'h00;
            reg_file[27684] <= 8'h00;
            reg_file[27685] <= 8'h00;
            reg_file[27686] <= 8'h00;
            reg_file[27687] <= 8'h00;
            reg_file[27688] <= 8'h00;
            reg_file[27689] <= 8'h00;
            reg_file[27690] <= 8'h00;
            reg_file[27691] <= 8'h00;
            reg_file[27692] <= 8'h00;
            reg_file[27693] <= 8'h00;
            reg_file[27694] <= 8'h00;
            reg_file[27695] <= 8'h00;
            reg_file[27696] <= 8'h00;
            reg_file[27697] <= 8'h00;
            reg_file[27698] <= 8'h00;
            reg_file[27699] <= 8'h00;
            reg_file[27700] <= 8'h00;
            reg_file[27701] <= 8'h00;
            reg_file[27702] <= 8'h00;
            reg_file[27703] <= 8'h00;
            reg_file[27704] <= 8'h00;
            reg_file[27705] <= 8'h00;
            reg_file[27706] <= 8'h00;
            reg_file[27707] <= 8'h00;
            reg_file[27708] <= 8'h00;
            reg_file[27709] <= 8'h00;
            reg_file[27710] <= 8'h00;
            reg_file[27711] <= 8'h00;
            reg_file[27712] <= 8'h00;
            reg_file[27713] <= 8'h00;
            reg_file[27714] <= 8'h00;
            reg_file[27715] <= 8'h00;
            reg_file[27716] <= 8'h00;
            reg_file[27717] <= 8'h00;
            reg_file[27718] <= 8'h00;
            reg_file[27719] <= 8'h00;
            reg_file[27720] <= 8'h00;
            reg_file[27721] <= 8'h00;
            reg_file[27722] <= 8'h00;
            reg_file[27723] <= 8'h00;
            reg_file[27724] <= 8'h00;
            reg_file[27725] <= 8'h00;
            reg_file[27726] <= 8'h00;
            reg_file[27727] <= 8'h00;
            reg_file[27728] <= 8'h00;
            reg_file[27729] <= 8'h00;
            reg_file[27730] <= 8'h00;
            reg_file[27731] <= 8'h00;
            reg_file[27732] <= 8'h00;
            reg_file[27733] <= 8'h00;
            reg_file[27734] <= 8'h00;
            reg_file[27735] <= 8'h00;
            reg_file[27736] <= 8'h00;
            reg_file[27737] <= 8'h00;
            reg_file[27738] <= 8'h00;
            reg_file[27739] <= 8'h00;
            reg_file[27740] <= 8'h00;
            reg_file[27741] <= 8'h00;
            reg_file[27742] <= 8'h00;
            reg_file[27743] <= 8'h00;
            reg_file[27744] <= 8'h00;
            reg_file[27745] <= 8'h00;
            reg_file[27746] <= 8'h00;
            reg_file[27747] <= 8'h00;
            reg_file[27748] <= 8'h00;
            reg_file[27749] <= 8'h00;
            reg_file[27750] <= 8'h00;
            reg_file[27751] <= 8'h00;
            reg_file[27752] <= 8'h00;
            reg_file[27753] <= 8'h00;
            reg_file[27754] <= 8'h00;
            reg_file[27755] <= 8'h00;
            reg_file[27756] <= 8'h00;
            reg_file[27757] <= 8'h00;
            reg_file[27758] <= 8'h00;
            reg_file[27759] <= 8'h00;
            reg_file[27760] <= 8'h00;
            reg_file[27761] <= 8'h00;
            reg_file[27762] <= 8'h00;
            reg_file[27763] <= 8'h00;
            reg_file[27764] <= 8'h00;
            reg_file[27765] <= 8'h00;
            reg_file[27766] <= 8'h00;
            reg_file[27767] <= 8'h00;
            reg_file[27768] <= 8'h00;
            reg_file[27769] <= 8'h00;
            reg_file[27770] <= 8'h00;
            reg_file[27771] <= 8'h00;
            reg_file[27772] <= 8'h00;
            reg_file[27773] <= 8'h00;
            reg_file[27774] <= 8'h00;
            reg_file[27775] <= 8'h00;
            reg_file[27776] <= 8'h00;
            reg_file[27777] <= 8'h00;
            reg_file[27778] <= 8'h00;
            reg_file[27779] <= 8'h00;
            reg_file[27780] <= 8'h00;
            reg_file[27781] <= 8'h00;
            reg_file[27782] <= 8'h00;
            reg_file[27783] <= 8'h00;
            reg_file[27784] <= 8'h00;
            reg_file[27785] <= 8'h00;
            reg_file[27786] <= 8'h00;
            reg_file[27787] <= 8'h00;
            reg_file[27788] <= 8'h00;
            reg_file[27789] <= 8'h00;
            reg_file[27790] <= 8'h00;
            reg_file[27791] <= 8'h00;
            reg_file[27792] <= 8'h00;
            reg_file[27793] <= 8'h00;
            reg_file[27794] <= 8'h00;
            reg_file[27795] <= 8'h00;
            reg_file[27796] <= 8'h00;
            reg_file[27797] <= 8'h00;
            reg_file[27798] <= 8'h00;
            reg_file[27799] <= 8'h00;
            reg_file[27800] <= 8'h00;
            reg_file[27801] <= 8'h00;
            reg_file[27802] <= 8'h00;
            reg_file[27803] <= 8'h00;
            reg_file[27804] <= 8'h00;
            reg_file[27805] <= 8'h00;
            reg_file[27806] <= 8'h00;
            reg_file[27807] <= 8'h00;
            reg_file[27808] <= 8'h00;
            reg_file[27809] <= 8'h00;
            reg_file[27810] <= 8'h00;
            reg_file[27811] <= 8'h00;
            reg_file[27812] <= 8'h00;
            reg_file[27813] <= 8'h00;
            reg_file[27814] <= 8'h00;
            reg_file[27815] <= 8'h00;
            reg_file[27816] <= 8'h00;
            reg_file[27817] <= 8'h00;
            reg_file[27818] <= 8'h00;
            reg_file[27819] <= 8'h00;
            reg_file[27820] <= 8'h00;
            reg_file[27821] <= 8'h00;
            reg_file[27822] <= 8'h00;
            reg_file[27823] <= 8'h00;
            reg_file[27824] <= 8'h00;
            reg_file[27825] <= 8'h00;
            reg_file[27826] <= 8'h00;
            reg_file[27827] <= 8'h00;
            reg_file[27828] <= 8'h00;
            reg_file[27829] <= 8'h00;
            reg_file[27830] <= 8'h00;
            reg_file[27831] <= 8'h00;
            reg_file[27832] <= 8'h00;
            reg_file[27833] <= 8'h00;
            reg_file[27834] <= 8'h00;
            reg_file[27835] <= 8'h00;
            reg_file[27836] <= 8'h00;
            reg_file[27837] <= 8'h00;
            reg_file[27838] <= 8'h00;
            reg_file[27839] <= 8'h00;
            reg_file[27840] <= 8'h00;
            reg_file[27841] <= 8'h00;
            reg_file[27842] <= 8'h00;
            reg_file[27843] <= 8'h00;
            reg_file[27844] <= 8'h00;
            reg_file[27845] <= 8'h00;
            reg_file[27846] <= 8'h00;
            reg_file[27847] <= 8'h00;
            reg_file[27848] <= 8'h00;
            reg_file[27849] <= 8'h00;
            reg_file[27850] <= 8'h00;
            reg_file[27851] <= 8'h00;
            reg_file[27852] <= 8'h00;
            reg_file[27853] <= 8'h00;
            reg_file[27854] <= 8'h00;
            reg_file[27855] <= 8'h00;
            reg_file[27856] <= 8'h00;
            reg_file[27857] <= 8'h00;
            reg_file[27858] <= 8'h00;
            reg_file[27859] <= 8'h00;
            reg_file[27860] <= 8'h00;
            reg_file[27861] <= 8'h00;
            reg_file[27862] <= 8'h00;
            reg_file[27863] <= 8'h00;
            reg_file[27864] <= 8'h00;
            reg_file[27865] <= 8'h00;
            reg_file[27866] <= 8'h00;
            reg_file[27867] <= 8'h00;
            reg_file[27868] <= 8'h00;
            reg_file[27869] <= 8'h00;
            reg_file[27870] <= 8'h00;
            reg_file[27871] <= 8'h00;
            reg_file[27872] <= 8'h00;
            reg_file[27873] <= 8'h00;
            reg_file[27874] <= 8'h00;
            reg_file[27875] <= 8'h00;
            reg_file[27876] <= 8'h00;
            reg_file[27877] <= 8'h00;
            reg_file[27878] <= 8'h00;
            reg_file[27879] <= 8'h00;
            reg_file[27880] <= 8'h00;
            reg_file[27881] <= 8'h00;
            reg_file[27882] <= 8'h00;
            reg_file[27883] <= 8'h00;
            reg_file[27884] <= 8'h00;
            reg_file[27885] <= 8'h00;
            reg_file[27886] <= 8'h00;
            reg_file[27887] <= 8'h00;
            reg_file[27888] <= 8'h00;
            reg_file[27889] <= 8'h00;
            reg_file[27890] <= 8'h00;
            reg_file[27891] <= 8'h00;
            reg_file[27892] <= 8'h00;
            reg_file[27893] <= 8'h00;
            reg_file[27894] <= 8'h00;
            reg_file[27895] <= 8'h00;
            reg_file[27896] <= 8'h00;
            reg_file[27897] <= 8'h00;
            reg_file[27898] <= 8'h00;
            reg_file[27899] <= 8'h00;
            reg_file[27900] <= 8'h00;
            reg_file[27901] <= 8'h00;
            reg_file[27902] <= 8'h00;
            reg_file[27903] <= 8'h00;
            reg_file[27904] <= 8'h00;
            reg_file[27905] <= 8'h00;
            reg_file[27906] <= 8'h00;
            reg_file[27907] <= 8'h00;
            reg_file[27908] <= 8'h00;
            reg_file[27909] <= 8'h00;
            reg_file[27910] <= 8'h00;
            reg_file[27911] <= 8'h00;
            reg_file[27912] <= 8'h00;
            reg_file[27913] <= 8'h00;
            reg_file[27914] <= 8'h00;
            reg_file[27915] <= 8'h00;
            reg_file[27916] <= 8'h00;
            reg_file[27917] <= 8'h00;
            reg_file[27918] <= 8'h00;
            reg_file[27919] <= 8'h00;
            reg_file[27920] <= 8'h00;
            reg_file[27921] <= 8'h00;
            reg_file[27922] <= 8'h00;
            reg_file[27923] <= 8'h00;
            reg_file[27924] <= 8'h00;
            reg_file[27925] <= 8'h00;
            reg_file[27926] <= 8'h00;
            reg_file[27927] <= 8'h00;
            reg_file[27928] <= 8'h00;
            reg_file[27929] <= 8'h00;
            reg_file[27930] <= 8'h00;
            reg_file[27931] <= 8'h00;
            reg_file[27932] <= 8'h00;
            reg_file[27933] <= 8'h00;
            reg_file[27934] <= 8'h00;
            reg_file[27935] <= 8'h00;
            reg_file[27936] <= 8'h00;
            reg_file[27937] <= 8'h00;
            reg_file[27938] <= 8'h00;
            reg_file[27939] <= 8'h00;
            reg_file[27940] <= 8'h00;
            reg_file[27941] <= 8'h00;
            reg_file[27942] <= 8'h00;
            reg_file[27943] <= 8'h00;
            reg_file[27944] <= 8'h00;
            reg_file[27945] <= 8'h00;
            reg_file[27946] <= 8'h00;
            reg_file[27947] <= 8'h00;
            reg_file[27948] <= 8'h00;
            reg_file[27949] <= 8'h00;
            reg_file[27950] <= 8'h00;
            reg_file[27951] <= 8'h00;
            reg_file[27952] <= 8'h00;
            reg_file[27953] <= 8'h00;
            reg_file[27954] <= 8'h00;
            reg_file[27955] <= 8'h00;
            reg_file[27956] <= 8'h00;
            reg_file[27957] <= 8'h00;
            reg_file[27958] <= 8'h00;
            reg_file[27959] <= 8'h00;
            reg_file[27960] <= 8'h00;
            reg_file[27961] <= 8'h00;
            reg_file[27962] <= 8'h00;
            reg_file[27963] <= 8'h00;
            reg_file[27964] <= 8'h00;
            reg_file[27965] <= 8'h00;
            reg_file[27966] <= 8'h00;
            reg_file[27967] <= 8'h00;
            reg_file[27968] <= 8'h00;
            reg_file[27969] <= 8'h00;
            reg_file[27970] <= 8'h00;
            reg_file[27971] <= 8'h00;
            reg_file[27972] <= 8'h00;
            reg_file[27973] <= 8'h00;
            reg_file[27974] <= 8'h00;
            reg_file[27975] <= 8'h00;
            reg_file[27976] <= 8'h00;
            reg_file[27977] <= 8'h00;
            reg_file[27978] <= 8'h00;
            reg_file[27979] <= 8'h00;
            reg_file[27980] <= 8'h00;
            reg_file[27981] <= 8'h00;
            reg_file[27982] <= 8'h00;
            reg_file[27983] <= 8'h00;
            reg_file[27984] <= 8'h00;
            reg_file[27985] <= 8'h00;
            reg_file[27986] <= 8'h00;
            reg_file[27987] <= 8'h00;
            reg_file[27988] <= 8'h00;
            reg_file[27989] <= 8'h00;
            reg_file[27990] <= 8'h00;
            reg_file[27991] <= 8'h00;
            reg_file[27992] <= 8'h00;
            reg_file[27993] <= 8'h00;
            reg_file[27994] <= 8'h00;
            reg_file[27995] <= 8'h00;
            reg_file[27996] <= 8'h00;
            reg_file[27997] <= 8'h00;
            reg_file[27998] <= 8'h00;
            reg_file[27999] <= 8'h00;
            reg_file[28000] <= 8'h00;
            reg_file[28001] <= 8'h00;
            reg_file[28002] <= 8'h00;
            reg_file[28003] <= 8'h00;
            reg_file[28004] <= 8'h00;
            reg_file[28005] <= 8'h00;
            reg_file[28006] <= 8'h00;
            reg_file[28007] <= 8'h00;
            reg_file[28008] <= 8'h00;
            reg_file[28009] <= 8'h00;
            reg_file[28010] <= 8'h00;
            reg_file[28011] <= 8'h00;
            reg_file[28012] <= 8'h00;
            reg_file[28013] <= 8'h00;
            reg_file[28014] <= 8'h00;
            reg_file[28015] <= 8'h00;
            reg_file[28016] <= 8'h00;
            reg_file[28017] <= 8'h00;
            reg_file[28018] <= 8'h00;
            reg_file[28019] <= 8'h00;
            reg_file[28020] <= 8'h00;
            reg_file[28021] <= 8'h00;
            reg_file[28022] <= 8'h00;
            reg_file[28023] <= 8'h00;
            reg_file[28024] <= 8'h00;
            reg_file[28025] <= 8'h00;
            reg_file[28026] <= 8'h00;
            reg_file[28027] <= 8'h00;
            reg_file[28028] <= 8'h00;
            reg_file[28029] <= 8'h00;
            reg_file[28030] <= 8'h00;
            reg_file[28031] <= 8'h00;
            reg_file[28032] <= 8'h00;
            reg_file[28033] <= 8'h00;
            reg_file[28034] <= 8'h00;
            reg_file[28035] <= 8'h00;
            reg_file[28036] <= 8'h00;
            reg_file[28037] <= 8'h00;
            reg_file[28038] <= 8'h00;
            reg_file[28039] <= 8'h00;
            reg_file[28040] <= 8'h00;
            reg_file[28041] <= 8'h00;
            reg_file[28042] <= 8'h00;
            reg_file[28043] <= 8'h00;
            reg_file[28044] <= 8'h00;
            reg_file[28045] <= 8'h00;
            reg_file[28046] <= 8'h00;
            reg_file[28047] <= 8'h00;
            reg_file[28048] <= 8'h00;
            reg_file[28049] <= 8'h00;
            reg_file[28050] <= 8'h00;
            reg_file[28051] <= 8'h00;
            reg_file[28052] <= 8'h00;
            reg_file[28053] <= 8'h00;
            reg_file[28054] <= 8'h00;
            reg_file[28055] <= 8'h00;
            reg_file[28056] <= 8'h00;
            reg_file[28057] <= 8'h00;
            reg_file[28058] <= 8'h00;
            reg_file[28059] <= 8'h00;
            reg_file[28060] <= 8'h00;
            reg_file[28061] <= 8'h00;
            reg_file[28062] <= 8'h00;
            reg_file[28063] <= 8'h00;
            reg_file[28064] <= 8'h00;
            reg_file[28065] <= 8'h00;
            reg_file[28066] <= 8'h00;
            reg_file[28067] <= 8'h00;
            reg_file[28068] <= 8'h00;
            reg_file[28069] <= 8'h00;
            reg_file[28070] <= 8'h00;
            reg_file[28071] <= 8'h00;
            reg_file[28072] <= 8'h00;
            reg_file[28073] <= 8'h00;
            reg_file[28074] <= 8'h00;
            reg_file[28075] <= 8'h00;
            reg_file[28076] <= 8'h00;
            reg_file[28077] <= 8'h00;
            reg_file[28078] <= 8'h00;
            reg_file[28079] <= 8'h00;
            reg_file[28080] <= 8'h00;
            reg_file[28081] <= 8'h00;
            reg_file[28082] <= 8'h00;
            reg_file[28083] <= 8'h00;
            reg_file[28084] <= 8'h00;
            reg_file[28085] <= 8'h00;
            reg_file[28086] <= 8'h00;
            reg_file[28087] <= 8'h00;
            reg_file[28088] <= 8'h00;
            reg_file[28089] <= 8'h00;
            reg_file[28090] <= 8'h00;
            reg_file[28091] <= 8'h00;
            reg_file[28092] <= 8'h00;
            reg_file[28093] <= 8'h00;
            reg_file[28094] <= 8'h00;
            reg_file[28095] <= 8'h00;
            reg_file[28096] <= 8'h00;
            reg_file[28097] <= 8'h00;
            reg_file[28098] <= 8'h00;
            reg_file[28099] <= 8'h00;
            reg_file[28100] <= 8'h00;
            reg_file[28101] <= 8'h00;
            reg_file[28102] <= 8'h00;
            reg_file[28103] <= 8'h00;
            reg_file[28104] <= 8'h00;
            reg_file[28105] <= 8'h00;
            reg_file[28106] <= 8'h00;
            reg_file[28107] <= 8'h00;
            reg_file[28108] <= 8'h00;
            reg_file[28109] <= 8'h00;
            reg_file[28110] <= 8'h00;
            reg_file[28111] <= 8'h00;
            reg_file[28112] <= 8'h00;
            reg_file[28113] <= 8'h00;
            reg_file[28114] <= 8'h00;
            reg_file[28115] <= 8'h00;
            reg_file[28116] <= 8'h00;
            reg_file[28117] <= 8'h00;
            reg_file[28118] <= 8'h00;
            reg_file[28119] <= 8'h00;
            reg_file[28120] <= 8'h00;
            reg_file[28121] <= 8'h00;
            reg_file[28122] <= 8'h00;
            reg_file[28123] <= 8'h00;
            reg_file[28124] <= 8'h00;
            reg_file[28125] <= 8'h00;
            reg_file[28126] <= 8'h00;
            reg_file[28127] <= 8'h00;
            reg_file[28128] <= 8'h00;
            reg_file[28129] <= 8'h00;
            reg_file[28130] <= 8'h00;
            reg_file[28131] <= 8'h00;
            reg_file[28132] <= 8'h00;
            reg_file[28133] <= 8'h00;
            reg_file[28134] <= 8'h00;
            reg_file[28135] <= 8'h00;
            reg_file[28136] <= 8'h00;
            reg_file[28137] <= 8'h00;
            reg_file[28138] <= 8'h00;
            reg_file[28139] <= 8'h00;
            reg_file[28140] <= 8'h00;
            reg_file[28141] <= 8'h00;
            reg_file[28142] <= 8'h00;
            reg_file[28143] <= 8'h00;
            reg_file[28144] <= 8'h00;
            reg_file[28145] <= 8'h00;
            reg_file[28146] <= 8'h00;
            reg_file[28147] <= 8'h00;
            reg_file[28148] <= 8'h00;
            reg_file[28149] <= 8'h00;
            reg_file[28150] <= 8'h00;
            reg_file[28151] <= 8'h00;
            reg_file[28152] <= 8'h00;
            reg_file[28153] <= 8'h00;
            reg_file[28154] <= 8'h00;
            reg_file[28155] <= 8'h00;
            reg_file[28156] <= 8'h00;
            reg_file[28157] <= 8'h00;
            reg_file[28158] <= 8'h00;
            reg_file[28159] <= 8'h00;
            reg_file[28160] <= 8'h00;
            reg_file[28161] <= 8'h00;
            reg_file[28162] <= 8'h00;
            reg_file[28163] <= 8'h00;
            reg_file[28164] <= 8'h00;
            reg_file[28165] <= 8'h00;
            reg_file[28166] <= 8'h00;
            reg_file[28167] <= 8'h00;
            reg_file[28168] <= 8'h00;
            reg_file[28169] <= 8'h00;
            reg_file[28170] <= 8'h00;
            reg_file[28171] <= 8'h00;
            reg_file[28172] <= 8'h00;
            reg_file[28173] <= 8'h00;
            reg_file[28174] <= 8'h00;
            reg_file[28175] <= 8'h00;
            reg_file[28176] <= 8'h00;
            reg_file[28177] <= 8'h00;
            reg_file[28178] <= 8'h00;
            reg_file[28179] <= 8'h00;
            reg_file[28180] <= 8'h00;
            reg_file[28181] <= 8'h00;
            reg_file[28182] <= 8'h00;
            reg_file[28183] <= 8'h00;
            reg_file[28184] <= 8'h00;
            reg_file[28185] <= 8'h00;
            reg_file[28186] <= 8'h00;
            reg_file[28187] <= 8'h00;
            reg_file[28188] <= 8'h00;
            reg_file[28189] <= 8'h00;
            reg_file[28190] <= 8'h00;
            reg_file[28191] <= 8'h00;
            reg_file[28192] <= 8'h00;
            reg_file[28193] <= 8'h00;
            reg_file[28194] <= 8'h00;
            reg_file[28195] <= 8'h00;
            reg_file[28196] <= 8'h00;
            reg_file[28197] <= 8'h00;
            reg_file[28198] <= 8'h00;
            reg_file[28199] <= 8'h00;
            reg_file[28200] <= 8'h00;
            reg_file[28201] <= 8'h00;
            reg_file[28202] <= 8'h00;
            reg_file[28203] <= 8'h00;
            reg_file[28204] <= 8'h00;
            reg_file[28205] <= 8'h00;
            reg_file[28206] <= 8'h00;
            reg_file[28207] <= 8'h00;
            reg_file[28208] <= 8'h00;
            reg_file[28209] <= 8'h00;
            reg_file[28210] <= 8'h00;
            reg_file[28211] <= 8'h00;
            reg_file[28212] <= 8'h00;
            reg_file[28213] <= 8'h00;
            reg_file[28214] <= 8'h00;
            reg_file[28215] <= 8'h00;
            reg_file[28216] <= 8'h00;
            reg_file[28217] <= 8'h00;
            reg_file[28218] <= 8'h00;
            reg_file[28219] <= 8'h00;
            reg_file[28220] <= 8'h00;
            reg_file[28221] <= 8'h00;
            reg_file[28222] <= 8'h00;
            reg_file[28223] <= 8'h00;
            reg_file[28224] <= 8'h00;
            reg_file[28225] <= 8'h00;
            reg_file[28226] <= 8'h00;
            reg_file[28227] <= 8'h00;
            reg_file[28228] <= 8'h00;
            reg_file[28229] <= 8'h00;
            reg_file[28230] <= 8'h00;
            reg_file[28231] <= 8'h00;
            reg_file[28232] <= 8'h00;
            reg_file[28233] <= 8'h00;
            reg_file[28234] <= 8'h00;
            reg_file[28235] <= 8'h00;
            reg_file[28236] <= 8'h00;
            reg_file[28237] <= 8'h00;
            reg_file[28238] <= 8'h00;
            reg_file[28239] <= 8'h00;
            reg_file[28240] <= 8'h00;
            reg_file[28241] <= 8'h00;
            reg_file[28242] <= 8'h00;
            reg_file[28243] <= 8'h00;
            reg_file[28244] <= 8'h00;
            reg_file[28245] <= 8'h00;
            reg_file[28246] <= 8'h00;
            reg_file[28247] <= 8'h00;
            reg_file[28248] <= 8'h00;
            reg_file[28249] <= 8'h00;
            reg_file[28250] <= 8'h00;
            reg_file[28251] <= 8'h00;
            reg_file[28252] <= 8'h00;
            reg_file[28253] <= 8'h00;
            reg_file[28254] <= 8'h00;
            reg_file[28255] <= 8'h00;
            reg_file[28256] <= 8'h00;
            reg_file[28257] <= 8'h00;
            reg_file[28258] <= 8'h00;
            reg_file[28259] <= 8'h00;
            reg_file[28260] <= 8'h00;
            reg_file[28261] <= 8'h00;
            reg_file[28262] <= 8'h00;
            reg_file[28263] <= 8'h00;
            reg_file[28264] <= 8'h00;
            reg_file[28265] <= 8'h00;
            reg_file[28266] <= 8'h00;
            reg_file[28267] <= 8'h00;
            reg_file[28268] <= 8'h00;
            reg_file[28269] <= 8'h00;
            reg_file[28270] <= 8'h00;
            reg_file[28271] <= 8'h00;
            reg_file[28272] <= 8'h00;
            reg_file[28273] <= 8'h00;
            reg_file[28274] <= 8'h00;
            reg_file[28275] <= 8'h00;
            reg_file[28276] <= 8'h00;
            reg_file[28277] <= 8'h00;
            reg_file[28278] <= 8'h00;
            reg_file[28279] <= 8'h00;
            reg_file[28280] <= 8'h00;
            reg_file[28281] <= 8'h00;
            reg_file[28282] <= 8'h00;
            reg_file[28283] <= 8'h00;
            reg_file[28284] <= 8'h00;
            reg_file[28285] <= 8'h00;
            reg_file[28286] <= 8'h00;
            reg_file[28287] <= 8'h00;
            reg_file[28288] <= 8'h00;
            reg_file[28289] <= 8'h00;
            reg_file[28290] <= 8'h00;
            reg_file[28291] <= 8'h00;
            reg_file[28292] <= 8'h00;
            reg_file[28293] <= 8'h00;
            reg_file[28294] <= 8'h00;
            reg_file[28295] <= 8'h00;
            reg_file[28296] <= 8'h00;
            reg_file[28297] <= 8'h00;
            reg_file[28298] <= 8'h00;
            reg_file[28299] <= 8'h00;
            reg_file[28300] <= 8'h00;
            reg_file[28301] <= 8'h00;
            reg_file[28302] <= 8'h00;
            reg_file[28303] <= 8'h00;
            reg_file[28304] <= 8'h00;
            reg_file[28305] <= 8'h00;
            reg_file[28306] <= 8'h00;
            reg_file[28307] <= 8'h00;
            reg_file[28308] <= 8'h00;
            reg_file[28309] <= 8'h00;
            reg_file[28310] <= 8'h00;
            reg_file[28311] <= 8'h00;
            reg_file[28312] <= 8'h00;
            reg_file[28313] <= 8'h00;
            reg_file[28314] <= 8'h00;
            reg_file[28315] <= 8'h00;
            reg_file[28316] <= 8'h00;
            reg_file[28317] <= 8'h00;
            reg_file[28318] <= 8'h00;
            reg_file[28319] <= 8'h00;
            reg_file[28320] <= 8'h00;
            reg_file[28321] <= 8'h00;
            reg_file[28322] <= 8'h00;
            reg_file[28323] <= 8'h00;
            reg_file[28324] <= 8'h00;
            reg_file[28325] <= 8'h00;
            reg_file[28326] <= 8'h00;
            reg_file[28327] <= 8'h00;
            reg_file[28328] <= 8'h00;
            reg_file[28329] <= 8'h00;
            reg_file[28330] <= 8'h00;
            reg_file[28331] <= 8'h00;
            reg_file[28332] <= 8'h00;
            reg_file[28333] <= 8'h00;
            reg_file[28334] <= 8'h00;
            reg_file[28335] <= 8'h00;
            reg_file[28336] <= 8'h00;
            reg_file[28337] <= 8'h00;
            reg_file[28338] <= 8'h00;
            reg_file[28339] <= 8'h00;
            reg_file[28340] <= 8'h00;
            reg_file[28341] <= 8'h00;
            reg_file[28342] <= 8'h00;
            reg_file[28343] <= 8'h00;
            reg_file[28344] <= 8'h00;
            reg_file[28345] <= 8'h00;
            reg_file[28346] <= 8'h00;
            reg_file[28347] <= 8'h00;
            reg_file[28348] <= 8'h00;
            reg_file[28349] <= 8'h00;
            reg_file[28350] <= 8'h00;
            reg_file[28351] <= 8'h00;
            reg_file[28352] <= 8'h00;
            reg_file[28353] <= 8'h00;
            reg_file[28354] <= 8'h00;
            reg_file[28355] <= 8'h00;
            reg_file[28356] <= 8'h00;
            reg_file[28357] <= 8'h00;
            reg_file[28358] <= 8'h00;
            reg_file[28359] <= 8'h00;
            reg_file[28360] <= 8'h00;
            reg_file[28361] <= 8'h00;
            reg_file[28362] <= 8'h00;
            reg_file[28363] <= 8'h00;
            reg_file[28364] <= 8'h00;
            reg_file[28365] <= 8'h00;
            reg_file[28366] <= 8'h00;
            reg_file[28367] <= 8'h00;
            reg_file[28368] <= 8'h00;
            reg_file[28369] <= 8'h00;
            reg_file[28370] <= 8'h00;
            reg_file[28371] <= 8'h00;
            reg_file[28372] <= 8'h00;
            reg_file[28373] <= 8'h00;
            reg_file[28374] <= 8'h00;
            reg_file[28375] <= 8'h00;
            reg_file[28376] <= 8'h00;
            reg_file[28377] <= 8'h00;
            reg_file[28378] <= 8'h00;
            reg_file[28379] <= 8'h00;
            reg_file[28380] <= 8'h00;
            reg_file[28381] <= 8'h00;
            reg_file[28382] <= 8'h00;
            reg_file[28383] <= 8'h00;
            reg_file[28384] <= 8'h00;
            reg_file[28385] <= 8'h00;
            reg_file[28386] <= 8'h00;
            reg_file[28387] <= 8'h00;
            reg_file[28388] <= 8'h00;
            reg_file[28389] <= 8'h00;
            reg_file[28390] <= 8'h00;
            reg_file[28391] <= 8'h00;
            reg_file[28392] <= 8'h00;
            reg_file[28393] <= 8'h00;
            reg_file[28394] <= 8'h00;
            reg_file[28395] <= 8'h00;
            reg_file[28396] <= 8'h00;
            reg_file[28397] <= 8'h00;
            reg_file[28398] <= 8'h00;
            reg_file[28399] <= 8'h00;
            reg_file[28400] <= 8'h00;
            reg_file[28401] <= 8'h00;
            reg_file[28402] <= 8'h00;
            reg_file[28403] <= 8'h00;
            reg_file[28404] <= 8'h00;
            reg_file[28405] <= 8'h00;
            reg_file[28406] <= 8'h00;
            reg_file[28407] <= 8'h00;
            reg_file[28408] <= 8'h00;
            reg_file[28409] <= 8'h00;
            reg_file[28410] <= 8'h00;
            reg_file[28411] <= 8'h00;
            reg_file[28412] <= 8'h00;
            reg_file[28413] <= 8'h00;
            reg_file[28414] <= 8'h00;
            reg_file[28415] <= 8'h00;
            reg_file[28416] <= 8'h00;
            reg_file[28417] <= 8'h00;
            reg_file[28418] <= 8'h00;
            reg_file[28419] <= 8'h00;
            reg_file[28420] <= 8'h00;
            reg_file[28421] <= 8'h00;
            reg_file[28422] <= 8'h00;
            reg_file[28423] <= 8'h00;
            reg_file[28424] <= 8'h00;
            reg_file[28425] <= 8'h00;
            reg_file[28426] <= 8'h00;
            reg_file[28427] <= 8'h00;
            reg_file[28428] <= 8'h00;
            reg_file[28429] <= 8'h00;
            reg_file[28430] <= 8'h00;
            reg_file[28431] <= 8'h00;
            reg_file[28432] <= 8'h00;
            reg_file[28433] <= 8'h00;
            reg_file[28434] <= 8'h00;
            reg_file[28435] <= 8'h00;
            reg_file[28436] <= 8'h00;
            reg_file[28437] <= 8'h00;
            reg_file[28438] <= 8'h00;
            reg_file[28439] <= 8'h00;
            reg_file[28440] <= 8'h00;
            reg_file[28441] <= 8'h00;
            reg_file[28442] <= 8'h00;
            reg_file[28443] <= 8'h00;
            reg_file[28444] <= 8'h00;
            reg_file[28445] <= 8'h00;
            reg_file[28446] <= 8'h00;
            reg_file[28447] <= 8'h00;
            reg_file[28448] <= 8'h00;
            reg_file[28449] <= 8'h00;
            reg_file[28450] <= 8'h00;
            reg_file[28451] <= 8'h00;
            reg_file[28452] <= 8'h00;
            reg_file[28453] <= 8'h00;
            reg_file[28454] <= 8'h00;
            reg_file[28455] <= 8'h00;
            reg_file[28456] <= 8'h00;
            reg_file[28457] <= 8'h00;
            reg_file[28458] <= 8'h00;
            reg_file[28459] <= 8'h00;
            reg_file[28460] <= 8'h00;
            reg_file[28461] <= 8'h00;
            reg_file[28462] <= 8'h00;
            reg_file[28463] <= 8'h00;
            reg_file[28464] <= 8'h00;
            reg_file[28465] <= 8'h00;
            reg_file[28466] <= 8'h00;
            reg_file[28467] <= 8'h00;
            reg_file[28468] <= 8'h00;
            reg_file[28469] <= 8'h00;
            reg_file[28470] <= 8'h00;
            reg_file[28471] <= 8'h00;
            reg_file[28472] <= 8'h00;
            reg_file[28473] <= 8'h00;
            reg_file[28474] <= 8'h00;
            reg_file[28475] <= 8'h00;
            reg_file[28476] <= 8'h00;
            reg_file[28477] <= 8'h00;
            reg_file[28478] <= 8'h00;
            reg_file[28479] <= 8'h00;
            reg_file[28480] <= 8'h00;
            reg_file[28481] <= 8'h00;
            reg_file[28482] <= 8'h00;
            reg_file[28483] <= 8'h00;
            reg_file[28484] <= 8'h00;
            reg_file[28485] <= 8'h00;
            reg_file[28486] <= 8'h00;
            reg_file[28487] <= 8'h00;
            reg_file[28488] <= 8'h00;
            reg_file[28489] <= 8'h00;
            reg_file[28490] <= 8'h00;
            reg_file[28491] <= 8'h00;
            reg_file[28492] <= 8'h00;
            reg_file[28493] <= 8'h00;
            reg_file[28494] <= 8'h00;
            reg_file[28495] <= 8'h00;
            reg_file[28496] <= 8'h00;
            reg_file[28497] <= 8'h00;
            reg_file[28498] <= 8'h00;
            reg_file[28499] <= 8'h00;
            reg_file[28500] <= 8'h00;
            reg_file[28501] <= 8'h00;
            reg_file[28502] <= 8'h00;
            reg_file[28503] <= 8'h00;
            reg_file[28504] <= 8'h00;
            reg_file[28505] <= 8'h00;
            reg_file[28506] <= 8'h00;
            reg_file[28507] <= 8'h00;
            reg_file[28508] <= 8'h00;
            reg_file[28509] <= 8'h00;
            reg_file[28510] <= 8'h00;
            reg_file[28511] <= 8'h00;
            reg_file[28512] <= 8'h00;
            reg_file[28513] <= 8'h00;
            reg_file[28514] <= 8'h00;
            reg_file[28515] <= 8'h00;
            reg_file[28516] <= 8'h00;
            reg_file[28517] <= 8'h00;
            reg_file[28518] <= 8'h00;
            reg_file[28519] <= 8'h00;
            reg_file[28520] <= 8'h00;
            reg_file[28521] <= 8'h00;
            reg_file[28522] <= 8'h00;
            reg_file[28523] <= 8'h00;
            reg_file[28524] <= 8'h00;
            reg_file[28525] <= 8'h00;
            reg_file[28526] <= 8'h00;
            reg_file[28527] <= 8'h00;
            reg_file[28528] <= 8'h00;
            reg_file[28529] <= 8'h00;
            reg_file[28530] <= 8'h00;
            reg_file[28531] <= 8'h00;
            reg_file[28532] <= 8'h00;
            reg_file[28533] <= 8'h00;
            reg_file[28534] <= 8'h00;
            reg_file[28535] <= 8'h00;
            reg_file[28536] <= 8'h00;
            reg_file[28537] <= 8'h00;
            reg_file[28538] <= 8'h00;
            reg_file[28539] <= 8'h00;
            reg_file[28540] <= 8'h00;
            reg_file[28541] <= 8'h00;
            reg_file[28542] <= 8'h00;
            reg_file[28543] <= 8'h00;
            reg_file[28544] <= 8'h00;
            reg_file[28545] <= 8'h00;
            reg_file[28546] <= 8'h00;
            reg_file[28547] <= 8'h00;
            reg_file[28548] <= 8'h00;
            reg_file[28549] <= 8'h00;
            reg_file[28550] <= 8'h00;
            reg_file[28551] <= 8'h00;
            reg_file[28552] <= 8'h00;
            reg_file[28553] <= 8'h00;
            reg_file[28554] <= 8'h00;
            reg_file[28555] <= 8'h00;
            reg_file[28556] <= 8'h00;
            reg_file[28557] <= 8'h00;
            reg_file[28558] <= 8'h00;
            reg_file[28559] <= 8'h00;
            reg_file[28560] <= 8'h00;
            reg_file[28561] <= 8'h00;
            reg_file[28562] <= 8'h00;
            reg_file[28563] <= 8'h00;
            reg_file[28564] <= 8'h00;
            reg_file[28565] <= 8'h00;
            reg_file[28566] <= 8'h00;
            reg_file[28567] <= 8'h00;
            reg_file[28568] <= 8'h00;
            reg_file[28569] <= 8'h00;
            reg_file[28570] <= 8'h00;
            reg_file[28571] <= 8'h00;
            reg_file[28572] <= 8'h00;
            reg_file[28573] <= 8'h00;
            reg_file[28574] <= 8'h00;
            reg_file[28575] <= 8'h00;
            reg_file[28576] <= 8'h00;
            reg_file[28577] <= 8'h00;
            reg_file[28578] <= 8'h00;
            reg_file[28579] <= 8'h00;
            reg_file[28580] <= 8'h00;
            reg_file[28581] <= 8'h00;
            reg_file[28582] <= 8'h00;
            reg_file[28583] <= 8'h00;
            reg_file[28584] <= 8'h00;
            reg_file[28585] <= 8'h00;
            reg_file[28586] <= 8'h00;
            reg_file[28587] <= 8'h00;
            reg_file[28588] <= 8'h00;
            reg_file[28589] <= 8'h00;
            reg_file[28590] <= 8'h00;
            reg_file[28591] <= 8'h00;
            reg_file[28592] <= 8'h00;
            reg_file[28593] <= 8'h00;
            reg_file[28594] <= 8'h00;
            reg_file[28595] <= 8'h00;
            reg_file[28596] <= 8'h00;
            reg_file[28597] <= 8'h00;
            reg_file[28598] <= 8'h00;
            reg_file[28599] <= 8'h00;
            reg_file[28600] <= 8'h00;
            reg_file[28601] <= 8'h00;
            reg_file[28602] <= 8'h00;
            reg_file[28603] <= 8'h00;
            reg_file[28604] <= 8'h00;
            reg_file[28605] <= 8'h00;
            reg_file[28606] <= 8'h00;
            reg_file[28607] <= 8'h00;
            reg_file[28608] <= 8'h00;
            reg_file[28609] <= 8'h00;
            reg_file[28610] <= 8'h00;
            reg_file[28611] <= 8'h00;
            reg_file[28612] <= 8'h00;
            reg_file[28613] <= 8'h00;
            reg_file[28614] <= 8'h00;
            reg_file[28615] <= 8'h00;
            reg_file[28616] <= 8'h00;
            reg_file[28617] <= 8'h00;
            reg_file[28618] <= 8'h00;
            reg_file[28619] <= 8'h00;
            reg_file[28620] <= 8'h00;
            reg_file[28621] <= 8'h00;
            reg_file[28622] <= 8'h00;
            reg_file[28623] <= 8'h00;
            reg_file[28624] <= 8'h00;
            reg_file[28625] <= 8'h00;
            reg_file[28626] <= 8'h00;
            reg_file[28627] <= 8'h00;
            reg_file[28628] <= 8'h00;
            reg_file[28629] <= 8'h00;
            reg_file[28630] <= 8'h00;
            reg_file[28631] <= 8'h00;
            reg_file[28632] <= 8'h00;
            reg_file[28633] <= 8'h00;
            reg_file[28634] <= 8'h00;
            reg_file[28635] <= 8'h00;
            reg_file[28636] <= 8'h00;
            reg_file[28637] <= 8'h00;
            reg_file[28638] <= 8'h00;
            reg_file[28639] <= 8'h00;
            reg_file[28640] <= 8'h00;
            reg_file[28641] <= 8'h00;
            reg_file[28642] <= 8'h00;
            reg_file[28643] <= 8'h00;
            reg_file[28644] <= 8'h00;
            reg_file[28645] <= 8'h00;
            reg_file[28646] <= 8'h00;
            reg_file[28647] <= 8'h00;
            reg_file[28648] <= 8'h00;
            reg_file[28649] <= 8'h00;
            reg_file[28650] <= 8'h00;
            reg_file[28651] <= 8'h00;
            reg_file[28652] <= 8'h00;
            reg_file[28653] <= 8'h00;
            reg_file[28654] <= 8'h00;
            reg_file[28655] <= 8'h00;
            reg_file[28656] <= 8'h00;
            reg_file[28657] <= 8'h00;
            reg_file[28658] <= 8'h00;
            reg_file[28659] <= 8'h00;
            reg_file[28660] <= 8'h00;
            reg_file[28661] <= 8'h00;
            reg_file[28662] <= 8'h00;
            reg_file[28663] <= 8'h00;
            reg_file[28664] <= 8'h00;
            reg_file[28665] <= 8'h00;
            reg_file[28666] <= 8'h00;
            reg_file[28667] <= 8'h00;
            reg_file[28668] <= 8'h00;
            reg_file[28669] <= 8'h00;
            reg_file[28670] <= 8'h00;
            reg_file[28671] <= 8'h00;
            reg_file[28672] <= 8'h00;
            reg_file[28673] <= 8'h00;
            reg_file[28674] <= 8'h00;
            reg_file[28675] <= 8'h00;
            reg_file[28676] <= 8'h00;
            reg_file[28677] <= 8'h00;
            reg_file[28678] <= 8'h00;
            reg_file[28679] <= 8'h00;
            reg_file[28680] <= 8'h00;
            reg_file[28681] <= 8'h00;
            reg_file[28682] <= 8'h00;
            reg_file[28683] <= 8'h00;
            reg_file[28684] <= 8'h00;
            reg_file[28685] <= 8'h00;
            reg_file[28686] <= 8'h00;
            reg_file[28687] <= 8'h00;
            reg_file[28688] <= 8'h00;
            reg_file[28689] <= 8'h00;
            reg_file[28690] <= 8'h00;
            reg_file[28691] <= 8'h00;
            reg_file[28692] <= 8'h00;
            reg_file[28693] <= 8'h00;
            reg_file[28694] <= 8'h00;
            reg_file[28695] <= 8'h00;
            reg_file[28696] <= 8'h00;
            reg_file[28697] <= 8'h00;
            reg_file[28698] <= 8'h00;
            reg_file[28699] <= 8'h00;
            reg_file[28700] <= 8'h00;
            reg_file[28701] <= 8'h00;
            reg_file[28702] <= 8'h00;
            reg_file[28703] <= 8'h00;
            reg_file[28704] <= 8'h00;
            reg_file[28705] <= 8'h00;
            reg_file[28706] <= 8'h00;
            reg_file[28707] <= 8'h00;
            reg_file[28708] <= 8'h00;
            reg_file[28709] <= 8'h00;
            reg_file[28710] <= 8'h00;
            reg_file[28711] <= 8'h00;
            reg_file[28712] <= 8'h00;
            reg_file[28713] <= 8'h00;
            reg_file[28714] <= 8'h00;
            reg_file[28715] <= 8'h00;
            reg_file[28716] <= 8'h00;
            reg_file[28717] <= 8'h00;
            reg_file[28718] <= 8'h00;
            reg_file[28719] <= 8'h00;
            reg_file[28720] <= 8'h00;
            reg_file[28721] <= 8'h00;
            reg_file[28722] <= 8'h00;
            reg_file[28723] <= 8'h00;
            reg_file[28724] <= 8'h00;
            reg_file[28725] <= 8'h00;
            reg_file[28726] <= 8'h00;
            reg_file[28727] <= 8'h00;
            reg_file[28728] <= 8'h00;
            reg_file[28729] <= 8'h00;
            reg_file[28730] <= 8'h00;
            reg_file[28731] <= 8'h00;
            reg_file[28732] <= 8'h00;
            reg_file[28733] <= 8'h00;
            reg_file[28734] <= 8'h00;
            reg_file[28735] <= 8'h00;
            reg_file[28736] <= 8'h00;
            reg_file[28737] <= 8'h00;
            reg_file[28738] <= 8'h00;
            reg_file[28739] <= 8'h00;
            reg_file[28740] <= 8'h00;
            reg_file[28741] <= 8'h00;
            reg_file[28742] <= 8'h00;
            reg_file[28743] <= 8'h00;
            reg_file[28744] <= 8'h00;
            reg_file[28745] <= 8'h00;
            reg_file[28746] <= 8'h00;
            reg_file[28747] <= 8'h00;
            reg_file[28748] <= 8'h00;
            reg_file[28749] <= 8'h00;
            reg_file[28750] <= 8'h00;
            reg_file[28751] <= 8'h00;
            reg_file[28752] <= 8'h00;
            reg_file[28753] <= 8'h00;
            reg_file[28754] <= 8'h00;
            reg_file[28755] <= 8'h00;
            reg_file[28756] <= 8'h00;
            reg_file[28757] <= 8'h00;
            reg_file[28758] <= 8'h00;
            reg_file[28759] <= 8'h00;
            reg_file[28760] <= 8'h00;
            reg_file[28761] <= 8'h00;
            reg_file[28762] <= 8'h00;
            reg_file[28763] <= 8'h00;
            reg_file[28764] <= 8'h00;
            reg_file[28765] <= 8'h00;
            reg_file[28766] <= 8'h00;
            reg_file[28767] <= 8'h00;
            reg_file[28768] <= 8'h00;
            reg_file[28769] <= 8'h00;
            reg_file[28770] <= 8'h00;
            reg_file[28771] <= 8'h00;
            reg_file[28772] <= 8'h00;
            reg_file[28773] <= 8'h00;
            reg_file[28774] <= 8'h00;
            reg_file[28775] <= 8'h00;
            reg_file[28776] <= 8'h00;
            reg_file[28777] <= 8'h00;
            reg_file[28778] <= 8'h00;
            reg_file[28779] <= 8'h00;
            reg_file[28780] <= 8'h00;
            reg_file[28781] <= 8'h00;
            reg_file[28782] <= 8'h00;
            reg_file[28783] <= 8'h00;
            reg_file[28784] <= 8'h00;
            reg_file[28785] <= 8'h00;
            reg_file[28786] <= 8'h00;
            reg_file[28787] <= 8'h00;
            reg_file[28788] <= 8'h00;
            reg_file[28789] <= 8'h00;
            reg_file[28790] <= 8'h00;
            reg_file[28791] <= 8'h00;
            reg_file[28792] <= 8'h00;
            reg_file[28793] <= 8'h00;
            reg_file[28794] <= 8'h00;
            reg_file[28795] <= 8'h00;
            reg_file[28796] <= 8'h00;
            reg_file[28797] <= 8'h00;
            reg_file[28798] <= 8'h00;
            reg_file[28799] <= 8'h00;
            reg_file[28800] <= 8'h00;
            reg_file[28801] <= 8'h00;
            reg_file[28802] <= 8'h00;
            reg_file[28803] <= 8'h00;
            reg_file[28804] <= 8'h00;
            reg_file[28805] <= 8'h00;
            reg_file[28806] <= 8'h00;
            reg_file[28807] <= 8'h00;
            reg_file[28808] <= 8'h00;
            reg_file[28809] <= 8'h00;
            reg_file[28810] <= 8'h00;
            reg_file[28811] <= 8'h00;
            reg_file[28812] <= 8'h00;
            reg_file[28813] <= 8'h00;
            reg_file[28814] <= 8'h00;
            reg_file[28815] <= 8'h00;
            reg_file[28816] <= 8'h00;
            reg_file[28817] <= 8'h00;
            reg_file[28818] <= 8'h00;
            reg_file[28819] <= 8'h00;
            reg_file[28820] <= 8'h00;
            reg_file[28821] <= 8'h00;
            reg_file[28822] <= 8'h00;
            reg_file[28823] <= 8'h00;
            reg_file[28824] <= 8'h00;
            reg_file[28825] <= 8'h00;
            reg_file[28826] <= 8'h00;
            reg_file[28827] <= 8'h00;
            reg_file[28828] <= 8'h00;
            reg_file[28829] <= 8'h00;
            reg_file[28830] <= 8'h00;
            reg_file[28831] <= 8'h00;
            reg_file[28832] <= 8'h00;
            reg_file[28833] <= 8'h00;
            reg_file[28834] <= 8'h00;
            reg_file[28835] <= 8'h00;
            reg_file[28836] <= 8'h00;
            reg_file[28837] <= 8'h00;
            reg_file[28838] <= 8'h00;
            reg_file[28839] <= 8'h00;
            reg_file[28840] <= 8'h00;
            reg_file[28841] <= 8'h00;
            reg_file[28842] <= 8'h00;
            reg_file[28843] <= 8'h00;
            reg_file[28844] <= 8'h00;
            reg_file[28845] <= 8'h00;
            reg_file[28846] <= 8'h00;
            reg_file[28847] <= 8'h00;
            reg_file[28848] <= 8'h00;
            reg_file[28849] <= 8'h00;
            reg_file[28850] <= 8'h00;
            reg_file[28851] <= 8'h00;
            reg_file[28852] <= 8'h00;
            reg_file[28853] <= 8'h00;
            reg_file[28854] <= 8'h00;
            reg_file[28855] <= 8'h00;
            reg_file[28856] <= 8'h00;
            reg_file[28857] <= 8'h00;
            reg_file[28858] <= 8'h00;
            reg_file[28859] <= 8'h00;
            reg_file[28860] <= 8'h00;
            reg_file[28861] <= 8'h00;
            reg_file[28862] <= 8'h00;
            reg_file[28863] <= 8'h00;
            reg_file[28864] <= 8'h00;
            reg_file[28865] <= 8'h00;
            reg_file[28866] <= 8'h00;
            reg_file[28867] <= 8'h00;
            reg_file[28868] <= 8'h00;
            reg_file[28869] <= 8'h00;
            reg_file[28870] <= 8'h00;
            reg_file[28871] <= 8'h00;
            reg_file[28872] <= 8'h00;
            reg_file[28873] <= 8'h00;
            reg_file[28874] <= 8'h00;
            reg_file[28875] <= 8'h00;
            reg_file[28876] <= 8'h00;
            reg_file[28877] <= 8'h00;
            reg_file[28878] <= 8'h00;
            reg_file[28879] <= 8'h00;
            reg_file[28880] <= 8'h00;
            reg_file[28881] <= 8'h00;
            reg_file[28882] <= 8'h00;
            reg_file[28883] <= 8'h00;
            reg_file[28884] <= 8'h00;
            reg_file[28885] <= 8'h00;
            reg_file[28886] <= 8'h00;
            reg_file[28887] <= 8'h00;
            reg_file[28888] <= 8'h00;
            reg_file[28889] <= 8'h00;
            reg_file[28890] <= 8'h00;
            reg_file[28891] <= 8'h00;
            reg_file[28892] <= 8'h00;
            reg_file[28893] <= 8'h00;
            reg_file[28894] <= 8'h00;
            reg_file[28895] <= 8'h00;
            reg_file[28896] <= 8'h00;
            reg_file[28897] <= 8'h00;
            reg_file[28898] <= 8'h00;
            reg_file[28899] <= 8'h00;
            reg_file[28900] <= 8'h00;
            reg_file[28901] <= 8'h00;
            reg_file[28902] <= 8'h00;
            reg_file[28903] <= 8'h00;
            reg_file[28904] <= 8'h00;
            reg_file[28905] <= 8'h00;
            reg_file[28906] <= 8'h00;
            reg_file[28907] <= 8'h00;
            reg_file[28908] <= 8'h00;
            reg_file[28909] <= 8'h00;
            reg_file[28910] <= 8'h00;
            reg_file[28911] <= 8'h00;
            reg_file[28912] <= 8'h00;
            reg_file[28913] <= 8'h00;
            reg_file[28914] <= 8'h00;
            reg_file[28915] <= 8'h00;
            reg_file[28916] <= 8'h00;
            reg_file[28917] <= 8'h00;
            reg_file[28918] <= 8'h00;
            reg_file[28919] <= 8'h00;
            reg_file[28920] <= 8'h00;
            reg_file[28921] <= 8'h00;
            reg_file[28922] <= 8'h00;
            reg_file[28923] <= 8'h00;
            reg_file[28924] <= 8'h00;
            reg_file[28925] <= 8'h00;
            reg_file[28926] <= 8'h00;
            reg_file[28927] <= 8'h00;
            reg_file[28928] <= 8'h00;
            reg_file[28929] <= 8'h00;
            reg_file[28930] <= 8'h00;
            reg_file[28931] <= 8'h00;
            reg_file[28932] <= 8'h00;
            reg_file[28933] <= 8'h00;
            reg_file[28934] <= 8'h00;
            reg_file[28935] <= 8'h00;
            reg_file[28936] <= 8'h00;
            reg_file[28937] <= 8'h00;
            reg_file[28938] <= 8'h00;
            reg_file[28939] <= 8'h00;
            reg_file[28940] <= 8'h00;
            reg_file[28941] <= 8'h00;
            reg_file[28942] <= 8'h00;
            reg_file[28943] <= 8'h00;
            reg_file[28944] <= 8'h00;
            reg_file[28945] <= 8'h00;
            reg_file[28946] <= 8'h00;
            reg_file[28947] <= 8'h00;
            reg_file[28948] <= 8'h00;
            reg_file[28949] <= 8'h00;
            reg_file[28950] <= 8'h00;
            reg_file[28951] <= 8'h00;
            reg_file[28952] <= 8'h00;
            reg_file[28953] <= 8'h00;
            reg_file[28954] <= 8'h00;
            reg_file[28955] <= 8'h00;
            reg_file[28956] <= 8'h00;
            reg_file[28957] <= 8'h00;
            reg_file[28958] <= 8'h00;
            reg_file[28959] <= 8'h00;
            reg_file[28960] <= 8'h00;
            reg_file[28961] <= 8'h00;
            reg_file[28962] <= 8'h00;
            reg_file[28963] <= 8'h00;
            reg_file[28964] <= 8'h00;
            reg_file[28965] <= 8'h00;
            reg_file[28966] <= 8'h00;
            reg_file[28967] <= 8'h00;
            reg_file[28968] <= 8'h00;
            reg_file[28969] <= 8'h00;
            reg_file[28970] <= 8'h00;
            reg_file[28971] <= 8'h00;
            reg_file[28972] <= 8'h00;
            reg_file[28973] <= 8'h00;
            reg_file[28974] <= 8'h00;
            reg_file[28975] <= 8'h00;
            reg_file[28976] <= 8'h00;
            reg_file[28977] <= 8'h00;
            reg_file[28978] <= 8'h00;
            reg_file[28979] <= 8'h00;
            reg_file[28980] <= 8'h00;
            reg_file[28981] <= 8'h00;
            reg_file[28982] <= 8'h00;
            reg_file[28983] <= 8'h00;
            reg_file[28984] <= 8'h00;
            reg_file[28985] <= 8'h00;
            reg_file[28986] <= 8'h00;
            reg_file[28987] <= 8'h00;
            reg_file[28988] <= 8'h00;
            reg_file[28989] <= 8'h00;
            reg_file[28990] <= 8'h00;
            reg_file[28991] <= 8'h00;
            reg_file[28992] <= 8'h00;
            reg_file[28993] <= 8'h00;
            reg_file[28994] <= 8'h00;
            reg_file[28995] <= 8'h00;
            reg_file[28996] <= 8'h00;
            reg_file[28997] <= 8'h00;
            reg_file[28998] <= 8'h00;
            reg_file[28999] <= 8'h00;
            reg_file[29000] <= 8'h00;
            reg_file[29001] <= 8'h00;
            reg_file[29002] <= 8'h00;
            reg_file[29003] <= 8'h00;
            reg_file[29004] <= 8'h00;
            reg_file[29005] <= 8'h00;
            reg_file[29006] <= 8'h00;
            reg_file[29007] <= 8'h00;
            reg_file[29008] <= 8'h00;
            reg_file[29009] <= 8'h00;
            reg_file[29010] <= 8'h00;
            reg_file[29011] <= 8'h00;
            reg_file[29012] <= 8'h00;
            reg_file[29013] <= 8'h00;
            reg_file[29014] <= 8'h00;
            reg_file[29015] <= 8'h00;
            reg_file[29016] <= 8'h00;
            reg_file[29017] <= 8'h00;
            reg_file[29018] <= 8'h00;
            reg_file[29019] <= 8'h00;
            reg_file[29020] <= 8'h00;
            reg_file[29021] <= 8'h00;
            reg_file[29022] <= 8'h00;
            reg_file[29023] <= 8'h00;
            reg_file[29024] <= 8'h00;
            reg_file[29025] <= 8'h00;
            reg_file[29026] <= 8'h00;
            reg_file[29027] <= 8'h00;
            reg_file[29028] <= 8'h00;
            reg_file[29029] <= 8'h00;
            reg_file[29030] <= 8'h00;
            reg_file[29031] <= 8'h00;
            reg_file[29032] <= 8'h00;
            reg_file[29033] <= 8'h00;
            reg_file[29034] <= 8'h00;
            reg_file[29035] <= 8'h00;
            reg_file[29036] <= 8'h00;
            reg_file[29037] <= 8'h00;
            reg_file[29038] <= 8'h00;
            reg_file[29039] <= 8'h00;
            reg_file[29040] <= 8'h00;
            reg_file[29041] <= 8'h00;
            reg_file[29042] <= 8'h00;
            reg_file[29043] <= 8'h00;
            reg_file[29044] <= 8'h00;
            reg_file[29045] <= 8'h00;
            reg_file[29046] <= 8'h00;
            reg_file[29047] <= 8'h00;
            reg_file[29048] <= 8'h00;
            reg_file[29049] <= 8'h00;
            reg_file[29050] <= 8'h00;
            reg_file[29051] <= 8'h00;
            reg_file[29052] <= 8'h00;
            reg_file[29053] <= 8'h00;
            reg_file[29054] <= 8'h00;
            reg_file[29055] <= 8'h00;
            reg_file[29056] <= 8'h00;
            reg_file[29057] <= 8'h00;
            reg_file[29058] <= 8'h00;
            reg_file[29059] <= 8'h00;
            reg_file[29060] <= 8'h00;
            reg_file[29061] <= 8'h00;
            reg_file[29062] <= 8'h00;
            reg_file[29063] <= 8'h00;
            reg_file[29064] <= 8'h00;
            reg_file[29065] <= 8'h00;
            reg_file[29066] <= 8'h00;
            reg_file[29067] <= 8'h00;
            reg_file[29068] <= 8'h00;
            reg_file[29069] <= 8'h00;
            reg_file[29070] <= 8'h00;
            reg_file[29071] <= 8'h00;
            reg_file[29072] <= 8'h00;
            reg_file[29073] <= 8'h00;
            reg_file[29074] <= 8'h00;
            reg_file[29075] <= 8'h00;
            reg_file[29076] <= 8'h00;
            reg_file[29077] <= 8'h00;
            reg_file[29078] <= 8'h00;
            reg_file[29079] <= 8'h00;
            reg_file[29080] <= 8'h00;
            reg_file[29081] <= 8'h00;
            reg_file[29082] <= 8'h00;
            reg_file[29083] <= 8'h00;
            reg_file[29084] <= 8'h00;
            reg_file[29085] <= 8'h00;
            reg_file[29086] <= 8'h00;
            reg_file[29087] <= 8'h00;
            reg_file[29088] <= 8'h00;
            reg_file[29089] <= 8'h00;
            reg_file[29090] <= 8'h00;
            reg_file[29091] <= 8'h00;
            reg_file[29092] <= 8'h00;
            reg_file[29093] <= 8'h00;
            reg_file[29094] <= 8'h00;
            reg_file[29095] <= 8'h00;
            reg_file[29096] <= 8'h00;
            reg_file[29097] <= 8'h00;
            reg_file[29098] <= 8'h00;
            reg_file[29099] <= 8'h00;
            reg_file[29100] <= 8'h00;
            reg_file[29101] <= 8'h00;
            reg_file[29102] <= 8'h00;
            reg_file[29103] <= 8'h00;
            reg_file[29104] <= 8'h00;
            reg_file[29105] <= 8'h00;
            reg_file[29106] <= 8'h00;
            reg_file[29107] <= 8'h00;
            reg_file[29108] <= 8'h00;
            reg_file[29109] <= 8'h00;
            reg_file[29110] <= 8'h00;
            reg_file[29111] <= 8'h00;
            reg_file[29112] <= 8'h00;
            reg_file[29113] <= 8'h00;
            reg_file[29114] <= 8'h00;
            reg_file[29115] <= 8'h00;
            reg_file[29116] <= 8'h00;
            reg_file[29117] <= 8'h00;
            reg_file[29118] <= 8'h00;
            reg_file[29119] <= 8'h00;
            reg_file[29120] <= 8'h00;
            reg_file[29121] <= 8'h00;
            reg_file[29122] <= 8'h00;
            reg_file[29123] <= 8'h00;
            reg_file[29124] <= 8'h00;
            reg_file[29125] <= 8'h00;
            reg_file[29126] <= 8'h00;
            reg_file[29127] <= 8'h00;
            reg_file[29128] <= 8'h00;
            reg_file[29129] <= 8'h00;
            reg_file[29130] <= 8'h00;
            reg_file[29131] <= 8'h00;
            reg_file[29132] <= 8'h00;
            reg_file[29133] <= 8'h00;
            reg_file[29134] <= 8'h00;
            reg_file[29135] <= 8'h00;
            reg_file[29136] <= 8'h00;
            reg_file[29137] <= 8'h00;
            reg_file[29138] <= 8'h00;
            reg_file[29139] <= 8'h00;
            reg_file[29140] <= 8'h00;
            reg_file[29141] <= 8'h00;
            reg_file[29142] <= 8'h00;
            reg_file[29143] <= 8'h00;
            reg_file[29144] <= 8'h00;
            reg_file[29145] <= 8'h00;
            reg_file[29146] <= 8'h00;
            reg_file[29147] <= 8'h00;
            reg_file[29148] <= 8'h00;
            reg_file[29149] <= 8'h00;
            reg_file[29150] <= 8'h00;
            reg_file[29151] <= 8'h00;
            reg_file[29152] <= 8'h00;
            reg_file[29153] <= 8'h00;
            reg_file[29154] <= 8'h00;
            reg_file[29155] <= 8'h00;
            reg_file[29156] <= 8'h00;
            reg_file[29157] <= 8'h00;
            reg_file[29158] <= 8'h00;
            reg_file[29159] <= 8'h00;
            reg_file[29160] <= 8'h00;
            reg_file[29161] <= 8'h00;
            reg_file[29162] <= 8'h00;
            reg_file[29163] <= 8'h00;
            reg_file[29164] <= 8'h00;
            reg_file[29165] <= 8'h00;
            reg_file[29166] <= 8'h00;
            reg_file[29167] <= 8'h00;
            reg_file[29168] <= 8'h00;
            reg_file[29169] <= 8'h00;
            reg_file[29170] <= 8'h00;
            reg_file[29171] <= 8'h00;
            reg_file[29172] <= 8'h00;
            reg_file[29173] <= 8'h00;
            reg_file[29174] <= 8'h00;
            reg_file[29175] <= 8'h00;
            reg_file[29176] <= 8'h00;
            reg_file[29177] <= 8'h00;
            reg_file[29178] <= 8'h00;
            reg_file[29179] <= 8'h00;
            reg_file[29180] <= 8'h00;
            reg_file[29181] <= 8'h00;
            reg_file[29182] <= 8'h00;
            reg_file[29183] <= 8'h00;
            reg_file[29184] <= 8'h00;
            reg_file[29185] <= 8'h00;
            reg_file[29186] <= 8'h00;
            reg_file[29187] <= 8'h00;
            reg_file[29188] <= 8'h00;
            reg_file[29189] <= 8'h00;
            reg_file[29190] <= 8'h00;
            reg_file[29191] <= 8'h00;
            reg_file[29192] <= 8'h00;
            reg_file[29193] <= 8'h00;
            reg_file[29194] <= 8'h00;
            reg_file[29195] <= 8'h00;
            reg_file[29196] <= 8'h00;
            reg_file[29197] <= 8'h00;
            reg_file[29198] <= 8'h00;
            reg_file[29199] <= 8'h00;
            reg_file[29200] <= 8'h00;
            reg_file[29201] <= 8'h00;
            reg_file[29202] <= 8'h00;
            reg_file[29203] <= 8'h00;
            reg_file[29204] <= 8'h00;
            reg_file[29205] <= 8'h00;
            reg_file[29206] <= 8'h00;
            reg_file[29207] <= 8'h00;
            reg_file[29208] <= 8'h00;
            reg_file[29209] <= 8'h00;
            reg_file[29210] <= 8'h00;
            reg_file[29211] <= 8'h00;
            reg_file[29212] <= 8'h00;
            reg_file[29213] <= 8'h00;
            reg_file[29214] <= 8'h00;
            reg_file[29215] <= 8'h00;
            reg_file[29216] <= 8'h00;
            reg_file[29217] <= 8'h00;
            reg_file[29218] <= 8'h00;
            reg_file[29219] <= 8'h00;
            reg_file[29220] <= 8'h00;
            reg_file[29221] <= 8'h00;
            reg_file[29222] <= 8'h00;
            reg_file[29223] <= 8'h00;
            reg_file[29224] <= 8'h00;
            reg_file[29225] <= 8'h00;
            reg_file[29226] <= 8'h00;
            reg_file[29227] <= 8'h00;
            reg_file[29228] <= 8'h00;
            reg_file[29229] <= 8'h00;
            reg_file[29230] <= 8'h00;
            reg_file[29231] <= 8'h00;
            reg_file[29232] <= 8'h00;
            reg_file[29233] <= 8'h00;
            reg_file[29234] <= 8'h00;
            reg_file[29235] <= 8'h00;
            reg_file[29236] <= 8'h00;
            reg_file[29237] <= 8'h00;
            reg_file[29238] <= 8'h00;
            reg_file[29239] <= 8'h00;
            reg_file[29240] <= 8'h00;
            reg_file[29241] <= 8'h00;
            reg_file[29242] <= 8'h00;
            reg_file[29243] <= 8'h00;
            reg_file[29244] <= 8'h00;
            reg_file[29245] <= 8'h00;
            reg_file[29246] <= 8'h00;
            reg_file[29247] <= 8'h00;
            reg_file[29248] <= 8'h00;
            reg_file[29249] <= 8'h00;
            reg_file[29250] <= 8'h00;
            reg_file[29251] <= 8'h00;
            reg_file[29252] <= 8'h00;
            reg_file[29253] <= 8'h00;
            reg_file[29254] <= 8'h00;
            reg_file[29255] <= 8'h00;
            reg_file[29256] <= 8'h00;
            reg_file[29257] <= 8'h00;
            reg_file[29258] <= 8'h00;
            reg_file[29259] <= 8'h00;
            reg_file[29260] <= 8'h00;
            reg_file[29261] <= 8'h00;
            reg_file[29262] <= 8'h00;
            reg_file[29263] <= 8'h00;
            reg_file[29264] <= 8'h00;
            reg_file[29265] <= 8'h00;
            reg_file[29266] <= 8'h00;
            reg_file[29267] <= 8'h00;
            reg_file[29268] <= 8'h00;
            reg_file[29269] <= 8'h00;
            reg_file[29270] <= 8'h00;
            reg_file[29271] <= 8'h00;
            reg_file[29272] <= 8'h00;
            reg_file[29273] <= 8'h00;
            reg_file[29274] <= 8'h00;
            reg_file[29275] <= 8'h00;
            reg_file[29276] <= 8'h00;
            reg_file[29277] <= 8'h00;
            reg_file[29278] <= 8'h00;
            reg_file[29279] <= 8'h00;
            reg_file[29280] <= 8'h00;
            reg_file[29281] <= 8'h00;
            reg_file[29282] <= 8'h00;
            reg_file[29283] <= 8'h00;
            reg_file[29284] <= 8'h00;
            reg_file[29285] <= 8'h00;
            reg_file[29286] <= 8'h00;
            reg_file[29287] <= 8'h00;
            reg_file[29288] <= 8'h00;
            reg_file[29289] <= 8'h00;
            reg_file[29290] <= 8'h00;
            reg_file[29291] <= 8'h00;
            reg_file[29292] <= 8'h00;
            reg_file[29293] <= 8'h00;
            reg_file[29294] <= 8'h00;
            reg_file[29295] <= 8'h00;
            reg_file[29296] <= 8'h00;
            reg_file[29297] <= 8'h00;
            reg_file[29298] <= 8'h00;
            reg_file[29299] <= 8'h00;
            reg_file[29300] <= 8'h00;
            reg_file[29301] <= 8'h00;
            reg_file[29302] <= 8'h00;
            reg_file[29303] <= 8'h00;
            reg_file[29304] <= 8'h00;
            reg_file[29305] <= 8'h00;
            reg_file[29306] <= 8'h00;
            reg_file[29307] <= 8'h00;
            reg_file[29308] <= 8'h00;
            reg_file[29309] <= 8'h00;
            reg_file[29310] <= 8'h00;
            reg_file[29311] <= 8'h00;
            reg_file[29312] <= 8'h00;
            reg_file[29313] <= 8'h00;
            reg_file[29314] <= 8'h00;
            reg_file[29315] <= 8'h00;
            reg_file[29316] <= 8'h00;
            reg_file[29317] <= 8'h00;
            reg_file[29318] <= 8'h00;
            reg_file[29319] <= 8'h00;
            reg_file[29320] <= 8'h00;
            reg_file[29321] <= 8'h00;
            reg_file[29322] <= 8'h00;
            reg_file[29323] <= 8'h00;
            reg_file[29324] <= 8'h00;
            reg_file[29325] <= 8'h00;
            reg_file[29326] <= 8'h00;
            reg_file[29327] <= 8'h00;
            reg_file[29328] <= 8'h00;
            reg_file[29329] <= 8'h00;
            reg_file[29330] <= 8'h00;
            reg_file[29331] <= 8'h00;
            reg_file[29332] <= 8'h00;
            reg_file[29333] <= 8'h00;
            reg_file[29334] <= 8'h00;
            reg_file[29335] <= 8'h00;
            reg_file[29336] <= 8'h00;
            reg_file[29337] <= 8'h00;
            reg_file[29338] <= 8'h00;
            reg_file[29339] <= 8'h00;
            reg_file[29340] <= 8'h00;
            reg_file[29341] <= 8'h00;
            reg_file[29342] <= 8'h00;
            reg_file[29343] <= 8'h00;
            reg_file[29344] <= 8'h00;
            reg_file[29345] <= 8'h00;
            reg_file[29346] <= 8'h00;
            reg_file[29347] <= 8'h00;
            reg_file[29348] <= 8'h00;
            reg_file[29349] <= 8'h00;
            reg_file[29350] <= 8'h00;
            reg_file[29351] <= 8'h00;
            reg_file[29352] <= 8'h00;
            reg_file[29353] <= 8'h00;
            reg_file[29354] <= 8'h00;
            reg_file[29355] <= 8'h00;
            reg_file[29356] <= 8'h00;
            reg_file[29357] <= 8'h00;
            reg_file[29358] <= 8'h00;
            reg_file[29359] <= 8'h00;
            reg_file[29360] <= 8'h00;
            reg_file[29361] <= 8'h00;
            reg_file[29362] <= 8'h00;
            reg_file[29363] <= 8'h00;
            reg_file[29364] <= 8'h00;
            reg_file[29365] <= 8'h00;
            reg_file[29366] <= 8'h00;
            reg_file[29367] <= 8'h00;
            reg_file[29368] <= 8'h00;
            reg_file[29369] <= 8'h00;
            reg_file[29370] <= 8'h00;
            reg_file[29371] <= 8'h00;
            reg_file[29372] <= 8'h00;
            reg_file[29373] <= 8'h00;
            reg_file[29374] <= 8'h00;
            reg_file[29375] <= 8'h00;
            reg_file[29376] <= 8'h00;
            reg_file[29377] <= 8'h00;
            reg_file[29378] <= 8'h00;
            reg_file[29379] <= 8'h00;
            reg_file[29380] <= 8'h00;
            reg_file[29381] <= 8'h00;
            reg_file[29382] <= 8'h00;
            reg_file[29383] <= 8'h00;
            reg_file[29384] <= 8'h00;
            reg_file[29385] <= 8'h00;
            reg_file[29386] <= 8'h00;
            reg_file[29387] <= 8'h00;
            reg_file[29388] <= 8'h00;
            reg_file[29389] <= 8'h00;
            reg_file[29390] <= 8'h00;
            reg_file[29391] <= 8'h00;
            reg_file[29392] <= 8'h00;
            reg_file[29393] <= 8'h00;
            reg_file[29394] <= 8'h00;
            reg_file[29395] <= 8'h00;
            reg_file[29396] <= 8'h00;
            reg_file[29397] <= 8'h00;
            reg_file[29398] <= 8'h00;
            reg_file[29399] <= 8'h00;
            reg_file[29400] <= 8'h00;
            reg_file[29401] <= 8'h00;
            reg_file[29402] <= 8'h00;
            reg_file[29403] <= 8'h00;
            reg_file[29404] <= 8'h00;
            reg_file[29405] <= 8'h00;
            reg_file[29406] <= 8'h00;
            reg_file[29407] <= 8'h00;
            reg_file[29408] <= 8'h00;
            reg_file[29409] <= 8'h00;
            reg_file[29410] <= 8'h00;
            reg_file[29411] <= 8'h00;
            reg_file[29412] <= 8'h00;
            reg_file[29413] <= 8'h00;
            reg_file[29414] <= 8'h00;
            reg_file[29415] <= 8'h00;
            reg_file[29416] <= 8'h00;
            reg_file[29417] <= 8'h00;
            reg_file[29418] <= 8'h00;
            reg_file[29419] <= 8'h00;
            reg_file[29420] <= 8'h00;
            reg_file[29421] <= 8'h00;
            reg_file[29422] <= 8'h00;
            reg_file[29423] <= 8'h00;
            reg_file[29424] <= 8'h00;
            reg_file[29425] <= 8'h00;
            reg_file[29426] <= 8'h00;
            reg_file[29427] <= 8'h00;
            reg_file[29428] <= 8'h00;
            reg_file[29429] <= 8'h00;
            reg_file[29430] <= 8'h00;
            reg_file[29431] <= 8'h00;
            reg_file[29432] <= 8'h00;
            reg_file[29433] <= 8'h00;
            reg_file[29434] <= 8'h00;
            reg_file[29435] <= 8'h00;
            reg_file[29436] <= 8'h00;
            reg_file[29437] <= 8'h00;
            reg_file[29438] <= 8'h00;
            reg_file[29439] <= 8'h00;
            reg_file[29440] <= 8'h00;
            reg_file[29441] <= 8'h00;
            reg_file[29442] <= 8'h00;
            reg_file[29443] <= 8'h00;
            reg_file[29444] <= 8'h00;
            reg_file[29445] <= 8'h00;
            reg_file[29446] <= 8'h00;
            reg_file[29447] <= 8'h00;
            reg_file[29448] <= 8'h00;
            reg_file[29449] <= 8'h00;
            reg_file[29450] <= 8'h00;
            reg_file[29451] <= 8'h00;
            reg_file[29452] <= 8'h00;
            reg_file[29453] <= 8'h00;
            reg_file[29454] <= 8'h00;
            reg_file[29455] <= 8'h00;
            reg_file[29456] <= 8'h00;
            reg_file[29457] <= 8'h00;
            reg_file[29458] <= 8'h00;
            reg_file[29459] <= 8'h00;
            reg_file[29460] <= 8'h00;
            reg_file[29461] <= 8'h00;
            reg_file[29462] <= 8'h00;
            reg_file[29463] <= 8'h00;
            reg_file[29464] <= 8'h00;
            reg_file[29465] <= 8'h00;
            reg_file[29466] <= 8'h00;
            reg_file[29467] <= 8'h00;
            reg_file[29468] <= 8'h00;
            reg_file[29469] <= 8'h00;
            reg_file[29470] <= 8'h00;
            reg_file[29471] <= 8'h00;
            reg_file[29472] <= 8'h00;
            reg_file[29473] <= 8'h00;
            reg_file[29474] <= 8'h00;
            reg_file[29475] <= 8'h00;
            reg_file[29476] <= 8'h00;
            reg_file[29477] <= 8'h00;
            reg_file[29478] <= 8'h00;
            reg_file[29479] <= 8'h00;
            reg_file[29480] <= 8'h00;
            reg_file[29481] <= 8'h00;
            reg_file[29482] <= 8'h00;
            reg_file[29483] <= 8'h00;
            reg_file[29484] <= 8'h00;
            reg_file[29485] <= 8'h00;
            reg_file[29486] <= 8'h00;
            reg_file[29487] <= 8'h00;
            reg_file[29488] <= 8'h00;
            reg_file[29489] <= 8'h00;
            reg_file[29490] <= 8'h00;
            reg_file[29491] <= 8'h00;
            reg_file[29492] <= 8'h00;
            reg_file[29493] <= 8'h00;
            reg_file[29494] <= 8'h00;
            reg_file[29495] <= 8'h00;
            reg_file[29496] <= 8'h00;
            reg_file[29497] <= 8'h00;
            reg_file[29498] <= 8'h00;
            reg_file[29499] <= 8'h00;
            reg_file[29500] <= 8'h00;
            reg_file[29501] <= 8'h00;
            reg_file[29502] <= 8'h00;
            reg_file[29503] <= 8'h00;
            reg_file[29504] <= 8'h00;
            reg_file[29505] <= 8'h00;
            reg_file[29506] <= 8'h00;
            reg_file[29507] <= 8'h00;
            reg_file[29508] <= 8'h00;
            reg_file[29509] <= 8'h00;
            reg_file[29510] <= 8'h00;
            reg_file[29511] <= 8'h00;
            reg_file[29512] <= 8'h00;
            reg_file[29513] <= 8'h00;
            reg_file[29514] <= 8'h00;
            reg_file[29515] <= 8'h00;
            reg_file[29516] <= 8'h00;
            reg_file[29517] <= 8'h00;
            reg_file[29518] <= 8'h00;
            reg_file[29519] <= 8'h00;
            reg_file[29520] <= 8'h00;
            reg_file[29521] <= 8'h00;
            reg_file[29522] <= 8'h00;
            reg_file[29523] <= 8'h00;
            reg_file[29524] <= 8'h00;
            reg_file[29525] <= 8'h00;
            reg_file[29526] <= 8'h00;
            reg_file[29527] <= 8'h00;
            reg_file[29528] <= 8'h00;
            reg_file[29529] <= 8'h00;
            reg_file[29530] <= 8'h00;
            reg_file[29531] <= 8'h00;
            reg_file[29532] <= 8'h00;
            reg_file[29533] <= 8'h00;
            reg_file[29534] <= 8'h00;
            reg_file[29535] <= 8'h00;
            reg_file[29536] <= 8'h00;
            reg_file[29537] <= 8'h00;
            reg_file[29538] <= 8'h00;
            reg_file[29539] <= 8'h00;
            reg_file[29540] <= 8'h00;
            reg_file[29541] <= 8'h00;
            reg_file[29542] <= 8'h00;
            reg_file[29543] <= 8'h00;
            reg_file[29544] <= 8'h00;
            reg_file[29545] <= 8'h00;
            reg_file[29546] <= 8'h00;
            reg_file[29547] <= 8'h00;
            reg_file[29548] <= 8'h00;
            reg_file[29549] <= 8'h00;
            reg_file[29550] <= 8'h00;
            reg_file[29551] <= 8'h00;
            reg_file[29552] <= 8'h00;
            reg_file[29553] <= 8'h00;
            reg_file[29554] <= 8'h00;
            reg_file[29555] <= 8'h00;
            reg_file[29556] <= 8'h00;
            reg_file[29557] <= 8'h00;
            reg_file[29558] <= 8'h00;
            reg_file[29559] <= 8'h00;
            reg_file[29560] <= 8'h00;
            reg_file[29561] <= 8'h00;
            reg_file[29562] <= 8'h00;
            reg_file[29563] <= 8'h00;
            reg_file[29564] <= 8'h00;
            reg_file[29565] <= 8'h00;
            reg_file[29566] <= 8'h00;
            reg_file[29567] <= 8'h00;
            reg_file[29568] <= 8'h00;
            reg_file[29569] <= 8'h00;
            reg_file[29570] <= 8'h00;
            reg_file[29571] <= 8'h00;
            reg_file[29572] <= 8'h00;
            reg_file[29573] <= 8'h00;
            reg_file[29574] <= 8'h00;
            reg_file[29575] <= 8'h00;
            reg_file[29576] <= 8'h00;
            reg_file[29577] <= 8'h00;
            reg_file[29578] <= 8'h00;
            reg_file[29579] <= 8'h00;
            reg_file[29580] <= 8'h00;
            reg_file[29581] <= 8'h00;
            reg_file[29582] <= 8'h00;
            reg_file[29583] <= 8'h00;
            reg_file[29584] <= 8'h00;
            reg_file[29585] <= 8'h00;
            reg_file[29586] <= 8'h00;
            reg_file[29587] <= 8'h00;
            reg_file[29588] <= 8'h00;
            reg_file[29589] <= 8'h00;
            reg_file[29590] <= 8'h00;
            reg_file[29591] <= 8'h00;
            reg_file[29592] <= 8'h00;
            reg_file[29593] <= 8'h00;
            reg_file[29594] <= 8'h00;
            reg_file[29595] <= 8'h00;
            reg_file[29596] <= 8'h00;
            reg_file[29597] <= 8'h00;
            reg_file[29598] <= 8'h00;
            reg_file[29599] <= 8'h00;
            reg_file[29600] <= 8'h00;
            reg_file[29601] <= 8'h00;
            reg_file[29602] <= 8'h00;
            reg_file[29603] <= 8'h00;
            reg_file[29604] <= 8'h00;
            reg_file[29605] <= 8'h00;
            reg_file[29606] <= 8'h00;
            reg_file[29607] <= 8'h00;
            reg_file[29608] <= 8'h00;
            reg_file[29609] <= 8'h00;
            reg_file[29610] <= 8'h00;
            reg_file[29611] <= 8'h00;
            reg_file[29612] <= 8'h00;
            reg_file[29613] <= 8'h00;
            reg_file[29614] <= 8'h00;
            reg_file[29615] <= 8'h00;
            reg_file[29616] <= 8'h00;
            reg_file[29617] <= 8'h00;
            reg_file[29618] <= 8'h00;
            reg_file[29619] <= 8'h00;
            reg_file[29620] <= 8'h00;
            reg_file[29621] <= 8'h00;
            reg_file[29622] <= 8'h00;
            reg_file[29623] <= 8'h00;
            reg_file[29624] <= 8'h00;
            reg_file[29625] <= 8'h00;
            reg_file[29626] <= 8'h00;
            reg_file[29627] <= 8'h00;
            reg_file[29628] <= 8'h00;
            reg_file[29629] <= 8'h00;
            reg_file[29630] <= 8'h00;
            reg_file[29631] <= 8'h00;
            reg_file[29632] <= 8'h00;
            reg_file[29633] <= 8'h00;
            reg_file[29634] <= 8'h00;
            reg_file[29635] <= 8'h00;
            reg_file[29636] <= 8'h00;
            reg_file[29637] <= 8'h00;
            reg_file[29638] <= 8'h00;
            reg_file[29639] <= 8'h00;
            reg_file[29640] <= 8'h00;
            reg_file[29641] <= 8'h00;
            reg_file[29642] <= 8'h00;
            reg_file[29643] <= 8'h00;
            reg_file[29644] <= 8'h00;
            reg_file[29645] <= 8'h00;
            reg_file[29646] <= 8'h00;
            reg_file[29647] <= 8'h00;
            reg_file[29648] <= 8'h00;
            reg_file[29649] <= 8'h00;
            reg_file[29650] <= 8'h00;
            reg_file[29651] <= 8'h00;
            reg_file[29652] <= 8'h00;
            reg_file[29653] <= 8'h00;
            reg_file[29654] <= 8'h00;
            reg_file[29655] <= 8'h00;
            reg_file[29656] <= 8'h00;
            reg_file[29657] <= 8'h00;
            reg_file[29658] <= 8'h00;
            reg_file[29659] <= 8'h00;
            reg_file[29660] <= 8'h00;
            reg_file[29661] <= 8'h00;
            reg_file[29662] <= 8'h00;
            reg_file[29663] <= 8'h00;
            reg_file[29664] <= 8'h00;
            reg_file[29665] <= 8'h00;
            reg_file[29666] <= 8'h00;
            reg_file[29667] <= 8'h00;
            reg_file[29668] <= 8'h00;
            reg_file[29669] <= 8'h00;
            reg_file[29670] <= 8'h00;
            reg_file[29671] <= 8'h00;
            reg_file[29672] <= 8'h00;
            reg_file[29673] <= 8'h00;
            reg_file[29674] <= 8'h00;
            reg_file[29675] <= 8'h00;
            reg_file[29676] <= 8'h00;
            reg_file[29677] <= 8'h00;
            reg_file[29678] <= 8'h00;
            reg_file[29679] <= 8'h00;
            reg_file[29680] <= 8'h00;
            reg_file[29681] <= 8'h00;
            reg_file[29682] <= 8'h00;
            reg_file[29683] <= 8'h00;
            reg_file[29684] <= 8'h00;
            reg_file[29685] <= 8'h00;
            reg_file[29686] <= 8'h00;
            reg_file[29687] <= 8'h00;
            reg_file[29688] <= 8'h00;
            reg_file[29689] <= 8'h00;
            reg_file[29690] <= 8'h00;
            reg_file[29691] <= 8'h00;
            reg_file[29692] <= 8'h00;
            reg_file[29693] <= 8'h00;
            reg_file[29694] <= 8'h00;
            reg_file[29695] <= 8'h00;
            reg_file[29696] <= 8'h00;
            reg_file[29697] <= 8'h00;
            reg_file[29698] <= 8'h00;
            reg_file[29699] <= 8'h00;
            reg_file[29700] <= 8'h00;
            reg_file[29701] <= 8'h00;
            reg_file[29702] <= 8'h00;
            reg_file[29703] <= 8'h00;
            reg_file[29704] <= 8'h00;
            reg_file[29705] <= 8'h00;
            reg_file[29706] <= 8'h00;
            reg_file[29707] <= 8'h00;
            reg_file[29708] <= 8'h00;
            reg_file[29709] <= 8'h00;
            reg_file[29710] <= 8'h00;
            reg_file[29711] <= 8'h00;
            reg_file[29712] <= 8'h00;
            reg_file[29713] <= 8'h00;
            reg_file[29714] <= 8'h00;
            reg_file[29715] <= 8'h00;
            reg_file[29716] <= 8'h00;
            reg_file[29717] <= 8'h00;
            reg_file[29718] <= 8'h00;
            reg_file[29719] <= 8'h00;
            reg_file[29720] <= 8'h00;
            reg_file[29721] <= 8'h00;
            reg_file[29722] <= 8'h00;
            reg_file[29723] <= 8'h00;
            reg_file[29724] <= 8'h00;
            reg_file[29725] <= 8'h00;
            reg_file[29726] <= 8'h00;
            reg_file[29727] <= 8'h00;
            reg_file[29728] <= 8'h00;
            reg_file[29729] <= 8'h00;
            reg_file[29730] <= 8'h00;
            reg_file[29731] <= 8'h00;
            reg_file[29732] <= 8'h00;
            reg_file[29733] <= 8'h00;
            reg_file[29734] <= 8'h00;
            reg_file[29735] <= 8'h00;
            reg_file[29736] <= 8'h00;
            reg_file[29737] <= 8'h00;
            reg_file[29738] <= 8'h00;
            reg_file[29739] <= 8'h00;
            reg_file[29740] <= 8'h00;
            reg_file[29741] <= 8'h00;
            reg_file[29742] <= 8'h00;
            reg_file[29743] <= 8'h00;
            reg_file[29744] <= 8'h00;
            reg_file[29745] <= 8'h00;
            reg_file[29746] <= 8'h00;
            reg_file[29747] <= 8'h00;
            reg_file[29748] <= 8'h00;
            reg_file[29749] <= 8'h00;
            reg_file[29750] <= 8'h00;
            reg_file[29751] <= 8'h00;
            reg_file[29752] <= 8'h00;
            reg_file[29753] <= 8'h00;
            reg_file[29754] <= 8'h00;
            reg_file[29755] <= 8'h00;
            reg_file[29756] <= 8'h00;
            reg_file[29757] <= 8'h00;
            reg_file[29758] <= 8'h00;
            reg_file[29759] <= 8'h00;
            reg_file[29760] <= 8'h00;
            reg_file[29761] <= 8'h00;
            reg_file[29762] <= 8'h00;
            reg_file[29763] <= 8'h00;
            reg_file[29764] <= 8'h00;
            reg_file[29765] <= 8'h00;
            reg_file[29766] <= 8'h00;
            reg_file[29767] <= 8'h00;
            reg_file[29768] <= 8'h00;
            reg_file[29769] <= 8'h00;
            reg_file[29770] <= 8'h00;
            reg_file[29771] <= 8'h00;
            reg_file[29772] <= 8'h00;
            reg_file[29773] <= 8'h00;
            reg_file[29774] <= 8'h00;
            reg_file[29775] <= 8'h00;
            reg_file[29776] <= 8'h00;
            reg_file[29777] <= 8'h00;
            reg_file[29778] <= 8'h00;
            reg_file[29779] <= 8'h00;
            reg_file[29780] <= 8'h00;
            reg_file[29781] <= 8'h00;
            reg_file[29782] <= 8'h00;
            reg_file[29783] <= 8'h00;
            reg_file[29784] <= 8'h00;
            reg_file[29785] <= 8'h00;
            reg_file[29786] <= 8'h00;
            reg_file[29787] <= 8'h00;
            reg_file[29788] <= 8'h00;
            reg_file[29789] <= 8'h00;
            reg_file[29790] <= 8'h00;
            reg_file[29791] <= 8'h00;
            reg_file[29792] <= 8'h00;
            reg_file[29793] <= 8'h00;
            reg_file[29794] <= 8'h00;
            reg_file[29795] <= 8'h00;
            reg_file[29796] <= 8'h00;
            reg_file[29797] <= 8'h00;
            reg_file[29798] <= 8'h00;
            reg_file[29799] <= 8'h00;
            reg_file[29800] <= 8'h00;
            reg_file[29801] <= 8'h00;
            reg_file[29802] <= 8'h00;
            reg_file[29803] <= 8'h00;
            reg_file[29804] <= 8'h00;
            reg_file[29805] <= 8'h00;
            reg_file[29806] <= 8'h00;
            reg_file[29807] <= 8'h00;
            reg_file[29808] <= 8'h00;
            reg_file[29809] <= 8'h00;
            reg_file[29810] <= 8'h00;
            reg_file[29811] <= 8'h00;
            reg_file[29812] <= 8'h00;
            reg_file[29813] <= 8'h00;
            reg_file[29814] <= 8'h00;
            reg_file[29815] <= 8'h00;
            reg_file[29816] <= 8'h00;
            reg_file[29817] <= 8'h00;
            reg_file[29818] <= 8'h00;
            reg_file[29819] <= 8'h00;
            reg_file[29820] <= 8'h00;
            reg_file[29821] <= 8'h00;
            reg_file[29822] <= 8'h00;
            reg_file[29823] <= 8'h00;
            reg_file[29824] <= 8'h00;
            reg_file[29825] <= 8'h00;
            reg_file[29826] <= 8'h00;
            reg_file[29827] <= 8'h00;
            reg_file[29828] <= 8'h00;
            reg_file[29829] <= 8'h00;
            reg_file[29830] <= 8'h00;
            reg_file[29831] <= 8'h00;
            reg_file[29832] <= 8'h00;
            reg_file[29833] <= 8'h00;
            reg_file[29834] <= 8'h00;
            reg_file[29835] <= 8'h00;
            reg_file[29836] <= 8'h00;
            reg_file[29837] <= 8'h00;
            reg_file[29838] <= 8'h00;
            reg_file[29839] <= 8'h00;
            reg_file[29840] <= 8'h00;
            reg_file[29841] <= 8'h00;
            reg_file[29842] <= 8'h00;
            reg_file[29843] <= 8'h00;
            reg_file[29844] <= 8'h00;
            reg_file[29845] <= 8'h00;
            reg_file[29846] <= 8'h00;
            reg_file[29847] <= 8'h00;
            reg_file[29848] <= 8'h00;
            reg_file[29849] <= 8'h00;
            reg_file[29850] <= 8'h00;
            reg_file[29851] <= 8'h00;
            reg_file[29852] <= 8'h00;
            reg_file[29853] <= 8'h00;
            reg_file[29854] <= 8'h00;
            reg_file[29855] <= 8'h00;
            reg_file[29856] <= 8'h00;
            reg_file[29857] <= 8'h00;
            reg_file[29858] <= 8'h00;
            reg_file[29859] <= 8'h00;
            reg_file[29860] <= 8'h00;
            reg_file[29861] <= 8'h00;
            reg_file[29862] <= 8'h00;
            reg_file[29863] <= 8'h00;
            reg_file[29864] <= 8'h00;
            reg_file[29865] <= 8'h00;
            reg_file[29866] <= 8'h00;
            reg_file[29867] <= 8'h00;
            reg_file[29868] <= 8'h00;
            reg_file[29869] <= 8'h00;
            reg_file[29870] <= 8'h00;
            reg_file[29871] <= 8'h00;
            reg_file[29872] <= 8'h00;
            reg_file[29873] <= 8'h00;
            reg_file[29874] <= 8'h00;
            reg_file[29875] <= 8'h00;
            reg_file[29876] <= 8'h00;
            reg_file[29877] <= 8'h00;
            reg_file[29878] <= 8'h00;
            reg_file[29879] <= 8'h00;
            reg_file[29880] <= 8'h00;
            reg_file[29881] <= 8'h00;
            reg_file[29882] <= 8'h00;
            reg_file[29883] <= 8'h00;
            reg_file[29884] <= 8'h00;
            reg_file[29885] <= 8'h00;
            reg_file[29886] <= 8'h00;
            reg_file[29887] <= 8'h00;
            reg_file[29888] <= 8'h00;
            reg_file[29889] <= 8'h00;
            reg_file[29890] <= 8'h00;
            reg_file[29891] <= 8'h00;
            reg_file[29892] <= 8'h00;
            reg_file[29893] <= 8'h00;
            reg_file[29894] <= 8'h00;
            reg_file[29895] <= 8'h00;
            reg_file[29896] <= 8'h00;
            reg_file[29897] <= 8'h00;
            reg_file[29898] <= 8'h00;
            reg_file[29899] <= 8'h00;
            reg_file[29900] <= 8'h00;
            reg_file[29901] <= 8'h00;
            reg_file[29902] <= 8'h00;
            reg_file[29903] <= 8'h00;
            reg_file[29904] <= 8'h00;
            reg_file[29905] <= 8'h00;
            reg_file[29906] <= 8'h00;
            reg_file[29907] <= 8'h00;
            reg_file[29908] <= 8'h00;
            reg_file[29909] <= 8'h00;
            reg_file[29910] <= 8'h00;
            reg_file[29911] <= 8'h00;
            reg_file[29912] <= 8'h00;
            reg_file[29913] <= 8'h00;
            reg_file[29914] <= 8'h00;
            reg_file[29915] <= 8'h00;
            reg_file[29916] <= 8'h00;
            reg_file[29917] <= 8'h00;
            reg_file[29918] <= 8'h00;
            reg_file[29919] <= 8'h00;
            reg_file[29920] <= 8'h00;
            reg_file[29921] <= 8'h00;
            reg_file[29922] <= 8'h00;
            reg_file[29923] <= 8'h00;
            reg_file[29924] <= 8'h00;
            reg_file[29925] <= 8'h00;
            reg_file[29926] <= 8'h00;
            reg_file[29927] <= 8'h00;
            reg_file[29928] <= 8'h00;
            reg_file[29929] <= 8'h00;
            reg_file[29930] <= 8'h00;
            reg_file[29931] <= 8'h00;
            reg_file[29932] <= 8'h00;
            reg_file[29933] <= 8'h00;
            reg_file[29934] <= 8'h00;
            reg_file[29935] <= 8'h00;
            reg_file[29936] <= 8'h00;
            reg_file[29937] <= 8'h00;
            reg_file[29938] <= 8'h00;
            reg_file[29939] <= 8'h00;
            reg_file[29940] <= 8'h00;
            reg_file[29941] <= 8'h00;
            reg_file[29942] <= 8'h00;
            reg_file[29943] <= 8'h00;
            reg_file[29944] <= 8'h00;
            reg_file[29945] <= 8'h00;
            reg_file[29946] <= 8'h00;
            reg_file[29947] <= 8'h00;
            reg_file[29948] <= 8'h00;
            reg_file[29949] <= 8'h00;
            reg_file[29950] <= 8'h00;
            reg_file[29951] <= 8'h00;
            reg_file[29952] <= 8'h00;
            reg_file[29953] <= 8'h00;
            reg_file[29954] <= 8'h00;
            reg_file[29955] <= 8'h00;
            reg_file[29956] <= 8'h00;
            reg_file[29957] <= 8'h00;
            reg_file[29958] <= 8'h00;
            reg_file[29959] <= 8'h00;
            reg_file[29960] <= 8'h00;
            reg_file[29961] <= 8'h00;
            reg_file[29962] <= 8'h00;
            reg_file[29963] <= 8'h00;
            reg_file[29964] <= 8'h00;
            reg_file[29965] <= 8'h00;
            reg_file[29966] <= 8'h00;
            reg_file[29967] <= 8'h00;
            reg_file[29968] <= 8'h00;
            reg_file[29969] <= 8'h00;
            reg_file[29970] <= 8'h00;
            reg_file[29971] <= 8'h00;
            reg_file[29972] <= 8'h00;
            reg_file[29973] <= 8'h00;
            reg_file[29974] <= 8'h00;
            reg_file[29975] <= 8'h00;
            reg_file[29976] <= 8'h00;
            reg_file[29977] <= 8'h00;
            reg_file[29978] <= 8'h00;
            reg_file[29979] <= 8'h00;
            reg_file[29980] <= 8'h00;
            reg_file[29981] <= 8'h00;
            reg_file[29982] <= 8'h00;
            reg_file[29983] <= 8'h00;
            reg_file[29984] <= 8'h00;
            reg_file[29985] <= 8'h00;
            reg_file[29986] <= 8'h00;
            reg_file[29987] <= 8'h00;
            reg_file[29988] <= 8'h00;
            reg_file[29989] <= 8'h00;
            reg_file[29990] <= 8'h00;
            reg_file[29991] <= 8'h00;
            reg_file[29992] <= 8'h00;
            reg_file[29993] <= 8'h00;
            reg_file[29994] <= 8'h00;
            reg_file[29995] <= 8'h00;
            reg_file[29996] <= 8'h00;
            reg_file[29997] <= 8'h00;
            reg_file[29998] <= 8'h00;
            reg_file[29999] <= 8'h00;
            reg_file[30000] <= 8'h00;
            reg_file[30001] <= 8'h00;
            reg_file[30002] <= 8'h00;
            reg_file[30003] <= 8'h00;
            reg_file[30004] <= 8'h00;
            reg_file[30005] <= 8'h00;
            reg_file[30006] <= 8'h00;
            reg_file[30007] <= 8'h00;
            reg_file[30008] <= 8'h00;
            reg_file[30009] <= 8'h00;
            reg_file[30010] <= 8'h00;
            reg_file[30011] <= 8'h00;
            reg_file[30012] <= 8'h00;
            reg_file[30013] <= 8'h00;
            reg_file[30014] <= 8'h00;
            reg_file[30015] <= 8'h00;
            reg_file[30016] <= 8'h00;
            reg_file[30017] <= 8'h00;
            reg_file[30018] <= 8'h00;
            reg_file[30019] <= 8'h00;
            reg_file[30020] <= 8'h00;
            reg_file[30021] <= 8'h00;
            reg_file[30022] <= 8'h00;
            reg_file[30023] <= 8'h00;
            reg_file[30024] <= 8'h00;
            reg_file[30025] <= 8'h00;
            reg_file[30026] <= 8'h00;
            reg_file[30027] <= 8'h00;
            reg_file[30028] <= 8'h00;
            reg_file[30029] <= 8'h00;
            reg_file[30030] <= 8'h00;
            reg_file[30031] <= 8'h00;
            reg_file[30032] <= 8'h00;
            reg_file[30033] <= 8'h00;
            reg_file[30034] <= 8'h00;
            reg_file[30035] <= 8'h00;
            reg_file[30036] <= 8'h00;
            reg_file[30037] <= 8'h00;
            reg_file[30038] <= 8'h00;
            reg_file[30039] <= 8'h00;
            reg_file[30040] <= 8'h00;
            reg_file[30041] <= 8'h00;
            reg_file[30042] <= 8'h00;
            reg_file[30043] <= 8'h00;
            reg_file[30044] <= 8'h00;
            reg_file[30045] <= 8'h00;
            reg_file[30046] <= 8'h00;
            reg_file[30047] <= 8'h00;
            reg_file[30048] <= 8'h00;
            reg_file[30049] <= 8'h00;
            reg_file[30050] <= 8'h00;
            reg_file[30051] <= 8'h00;
            reg_file[30052] <= 8'h00;
            reg_file[30053] <= 8'h00;
            reg_file[30054] <= 8'h00;
            reg_file[30055] <= 8'h00;
            reg_file[30056] <= 8'h00;
            reg_file[30057] <= 8'h00;
            reg_file[30058] <= 8'h00;
            reg_file[30059] <= 8'h00;
            reg_file[30060] <= 8'h00;
            reg_file[30061] <= 8'h00;
            reg_file[30062] <= 8'h00;
            reg_file[30063] <= 8'h00;
            reg_file[30064] <= 8'h00;
            reg_file[30065] <= 8'h00;
            reg_file[30066] <= 8'h00;
            reg_file[30067] <= 8'h00;
            reg_file[30068] <= 8'h00;
            reg_file[30069] <= 8'h00;
            reg_file[30070] <= 8'h00;
            reg_file[30071] <= 8'h00;
            reg_file[30072] <= 8'h00;
            reg_file[30073] <= 8'h00;
            reg_file[30074] <= 8'h00;
            reg_file[30075] <= 8'h00;
            reg_file[30076] <= 8'h00;
            reg_file[30077] <= 8'h00;
            reg_file[30078] <= 8'h00;
            reg_file[30079] <= 8'h00;
            reg_file[30080] <= 8'h00;
            reg_file[30081] <= 8'h00;
            reg_file[30082] <= 8'h00;
            reg_file[30083] <= 8'h00;
            reg_file[30084] <= 8'h00;
            reg_file[30085] <= 8'h00;
            reg_file[30086] <= 8'h00;
            reg_file[30087] <= 8'h00;
            reg_file[30088] <= 8'h00;
            reg_file[30089] <= 8'h00;
            reg_file[30090] <= 8'h00;
            reg_file[30091] <= 8'h00;
            reg_file[30092] <= 8'h00;
            reg_file[30093] <= 8'h00;
            reg_file[30094] <= 8'h00;
            reg_file[30095] <= 8'h00;
            reg_file[30096] <= 8'h00;
            reg_file[30097] <= 8'h00;
            reg_file[30098] <= 8'h00;
            reg_file[30099] <= 8'h00;
            reg_file[30100] <= 8'h00;
            reg_file[30101] <= 8'h00;
            reg_file[30102] <= 8'h00;
            reg_file[30103] <= 8'h00;
            reg_file[30104] <= 8'h00;
            reg_file[30105] <= 8'h00;
            reg_file[30106] <= 8'h00;
            reg_file[30107] <= 8'h00;
            reg_file[30108] <= 8'h00;
            reg_file[30109] <= 8'h00;
            reg_file[30110] <= 8'h00;
            reg_file[30111] <= 8'h00;
            reg_file[30112] <= 8'h00;
            reg_file[30113] <= 8'h00;
            reg_file[30114] <= 8'h00;
            reg_file[30115] <= 8'h00;
            reg_file[30116] <= 8'h00;
            reg_file[30117] <= 8'h00;
            reg_file[30118] <= 8'h00;
            reg_file[30119] <= 8'h00;
            reg_file[30120] <= 8'h00;
            reg_file[30121] <= 8'h00;
            reg_file[30122] <= 8'h00;
            reg_file[30123] <= 8'h00;
            reg_file[30124] <= 8'h00;
            reg_file[30125] <= 8'h00;
            reg_file[30126] <= 8'h00;
            reg_file[30127] <= 8'h00;
            reg_file[30128] <= 8'h00;
            reg_file[30129] <= 8'h00;
            reg_file[30130] <= 8'h00;
            reg_file[30131] <= 8'h00;
            reg_file[30132] <= 8'h00;
            reg_file[30133] <= 8'h00;
            reg_file[30134] <= 8'h00;
            reg_file[30135] <= 8'h00;
            reg_file[30136] <= 8'h00;
            reg_file[30137] <= 8'h00;
            reg_file[30138] <= 8'h00;
            reg_file[30139] <= 8'h00;
            reg_file[30140] <= 8'h00;
            reg_file[30141] <= 8'h00;
            reg_file[30142] <= 8'h00;
            reg_file[30143] <= 8'h00;
            reg_file[30144] <= 8'h00;
            reg_file[30145] <= 8'h00;
            reg_file[30146] <= 8'h00;
            reg_file[30147] <= 8'h00;
            reg_file[30148] <= 8'h00;
            reg_file[30149] <= 8'h00;
            reg_file[30150] <= 8'h00;
            reg_file[30151] <= 8'h00;
            reg_file[30152] <= 8'h00;
            reg_file[30153] <= 8'h00;
            reg_file[30154] <= 8'h00;
            reg_file[30155] <= 8'h00;
            reg_file[30156] <= 8'h00;
            reg_file[30157] <= 8'h00;
            reg_file[30158] <= 8'h00;
            reg_file[30159] <= 8'h00;
            reg_file[30160] <= 8'h00;
            reg_file[30161] <= 8'h00;
            reg_file[30162] <= 8'h00;
            reg_file[30163] <= 8'h00;
            reg_file[30164] <= 8'h00;
            reg_file[30165] <= 8'h00;
            reg_file[30166] <= 8'h00;
            reg_file[30167] <= 8'h00;
            reg_file[30168] <= 8'h00;
            reg_file[30169] <= 8'h00;
            reg_file[30170] <= 8'h00;
            reg_file[30171] <= 8'h00;
            reg_file[30172] <= 8'h00;
            reg_file[30173] <= 8'h00;
            reg_file[30174] <= 8'h00;
            reg_file[30175] <= 8'h00;
            reg_file[30176] <= 8'h00;
            reg_file[30177] <= 8'h00;
            reg_file[30178] <= 8'h00;
            reg_file[30179] <= 8'h00;
            reg_file[30180] <= 8'h00;
            reg_file[30181] <= 8'h00;
            reg_file[30182] <= 8'h00;
            reg_file[30183] <= 8'h00;
            reg_file[30184] <= 8'h00;
            reg_file[30185] <= 8'h00;
            reg_file[30186] <= 8'h00;
            reg_file[30187] <= 8'h00;
            reg_file[30188] <= 8'h00;
            reg_file[30189] <= 8'h00;
            reg_file[30190] <= 8'h00;
            reg_file[30191] <= 8'h00;
            reg_file[30192] <= 8'h00;
            reg_file[30193] <= 8'h00;
            reg_file[30194] <= 8'h00;
            reg_file[30195] <= 8'h00;
            reg_file[30196] <= 8'h00;
            reg_file[30197] <= 8'h00;
            reg_file[30198] <= 8'h00;
            reg_file[30199] <= 8'h00;
            reg_file[30200] <= 8'h00;
            reg_file[30201] <= 8'h00;
            reg_file[30202] <= 8'h00;
            reg_file[30203] <= 8'h00;
            reg_file[30204] <= 8'h00;
            reg_file[30205] <= 8'h00;
            reg_file[30206] <= 8'h00;
            reg_file[30207] <= 8'h00;
            reg_file[30208] <= 8'h00;
            reg_file[30209] <= 8'h00;
            reg_file[30210] <= 8'h00;
            reg_file[30211] <= 8'h00;
            reg_file[30212] <= 8'h00;
            reg_file[30213] <= 8'h00;
            reg_file[30214] <= 8'h00;
            reg_file[30215] <= 8'h00;
            reg_file[30216] <= 8'h00;
            reg_file[30217] <= 8'h00;
            reg_file[30218] <= 8'h00;
            reg_file[30219] <= 8'h00;
            reg_file[30220] <= 8'h00;
            reg_file[30221] <= 8'h00;
            reg_file[30222] <= 8'h00;
            reg_file[30223] <= 8'h00;
            reg_file[30224] <= 8'h00;
            reg_file[30225] <= 8'h00;
            reg_file[30226] <= 8'h00;
            reg_file[30227] <= 8'h00;
            reg_file[30228] <= 8'h00;
            reg_file[30229] <= 8'h00;
            reg_file[30230] <= 8'h00;
            reg_file[30231] <= 8'h00;
            reg_file[30232] <= 8'h00;
            reg_file[30233] <= 8'h00;
            reg_file[30234] <= 8'h00;
            reg_file[30235] <= 8'h00;
            reg_file[30236] <= 8'h00;
            reg_file[30237] <= 8'h00;
            reg_file[30238] <= 8'h00;
            reg_file[30239] <= 8'h00;
            reg_file[30240] <= 8'h00;
            reg_file[30241] <= 8'h00;
            reg_file[30242] <= 8'h00;
            reg_file[30243] <= 8'h00;
            reg_file[30244] <= 8'h00;
            reg_file[30245] <= 8'h00;
            reg_file[30246] <= 8'h00;
            reg_file[30247] <= 8'h00;
            reg_file[30248] <= 8'h00;
            reg_file[30249] <= 8'h00;
            reg_file[30250] <= 8'h00;
            reg_file[30251] <= 8'h00;
            reg_file[30252] <= 8'h00;
            reg_file[30253] <= 8'h00;
            reg_file[30254] <= 8'h00;
            reg_file[30255] <= 8'h00;
            reg_file[30256] <= 8'h00;
            reg_file[30257] <= 8'h00;
            reg_file[30258] <= 8'h00;
            reg_file[30259] <= 8'h00;
            reg_file[30260] <= 8'h00;
            reg_file[30261] <= 8'h00;
            reg_file[30262] <= 8'h00;
            reg_file[30263] <= 8'h00;
            reg_file[30264] <= 8'h00;
            reg_file[30265] <= 8'h00;
            reg_file[30266] <= 8'h00;
            reg_file[30267] <= 8'h00;
            reg_file[30268] <= 8'h00;
            reg_file[30269] <= 8'h00;
            reg_file[30270] <= 8'h00;
            reg_file[30271] <= 8'h00;
            reg_file[30272] <= 8'h00;
            reg_file[30273] <= 8'h00;
            reg_file[30274] <= 8'h00;
            reg_file[30275] <= 8'h00;
            reg_file[30276] <= 8'h00;
            reg_file[30277] <= 8'h00;
            reg_file[30278] <= 8'h00;
            reg_file[30279] <= 8'h00;
            reg_file[30280] <= 8'h00;
            reg_file[30281] <= 8'h00;
            reg_file[30282] <= 8'h00;
            reg_file[30283] <= 8'h00;
            reg_file[30284] <= 8'h00;
            reg_file[30285] <= 8'h00;
            reg_file[30286] <= 8'h00;
            reg_file[30287] <= 8'h00;
            reg_file[30288] <= 8'h00;
            reg_file[30289] <= 8'h00;
            reg_file[30290] <= 8'h00;
            reg_file[30291] <= 8'h00;
            reg_file[30292] <= 8'h00;
            reg_file[30293] <= 8'h00;
            reg_file[30294] <= 8'h00;
            reg_file[30295] <= 8'h00;
            reg_file[30296] <= 8'h00;
            reg_file[30297] <= 8'h00;
            reg_file[30298] <= 8'h00;
            reg_file[30299] <= 8'h00;
            reg_file[30300] <= 8'h00;
            reg_file[30301] <= 8'h00;
            reg_file[30302] <= 8'h00;
            reg_file[30303] <= 8'h00;
            reg_file[30304] <= 8'h00;
            reg_file[30305] <= 8'h00;
            reg_file[30306] <= 8'h00;
            reg_file[30307] <= 8'h00;
            reg_file[30308] <= 8'h00;
            reg_file[30309] <= 8'h00;
            reg_file[30310] <= 8'h00;
            reg_file[30311] <= 8'h00;
            reg_file[30312] <= 8'h00;
            reg_file[30313] <= 8'h00;
            reg_file[30314] <= 8'h00;
            reg_file[30315] <= 8'h00;
            reg_file[30316] <= 8'h00;
            reg_file[30317] <= 8'h00;
            reg_file[30318] <= 8'h00;
            reg_file[30319] <= 8'h00;
            reg_file[30320] <= 8'h00;
            reg_file[30321] <= 8'h00;
            reg_file[30322] <= 8'h00;
            reg_file[30323] <= 8'h00;
            reg_file[30324] <= 8'h00;
            reg_file[30325] <= 8'h00;
            reg_file[30326] <= 8'h00;
            reg_file[30327] <= 8'h00;
            reg_file[30328] <= 8'h00;
            reg_file[30329] <= 8'h00;
            reg_file[30330] <= 8'h00;
            reg_file[30331] <= 8'h00;
            reg_file[30332] <= 8'h00;
            reg_file[30333] <= 8'h00;
            reg_file[30334] <= 8'h00;
            reg_file[30335] <= 8'h00;
            reg_file[30336] <= 8'h00;
            reg_file[30337] <= 8'h00;
            reg_file[30338] <= 8'h00;
            reg_file[30339] <= 8'h00;
            reg_file[30340] <= 8'h00;
            reg_file[30341] <= 8'h00;
            reg_file[30342] <= 8'h00;
            reg_file[30343] <= 8'h00;
            reg_file[30344] <= 8'h00;
            reg_file[30345] <= 8'h00;
            reg_file[30346] <= 8'h00;
            reg_file[30347] <= 8'h00;
            reg_file[30348] <= 8'h00;
            reg_file[30349] <= 8'h00;
            reg_file[30350] <= 8'h00;
            reg_file[30351] <= 8'h00;
            reg_file[30352] <= 8'h00;
            reg_file[30353] <= 8'h00;
            reg_file[30354] <= 8'h00;
            reg_file[30355] <= 8'h00;
            reg_file[30356] <= 8'h00;
            reg_file[30357] <= 8'h00;
            reg_file[30358] <= 8'h00;
            reg_file[30359] <= 8'h00;
            reg_file[30360] <= 8'h00;
            reg_file[30361] <= 8'h00;
            reg_file[30362] <= 8'h00;
            reg_file[30363] <= 8'h00;
            reg_file[30364] <= 8'h00;
            reg_file[30365] <= 8'h00;
            reg_file[30366] <= 8'h00;
            reg_file[30367] <= 8'h00;
            reg_file[30368] <= 8'h00;
            reg_file[30369] <= 8'h00;
            reg_file[30370] <= 8'h00;
            reg_file[30371] <= 8'h00;
            reg_file[30372] <= 8'h00;
            reg_file[30373] <= 8'h00;
            reg_file[30374] <= 8'h00;
            reg_file[30375] <= 8'h00;
            reg_file[30376] <= 8'h00;
            reg_file[30377] <= 8'h00;
            reg_file[30378] <= 8'h00;
            reg_file[30379] <= 8'h00;
            reg_file[30380] <= 8'h00;
            reg_file[30381] <= 8'h00;
            reg_file[30382] <= 8'h00;
            reg_file[30383] <= 8'h00;
            reg_file[30384] <= 8'h00;
            reg_file[30385] <= 8'h00;
            reg_file[30386] <= 8'h00;
            reg_file[30387] <= 8'h00;
            reg_file[30388] <= 8'h00;
            reg_file[30389] <= 8'h00;
            reg_file[30390] <= 8'h00;
            reg_file[30391] <= 8'h00;
            reg_file[30392] <= 8'h00;
            reg_file[30393] <= 8'h00;
            reg_file[30394] <= 8'h00;
            reg_file[30395] <= 8'h00;
            reg_file[30396] <= 8'h00;
            reg_file[30397] <= 8'h00;
            reg_file[30398] <= 8'h00;
            reg_file[30399] <= 8'h00;
            reg_file[30400] <= 8'h00;
            reg_file[30401] <= 8'h00;
            reg_file[30402] <= 8'h00;
            reg_file[30403] <= 8'h00;
            reg_file[30404] <= 8'h00;
            reg_file[30405] <= 8'h00;
            reg_file[30406] <= 8'h00;
            reg_file[30407] <= 8'h00;
            reg_file[30408] <= 8'h00;
            reg_file[30409] <= 8'h00;
            reg_file[30410] <= 8'h00;
            reg_file[30411] <= 8'h00;
            reg_file[30412] <= 8'h00;
            reg_file[30413] <= 8'h00;
            reg_file[30414] <= 8'h00;
            reg_file[30415] <= 8'h00;
            reg_file[30416] <= 8'h00;
            reg_file[30417] <= 8'h00;
            reg_file[30418] <= 8'h00;
            reg_file[30419] <= 8'h00;
            reg_file[30420] <= 8'h00;
            reg_file[30421] <= 8'h00;
            reg_file[30422] <= 8'h00;
            reg_file[30423] <= 8'h00;
            reg_file[30424] <= 8'h00;
            reg_file[30425] <= 8'h00;
            reg_file[30426] <= 8'h00;
            reg_file[30427] <= 8'h00;
            reg_file[30428] <= 8'h00;
            reg_file[30429] <= 8'h00;
            reg_file[30430] <= 8'h00;
            reg_file[30431] <= 8'h00;
            reg_file[30432] <= 8'h00;
            reg_file[30433] <= 8'h00;
            reg_file[30434] <= 8'h00;
            reg_file[30435] <= 8'h00;
            reg_file[30436] <= 8'h00;
            reg_file[30437] <= 8'h00;
            reg_file[30438] <= 8'h00;
            reg_file[30439] <= 8'h00;
            reg_file[30440] <= 8'h00;
            reg_file[30441] <= 8'h00;
            reg_file[30442] <= 8'h00;
            reg_file[30443] <= 8'h00;
            reg_file[30444] <= 8'h00;
            reg_file[30445] <= 8'h00;
            reg_file[30446] <= 8'h00;
            reg_file[30447] <= 8'h00;
            reg_file[30448] <= 8'h00;
            reg_file[30449] <= 8'h00;
            reg_file[30450] <= 8'h00;
            reg_file[30451] <= 8'h00;
            reg_file[30452] <= 8'h00;
            reg_file[30453] <= 8'h00;
            reg_file[30454] <= 8'h00;
            reg_file[30455] <= 8'h00;
            reg_file[30456] <= 8'h00;
            reg_file[30457] <= 8'h00;
            reg_file[30458] <= 8'h00;
            reg_file[30459] <= 8'h00;
            reg_file[30460] <= 8'h00;
            reg_file[30461] <= 8'h00;
            reg_file[30462] <= 8'h00;
            reg_file[30463] <= 8'h00;
            reg_file[30464] <= 8'h00;
            reg_file[30465] <= 8'h00;
            reg_file[30466] <= 8'h00;
            reg_file[30467] <= 8'h00;
            reg_file[30468] <= 8'h00;
            reg_file[30469] <= 8'h00;
            reg_file[30470] <= 8'h00;
            reg_file[30471] <= 8'h00;
            reg_file[30472] <= 8'h00;
            reg_file[30473] <= 8'h00;
            reg_file[30474] <= 8'h00;
            reg_file[30475] <= 8'h00;
            reg_file[30476] <= 8'h00;
            reg_file[30477] <= 8'h00;
            reg_file[30478] <= 8'h00;
            reg_file[30479] <= 8'h00;
            reg_file[30480] <= 8'h00;
            reg_file[30481] <= 8'h00;
            reg_file[30482] <= 8'h00;
            reg_file[30483] <= 8'h00;
            reg_file[30484] <= 8'h00;
            reg_file[30485] <= 8'h00;
            reg_file[30486] <= 8'h00;
            reg_file[30487] <= 8'h00;
            reg_file[30488] <= 8'h00;
            reg_file[30489] <= 8'h00;
            reg_file[30490] <= 8'h00;
            reg_file[30491] <= 8'h00;
            reg_file[30492] <= 8'h00;
            reg_file[30493] <= 8'h00;
            reg_file[30494] <= 8'h00;
            reg_file[30495] <= 8'h00;
            reg_file[30496] <= 8'h00;
            reg_file[30497] <= 8'h00;
            reg_file[30498] <= 8'h00;
            reg_file[30499] <= 8'h00;
            reg_file[30500] <= 8'h00;
            reg_file[30501] <= 8'h00;
            reg_file[30502] <= 8'h00;
            reg_file[30503] <= 8'h00;
            reg_file[30504] <= 8'h00;
            reg_file[30505] <= 8'h00;
            reg_file[30506] <= 8'h00;
            reg_file[30507] <= 8'h00;
            reg_file[30508] <= 8'h00;
            reg_file[30509] <= 8'h00;
            reg_file[30510] <= 8'h00;
            reg_file[30511] <= 8'h00;
            reg_file[30512] <= 8'h00;
            reg_file[30513] <= 8'h00;
            reg_file[30514] <= 8'h00;
            reg_file[30515] <= 8'h00;
            reg_file[30516] <= 8'h00;
            reg_file[30517] <= 8'h00;
            reg_file[30518] <= 8'h00;
            reg_file[30519] <= 8'h00;
            reg_file[30520] <= 8'h00;
            reg_file[30521] <= 8'h00;
            reg_file[30522] <= 8'h00;
            reg_file[30523] <= 8'h00;
            reg_file[30524] <= 8'h00;
            reg_file[30525] <= 8'h00;
            reg_file[30526] <= 8'h00;
            reg_file[30527] <= 8'h00;
            reg_file[30528] <= 8'h00;
            reg_file[30529] <= 8'h00;
            reg_file[30530] <= 8'h00;
            reg_file[30531] <= 8'h00;
            reg_file[30532] <= 8'h00;
            reg_file[30533] <= 8'h00;
            reg_file[30534] <= 8'h00;
            reg_file[30535] <= 8'h00;
            reg_file[30536] <= 8'h00;
            reg_file[30537] <= 8'h00;
            reg_file[30538] <= 8'h00;
            reg_file[30539] <= 8'h00;
            reg_file[30540] <= 8'h00;
            reg_file[30541] <= 8'h00;
            reg_file[30542] <= 8'h00;
            reg_file[30543] <= 8'h00;
            reg_file[30544] <= 8'h00;
            reg_file[30545] <= 8'h00;
            reg_file[30546] <= 8'h00;
            reg_file[30547] <= 8'h00;
            reg_file[30548] <= 8'h00;
            reg_file[30549] <= 8'h00;
            reg_file[30550] <= 8'h00;
            reg_file[30551] <= 8'h00;
            reg_file[30552] <= 8'h00;
            reg_file[30553] <= 8'h00;
            reg_file[30554] <= 8'h00;
            reg_file[30555] <= 8'h00;
            reg_file[30556] <= 8'h00;
            reg_file[30557] <= 8'h00;
            reg_file[30558] <= 8'h00;
            reg_file[30559] <= 8'h00;
            reg_file[30560] <= 8'h00;
            reg_file[30561] <= 8'h00;
            reg_file[30562] <= 8'h00;
            reg_file[30563] <= 8'h00;
            reg_file[30564] <= 8'h00;
            reg_file[30565] <= 8'h00;
            reg_file[30566] <= 8'h00;
            reg_file[30567] <= 8'h00;
            reg_file[30568] <= 8'h00;
            reg_file[30569] <= 8'h00;
            reg_file[30570] <= 8'h00;
            reg_file[30571] <= 8'h00;
            reg_file[30572] <= 8'h00;
            reg_file[30573] <= 8'h00;
            reg_file[30574] <= 8'h00;
            reg_file[30575] <= 8'h00;
            reg_file[30576] <= 8'h00;
            reg_file[30577] <= 8'h00;
            reg_file[30578] <= 8'h00;
            reg_file[30579] <= 8'h00;
            reg_file[30580] <= 8'h00;
            reg_file[30581] <= 8'h00;
            reg_file[30582] <= 8'h00;
            reg_file[30583] <= 8'h00;
            reg_file[30584] <= 8'h00;
            reg_file[30585] <= 8'h00;
            reg_file[30586] <= 8'h00;
            reg_file[30587] <= 8'h00;
            reg_file[30588] <= 8'h00;
            reg_file[30589] <= 8'h00;
            reg_file[30590] <= 8'h00;
            reg_file[30591] <= 8'h00;
            reg_file[30592] <= 8'h00;
            reg_file[30593] <= 8'h00;
            reg_file[30594] <= 8'h00;
            reg_file[30595] <= 8'h00;
            reg_file[30596] <= 8'h00;
            reg_file[30597] <= 8'h00;
            reg_file[30598] <= 8'h00;
            reg_file[30599] <= 8'h00;
            reg_file[30600] <= 8'h00;
            reg_file[30601] <= 8'h00;
            reg_file[30602] <= 8'h00;
            reg_file[30603] <= 8'h00;
            reg_file[30604] <= 8'h00;
            reg_file[30605] <= 8'h00;
            reg_file[30606] <= 8'h00;
            reg_file[30607] <= 8'h00;
            reg_file[30608] <= 8'h00;
            reg_file[30609] <= 8'h00;
            reg_file[30610] <= 8'h00;
            reg_file[30611] <= 8'h00;
            reg_file[30612] <= 8'h00;
            reg_file[30613] <= 8'h00;
            reg_file[30614] <= 8'h00;
            reg_file[30615] <= 8'h00;
            reg_file[30616] <= 8'h00;
            reg_file[30617] <= 8'h00;
            reg_file[30618] <= 8'h00;
            reg_file[30619] <= 8'h00;
            reg_file[30620] <= 8'h00;
            reg_file[30621] <= 8'h00;
            reg_file[30622] <= 8'h00;
            reg_file[30623] <= 8'h00;
            reg_file[30624] <= 8'h00;
            reg_file[30625] <= 8'h00;
            reg_file[30626] <= 8'h00;
            reg_file[30627] <= 8'h00;
            reg_file[30628] <= 8'h00;
            reg_file[30629] <= 8'h00;
            reg_file[30630] <= 8'h00;
            reg_file[30631] <= 8'h00;
            reg_file[30632] <= 8'h00;
            reg_file[30633] <= 8'h00;
            reg_file[30634] <= 8'h00;
            reg_file[30635] <= 8'h00;
            reg_file[30636] <= 8'h00;
            reg_file[30637] <= 8'h00;
            reg_file[30638] <= 8'h00;
            reg_file[30639] <= 8'h00;
            reg_file[30640] <= 8'h00;
            reg_file[30641] <= 8'h00;
            reg_file[30642] <= 8'h00;
            reg_file[30643] <= 8'h00;
            reg_file[30644] <= 8'h00;
            reg_file[30645] <= 8'h00;
            reg_file[30646] <= 8'h00;
            reg_file[30647] <= 8'h00;
            reg_file[30648] <= 8'h00;
            reg_file[30649] <= 8'h00;
            reg_file[30650] <= 8'h00;
            reg_file[30651] <= 8'h00;
            reg_file[30652] <= 8'h00;
            reg_file[30653] <= 8'h00;
            reg_file[30654] <= 8'h00;
            reg_file[30655] <= 8'h00;
            reg_file[30656] <= 8'h00;
            reg_file[30657] <= 8'h00;
            reg_file[30658] <= 8'h00;
            reg_file[30659] <= 8'h00;
            reg_file[30660] <= 8'h00;
            reg_file[30661] <= 8'h00;
            reg_file[30662] <= 8'h00;
            reg_file[30663] <= 8'h00;
            reg_file[30664] <= 8'h00;
            reg_file[30665] <= 8'h00;
            reg_file[30666] <= 8'h00;
            reg_file[30667] <= 8'h00;
            reg_file[30668] <= 8'h00;
            reg_file[30669] <= 8'h00;
            reg_file[30670] <= 8'h00;
            reg_file[30671] <= 8'h00;
            reg_file[30672] <= 8'h00;
            reg_file[30673] <= 8'h00;
            reg_file[30674] <= 8'h00;
            reg_file[30675] <= 8'h00;
            reg_file[30676] <= 8'h00;
            reg_file[30677] <= 8'h00;
            reg_file[30678] <= 8'h00;
            reg_file[30679] <= 8'h00;
            reg_file[30680] <= 8'h00;
            reg_file[30681] <= 8'h00;
            reg_file[30682] <= 8'h00;
            reg_file[30683] <= 8'h00;
            reg_file[30684] <= 8'h00;
            reg_file[30685] <= 8'h00;
            reg_file[30686] <= 8'h00;
            reg_file[30687] <= 8'h00;
            reg_file[30688] <= 8'h00;
            reg_file[30689] <= 8'h00;
            reg_file[30690] <= 8'h00;
            reg_file[30691] <= 8'h00;
            reg_file[30692] <= 8'h00;
            reg_file[30693] <= 8'h00;
            reg_file[30694] <= 8'h00;
            reg_file[30695] <= 8'h00;
            reg_file[30696] <= 8'h00;
            reg_file[30697] <= 8'h00;
            reg_file[30698] <= 8'h00;
            reg_file[30699] <= 8'h00;
            reg_file[30700] <= 8'h00;
            reg_file[30701] <= 8'h00;
            reg_file[30702] <= 8'h00;
            reg_file[30703] <= 8'h00;
            reg_file[30704] <= 8'h00;
            reg_file[30705] <= 8'h00;
            reg_file[30706] <= 8'h00;
            reg_file[30707] <= 8'h00;
            reg_file[30708] <= 8'h00;
            reg_file[30709] <= 8'h00;
            reg_file[30710] <= 8'h00;
            reg_file[30711] <= 8'h00;
            reg_file[30712] <= 8'h00;
            reg_file[30713] <= 8'h00;
            reg_file[30714] <= 8'h00;
            reg_file[30715] <= 8'h00;
            reg_file[30716] <= 8'h00;
            reg_file[30717] <= 8'h00;
            reg_file[30718] <= 8'h00;
            reg_file[30719] <= 8'h00;
            reg_file[30720] <= 8'h00;
            reg_file[30721] <= 8'h00;
            reg_file[30722] <= 8'h00;
            reg_file[30723] <= 8'h00;
            reg_file[30724] <= 8'h00;
            reg_file[30725] <= 8'h00;
            reg_file[30726] <= 8'h00;
            reg_file[30727] <= 8'h00;
            reg_file[30728] <= 8'h00;
            reg_file[30729] <= 8'h00;
            reg_file[30730] <= 8'h00;
            reg_file[30731] <= 8'h00;
            reg_file[30732] <= 8'h00;
            reg_file[30733] <= 8'h00;
            reg_file[30734] <= 8'h00;
            reg_file[30735] <= 8'h00;
            reg_file[30736] <= 8'h00;
            reg_file[30737] <= 8'h00;
            reg_file[30738] <= 8'h00;
            reg_file[30739] <= 8'h00;
            reg_file[30740] <= 8'h00;
            reg_file[30741] <= 8'h00;
            reg_file[30742] <= 8'h00;
            reg_file[30743] <= 8'h00;
            reg_file[30744] <= 8'h00;
            reg_file[30745] <= 8'h00;
            reg_file[30746] <= 8'h00;
            reg_file[30747] <= 8'h00;
            reg_file[30748] <= 8'h00;
            reg_file[30749] <= 8'h00;
            reg_file[30750] <= 8'h00;
            reg_file[30751] <= 8'h00;
            reg_file[30752] <= 8'h00;
            reg_file[30753] <= 8'h00;
            reg_file[30754] <= 8'h00;
            reg_file[30755] <= 8'h00;
            reg_file[30756] <= 8'h00;
            reg_file[30757] <= 8'h00;
            reg_file[30758] <= 8'h00;
            reg_file[30759] <= 8'h00;
            reg_file[30760] <= 8'h00;
            reg_file[30761] <= 8'h00;
            reg_file[30762] <= 8'h00;
            reg_file[30763] <= 8'h00;
            reg_file[30764] <= 8'h00;
            reg_file[30765] <= 8'h00;
            reg_file[30766] <= 8'h00;
            reg_file[30767] <= 8'h00;
            reg_file[30768] <= 8'h00;
            reg_file[30769] <= 8'h00;
            reg_file[30770] <= 8'h00;
            reg_file[30771] <= 8'h00;
            reg_file[30772] <= 8'h00;
            reg_file[30773] <= 8'h00;
            reg_file[30774] <= 8'h00;
            reg_file[30775] <= 8'h00;
            reg_file[30776] <= 8'h00;
            reg_file[30777] <= 8'h00;
            reg_file[30778] <= 8'h00;
            reg_file[30779] <= 8'h00;
            reg_file[30780] <= 8'h00;
            reg_file[30781] <= 8'h00;
            reg_file[30782] <= 8'h00;
            reg_file[30783] <= 8'h00;
            reg_file[30784] <= 8'h00;
            reg_file[30785] <= 8'h00;
            reg_file[30786] <= 8'h00;
            reg_file[30787] <= 8'h00;
            reg_file[30788] <= 8'h00;
            reg_file[30789] <= 8'h00;
            reg_file[30790] <= 8'h00;
            reg_file[30791] <= 8'h00;
            reg_file[30792] <= 8'h00;
            reg_file[30793] <= 8'h00;
            reg_file[30794] <= 8'h00;
            reg_file[30795] <= 8'h00;
            reg_file[30796] <= 8'h00;
            reg_file[30797] <= 8'h00;
            reg_file[30798] <= 8'h00;
            reg_file[30799] <= 8'h00;
            reg_file[30800] <= 8'h00;
            reg_file[30801] <= 8'h00;
            reg_file[30802] <= 8'h00;
            reg_file[30803] <= 8'h00;
            reg_file[30804] <= 8'h00;
            reg_file[30805] <= 8'h00;
            reg_file[30806] <= 8'h00;
            reg_file[30807] <= 8'h00;
            reg_file[30808] <= 8'h00;
            reg_file[30809] <= 8'h00;
            reg_file[30810] <= 8'h00;
            reg_file[30811] <= 8'h00;
            reg_file[30812] <= 8'h00;
            reg_file[30813] <= 8'h00;
            reg_file[30814] <= 8'h00;
            reg_file[30815] <= 8'h00;
            reg_file[30816] <= 8'h00;
            reg_file[30817] <= 8'h00;
            reg_file[30818] <= 8'h00;
            reg_file[30819] <= 8'h00;
            reg_file[30820] <= 8'h00;
            reg_file[30821] <= 8'h00;
            reg_file[30822] <= 8'h00;
            reg_file[30823] <= 8'h00;
            reg_file[30824] <= 8'h00;
            reg_file[30825] <= 8'h00;
            reg_file[30826] <= 8'h00;
            reg_file[30827] <= 8'h00;
            reg_file[30828] <= 8'h00;
            reg_file[30829] <= 8'h00;
            reg_file[30830] <= 8'h00;
            reg_file[30831] <= 8'h00;
            reg_file[30832] <= 8'h00;
            reg_file[30833] <= 8'h00;
            reg_file[30834] <= 8'h00;
            reg_file[30835] <= 8'h00;
            reg_file[30836] <= 8'h00;
            reg_file[30837] <= 8'h00;
            reg_file[30838] <= 8'h00;
            reg_file[30839] <= 8'h00;
            reg_file[30840] <= 8'h00;
            reg_file[30841] <= 8'h00;
            reg_file[30842] <= 8'h00;
            reg_file[30843] <= 8'h00;
            reg_file[30844] <= 8'h00;
            reg_file[30845] <= 8'h00;
            reg_file[30846] <= 8'h00;
            reg_file[30847] <= 8'h00;
            reg_file[30848] <= 8'h00;
            reg_file[30849] <= 8'h00;
            reg_file[30850] <= 8'h00;
            reg_file[30851] <= 8'h00;
            reg_file[30852] <= 8'h00;
            reg_file[30853] <= 8'h00;
            reg_file[30854] <= 8'h00;
            reg_file[30855] <= 8'h00;
            reg_file[30856] <= 8'h00;
            reg_file[30857] <= 8'h00;
            reg_file[30858] <= 8'h00;
            reg_file[30859] <= 8'h00;
            reg_file[30860] <= 8'h00;
            reg_file[30861] <= 8'h00;
            reg_file[30862] <= 8'h00;
            reg_file[30863] <= 8'h00;
            reg_file[30864] <= 8'h00;
            reg_file[30865] <= 8'h00;
            reg_file[30866] <= 8'h00;
            reg_file[30867] <= 8'h00;
            reg_file[30868] <= 8'h00;
            reg_file[30869] <= 8'h00;
            reg_file[30870] <= 8'h00;
            reg_file[30871] <= 8'h00;
            reg_file[30872] <= 8'h00;
            reg_file[30873] <= 8'h00;
            reg_file[30874] <= 8'h00;
            reg_file[30875] <= 8'h00;
            reg_file[30876] <= 8'h00;
            reg_file[30877] <= 8'h00;
            reg_file[30878] <= 8'h00;
            reg_file[30879] <= 8'h00;
            reg_file[30880] <= 8'h00;
            reg_file[30881] <= 8'h00;
            reg_file[30882] <= 8'h00;
            reg_file[30883] <= 8'h00;
            reg_file[30884] <= 8'h00;
            reg_file[30885] <= 8'h00;
            reg_file[30886] <= 8'h00;
            reg_file[30887] <= 8'h00;
            reg_file[30888] <= 8'h00;
            reg_file[30889] <= 8'h00;
            reg_file[30890] <= 8'h00;
            reg_file[30891] <= 8'h00;
            reg_file[30892] <= 8'h00;
            reg_file[30893] <= 8'h00;
            reg_file[30894] <= 8'h00;
            reg_file[30895] <= 8'h00;
            reg_file[30896] <= 8'h00;
            reg_file[30897] <= 8'h00;
            reg_file[30898] <= 8'h00;
            reg_file[30899] <= 8'h00;
            reg_file[30900] <= 8'h00;
            reg_file[30901] <= 8'h00;
            reg_file[30902] <= 8'h00;
            reg_file[30903] <= 8'h00;
            reg_file[30904] <= 8'h00;
            reg_file[30905] <= 8'h00;
            reg_file[30906] <= 8'h00;
            reg_file[30907] <= 8'h00;
            reg_file[30908] <= 8'h00;
            reg_file[30909] <= 8'h00;
            reg_file[30910] <= 8'h00;
            reg_file[30911] <= 8'h00;
            reg_file[30912] <= 8'h00;
            reg_file[30913] <= 8'h00;
            reg_file[30914] <= 8'h00;
            reg_file[30915] <= 8'h00;
            reg_file[30916] <= 8'h00;
            reg_file[30917] <= 8'h00;
            reg_file[30918] <= 8'h00;
            reg_file[30919] <= 8'h00;
            reg_file[30920] <= 8'h00;
            reg_file[30921] <= 8'h00;
            reg_file[30922] <= 8'h00;
            reg_file[30923] <= 8'h00;
            reg_file[30924] <= 8'h00;
            reg_file[30925] <= 8'h00;
            reg_file[30926] <= 8'h00;
            reg_file[30927] <= 8'h00;
            reg_file[30928] <= 8'h00;
            reg_file[30929] <= 8'h00;
            reg_file[30930] <= 8'h00;
            reg_file[30931] <= 8'h00;
            reg_file[30932] <= 8'h00;
            reg_file[30933] <= 8'h00;
            reg_file[30934] <= 8'h00;
            reg_file[30935] <= 8'h00;
            reg_file[30936] <= 8'h00;
            reg_file[30937] <= 8'h00;
            reg_file[30938] <= 8'h00;
            reg_file[30939] <= 8'h00;
            reg_file[30940] <= 8'h00;
            reg_file[30941] <= 8'h00;
            reg_file[30942] <= 8'h00;
            reg_file[30943] <= 8'h00;
            reg_file[30944] <= 8'h00;
            reg_file[30945] <= 8'h00;
            reg_file[30946] <= 8'h00;
            reg_file[30947] <= 8'h00;
            reg_file[30948] <= 8'h00;
            reg_file[30949] <= 8'h00;
            reg_file[30950] <= 8'h00;
            reg_file[30951] <= 8'h00;
            reg_file[30952] <= 8'h00;
            reg_file[30953] <= 8'h00;
            reg_file[30954] <= 8'h00;
            reg_file[30955] <= 8'h00;
            reg_file[30956] <= 8'h00;
            reg_file[30957] <= 8'h00;
            reg_file[30958] <= 8'h00;
            reg_file[30959] <= 8'h00;
            reg_file[30960] <= 8'h00;
            reg_file[30961] <= 8'h00;
            reg_file[30962] <= 8'h00;
            reg_file[30963] <= 8'h00;
            reg_file[30964] <= 8'h00;
            reg_file[30965] <= 8'h00;
            reg_file[30966] <= 8'h00;
            reg_file[30967] <= 8'h00;
            reg_file[30968] <= 8'h00;
            reg_file[30969] <= 8'h00;
            reg_file[30970] <= 8'h00;
            reg_file[30971] <= 8'h00;
            reg_file[30972] <= 8'h00;
            reg_file[30973] <= 8'h00;
            reg_file[30974] <= 8'h00;
            reg_file[30975] <= 8'h00;
            reg_file[30976] <= 8'h00;
            reg_file[30977] <= 8'h00;
            reg_file[30978] <= 8'h00;
            reg_file[30979] <= 8'h00;
            reg_file[30980] <= 8'h00;
            reg_file[30981] <= 8'h00;
            reg_file[30982] <= 8'h00;
            reg_file[30983] <= 8'h00;
            reg_file[30984] <= 8'h00;
            reg_file[30985] <= 8'h00;
            reg_file[30986] <= 8'h00;
            reg_file[30987] <= 8'h00;
            reg_file[30988] <= 8'h00;
            reg_file[30989] <= 8'h00;
            reg_file[30990] <= 8'h00;
            reg_file[30991] <= 8'h00;
            reg_file[30992] <= 8'h00;
            reg_file[30993] <= 8'h00;
            reg_file[30994] <= 8'h00;
            reg_file[30995] <= 8'h00;
            reg_file[30996] <= 8'h00;
            reg_file[30997] <= 8'h00;
            reg_file[30998] <= 8'h00;
            reg_file[30999] <= 8'h00;
            reg_file[31000] <= 8'h00;
            reg_file[31001] <= 8'h00;
            reg_file[31002] <= 8'h00;
            reg_file[31003] <= 8'h00;
            reg_file[31004] <= 8'h00;
            reg_file[31005] <= 8'h00;
            reg_file[31006] <= 8'h00;
            reg_file[31007] <= 8'h00;
            reg_file[31008] <= 8'h00;
            reg_file[31009] <= 8'h00;
            reg_file[31010] <= 8'h00;
            reg_file[31011] <= 8'h00;
            reg_file[31012] <= 8'h00;
            reg_file[31013] <= 8'h00;
            reg_file[31014] <= 8'h00;
            reg_file[31015] <= 8'h00;
            reg_file[31016] <= 8'h00;
            reg_file[31017] <= 8'h00;
            reg_file[31018] <= 8'h00;
            reg_file[31019] <= 8'h00;
            reg_file[31020] <= 8'h00;
            reg_file[31021] <= 8'h00;
            reg_file[31022] <= 8'h00;
            reg_file[31023] <= 8'h00;
            reg_file[31024] <= 8'h00;
            reg_file[31025] <= 8'h00;
            reg_file[31026] <= 8'h00;
            reg_file[31027] <= 8'h00;
            reg_file[31028] <= 8'h00;
            reg_file[31029] <= 8'h00;
            reg_file[31030] <= 8'h00;
            reg_file[31031] <= 8'h00;
            reg_file[31032] <= 8'h00;
            reg_file[31033] <= 8'h00;
            reg_file[31034] <= 8'h00;
            reg_file[31035] <= 8'h00;
            reg_file[31036] <= 8'h00;
            reg_file[31037] <= 8'h00;
            reg_file[31038] <= 8'h00;
            reg_file[31039] <= 8'h00;
            reg_file[31040] <= 8'h00;
            reg_file[31041] <= 8'h00;
            reg_file[31042] <= 8'h00;
            reg_file[31043] <= 8'h00;
            reg_file[31044] <= 8'h00;
            reg_file[31045] <= 8'h00;
            reg_file[31046] <= 8'h00;
            reg_file[31047] <= 8'h00;
            reg_file[31048] <= 8'h00;
            reg_file[31049] <= 8'h00;
            reg_file[31050] <= 8'h00;
            reg_file[31051] <= 8'h00;
            reg_file[31052] <= 8'h00;
            reg_file[31053] <= 8'h00;
            reg_file[31054] <= 8'h00;
            reg_file[31055] <= 8'h00;
            reg_file[31056] <= 8'h00;
            reg_file[31057] <= 8'h00;
            reg_file[31058] <= 8'h00;
            reg_file[31059] <= 8'h00;
            reg_file[31060] <= 8'h00;
            reg_file[31061] <= 8'h00;
            reg_file[31062] <= 8'h00;
            reg_file[31063] <= 8'h00;
            reg_file[31064] <= 8'h00;
            reg_file[31065] <= 8'h00;
            reg_file[31066] <= 8'h00;
            reg_file[31067] <= 8'h00;
            reg_file[31068] <= 8'h00;
            reg_file[31069] <= 8'h00;
            reg_file[31070] <= 8'h00;
            reg_file[31071] <= 8'h00;
            reg_file[31072] <= 8'h00;
            reg_file[31073] <= 8'h00;
            reg_file[31074] <= 8'h00;
            reg_file[31075] <= 8'h00;
            reg_file[31076] <= 8'h00;
            reg_file[31077] <= 8'h00;
            reg_file[31078] <= 8'h00;
            reg_file[31079] <= 8'h00;
            reg_file[31080] <= 8'h00;
            reg_file[31081] <= 8'h00;
            reg_file[31082] <= 8'h00;
            reg_file[31083] <= 8'h00;
            reg_file[31084] <= 8'h00;
            reg_file[31085] <= 8'h00;
            reg_file[31086] <= 8'h00;
            reg_file[31087] <= 8'h00;
            reg_file[31088] <= 8'h00;
            reg_file[31089] <= 8'h00;
            reg_file[31090] <= 8'h00;
            reg_file[31091] <= 8'h00;
            reg_file[31092] <= 8'h00;
            reg_file[31093] <= 8'h00;
            reg_file[31094] <= 8'h00;
            reg_file[31095] <= 8'h00;
            reg_file[31096] <= 8'h00;
            reg_file[31097] <= 8'h00;
            reg_file[31098] <= 8'h00;
            reg_file[31099] <= 8'h00;
            reg_file[31100] <= 8'h00;
            reg_file[31101] <= 8'h00;
            reg_file[31102] <= 8'h00;
            reg_file[31103] <= 8'h00;
            reg_file[31104] <= 8'h00;
            reg_file[31105] <= 8'h00;
            reg_file[31106] <= 8'h00;
            reg_file[31107] <= 8'h00;
            reg_file[31108] <= 8'h00;
            reg_file[31109] <= 8'h00;
            reg_file[31110] <= 8'h00;
            reg_file[31111] <= 8'h00;
            reg_file[31112] <= 8'h00;
            reg_file[31113] <= 8'h00;
            reg_file[31114] <= 8'h00;
            reg_file[31115] <= 8'h00;
            reg_file[31116] <= 8'h00;
            reg_file[31117] <= 8'h00;
            reg_file[31118] <= 8'h00;
            reg_file[31119] <= 8'h00;
            reg_file[31120] <= 8'h00;
            reg_file[31121] <= 8'h00;
            reg_file[31122] <= 8'h00;
            reg_file[31123] <= 8'h00;
            reg_file[31124] <= 8'h00;
            reg_file[31125] <= 8'h00;
            reg_file[31126] <= 8'h00;
            reg_file[31127] <= 8'h00;
            reg_file[31128] <= 8'h00;
            reg_file[31129] <= 8'h00;
            reg_file[31130] <= 8'h00;
            reg_file[31131] <= 8'h00;
            reg_file[31132] <= 8'h00;
            reg_file[31133] <= 8'h00;
            reg_file[31134] <= 8'h00;
            reg_file[31135] <= 8'h00;
            reg_file[31136] <= 8'h00;
            reg_file[31137] <= 8'h00;
            reg_file[31138] <= 8'h00;
            reg_file[31139] <= 8'h00;
            reg_file[31140] <= 8'h00;
            reg_file[31141] <= 8'h00;
            reg_file[31142] <= 8'h00;
            reg_file[31143] <= 8'h00;
            reg_file[31144] <= 8'h00;
            reg_file[31145] <= 8'h00;
            reg_file[31146] <= 8'h00;
            reg_file[31147] <= 8'h00;
            reg_file[31148] <= 8'h00;
            reg_file[31149] <= 8'h00;
            reg_file[31150] <= 8'h00;
            reg_file[31151] <= 8'h00;
            reg_file[31152] <= 8'h00;
            reg_file[31153] <= 8'h00;
            reg_file[31154] <= 8'h00;
            reg_file[31155] <= 8'h00;
            reg_file[31156] <= 8'h00;
            reg_file[31157] <= 8'h00;
            reg_file[31158] <= 8'h00;
            reg_file[31159] <= 8'h00;
            reg_file[31160] <= 8'h00;
            reg_file[31161] <= 8'h00;
            reg_file[31162] <= 8'h00;
            reg_file[31163] <= 8'h00;
            reg_file[31164] <= 8'h00;
            reg_file[31165] <= 8'h00;
            reg_file[31166] <= 8'h00;
            reg_file[31167] <= 8'h00;
            reg_file[31168] <= 8'h00;
            reg_file[31169] <= 8'h00;
            reg_file[31170] <= 8'h00;
            reg_file[31171] <= 8'h00;
            reg_file[31172] <= 8'h00;
            reg_file[31173] <= 8'h00;
            reg_file[31174] <= 8'h00;
            reg_file[31175] <= 8'h00;
            reg_file[31176] <= 8'h00;
            reg_file[31177] <= 8'h00;
            reg_file[31178] <= 8'h00;
            reg_file[31179] <= 8'h00;
            reg_file[31180] <= 8'h00;
            reg_file[31181] <= 8'h00;
            reg_file[31182] <= 8'h00;
            reg_file[31183] <= 8'h00;
            reg_file[31184] <= 8'h00;
            reg_file[31185] <= 8'h00;
            reg_file[31186] <= 8'h00;
            reg_file[31187] <= 8'h00;
            reg_file[31188] <= 8'h00;
            reg_file[31189] <= 8'h00;
            reg_file[31190] <= 8'h00;
            reg_file[31191] <= 8'h00;
            reg_file[31192] <= 8'h00;
            reg_file[31193] <= 8'h00;
            reg_file[31194] <= 8'h00;
            reg_file[31195] <= 8'h00;
            reg_file[31196] <= 8'h00;
            reg_file[31197] <= 8'h00;
            reg_file[31198] <= 8'h00;
            reg_file[31199] <= 8'h00;
            reg_file[31200] <= 8'h00;
            reg_file[31201] <= 8'h00;
            reg_file[31202] <= 8'h00;
            reg_file[31203] <= 8'h00;
            reg_file[31204] <= 8'h00;
            reg_file[31205] <= 8'h00;
            reg_file[31206] <= 8'h00;
            reg_file[31207] <= 8'h00;
            reg_file[31208] <= 8'h00;
            reg_file[31209] <= 8'h00;
            reg_file[31210] <= 8'h00;
            reg_file[31211] <= 8'h00;
            reg_file[31212] <= 8'h00;
            reg_file[31213] <= 8'h00;
            reg_file[31214] <= 8'h00;
            reg_file[31215] <= 8'h00;
            reg_file[31216] <= 8'h00;
            reg_file[31217] <= 8'h00;
            reg_file[31218] <= 8'h00;
            reg_file[31219] <= 8'h00;
            reg_file[31220] <= 8'h00;
            reg_file[31221] <= 8'h00;
            reg_file[31222] <= 8'h00;
            reg_file[31223] <= 8'h00;
            reg_file[31224] <= 8'h00;
            reg_file[31225] <= 8'h00;
            reg_file[31226] <= 8'h00;
            reg_file[31227] <= 8'h00;
            reg_file[31228] <= 8'h00;
            reg_file[31229] <= 8'h00;
            reg_file[31230] <= 8'h00;
            reg_file[31231] <= 8'h00;
            reg_file[31232] <= 8'h00;
            reg_file[31233] <= 8'h00;
            reg_file[31234] <= 8'h00;
            reg_file[31235] <= 8'h00;
            reg_file[31236] <= 8'h00;
            reg_file[31237] <= 8'h00;
            reg_file[31238] <= 8'h00;
            reg_file[31239] <= 8'h00;
            reg_file[31240] <= 8'h00;
            reg_file[31241] <= 8'h00;
            reg_file[31242] <= 8'h00;
            reg_file[31243] <= 8'h00;
            reg_file[31244] <= 8'h00;
            reg_file[31245] <= 8'h00;
            reg_file[31246] <= 8'h00;
            reg_file[31247] <= 8'h00;
            reg_file[31248] <= 8'h00;
            reg_file[31249] <= 8'h00;
            reg_file[31250] <= 8'h00;
            reg_file[31251] <= 8'h00;
            reg_file[31252] <= 8'h00;
            reg_file[31253] <= 8'h00;
            reg_file[31254] <= 8'h00;
            reg_file[31255] <= 8'h00;
            reg_file[31256] <= 8'h00;
            reg_file[31257] <= 8'h00;
            reg_file[31258] <= 8'h00;
            reg_file[31259] <= 8'h00;
            reg_file[31260] <= 8'h00;
            reg_file[31261] <= 8'h00;
            reg_file[31262] <= 8'h00;
            reg_file[31263] <= 8'h00;
            reg_file[31264] <= 8'h00;
            reg_file[31265] <= 8'h00;
            reg_file[31266] <= 8'h00;
            reg_file[31267] <= 8'h00;
            reg_file[31268] <= 8'h00;
            reg_file[31269] <= 8'h00;
            reg_file[31270] <= 8'h00;
            reg_file[31271] <= 8'h00;
            reg_file[31272] <= 8'h00;
            reg_file[31273] <= 8'h00;
            reg_file[31274] <= 8'h00;
            reg_file[31275] <= 8'h00;
            reg_file[31276] <= 8'h00;
            reg_file[31277] <= 8'h00;
            reg_file[31278] <= 8'h00;
            reg_file[31279] <= 8'h00;
            reg_file[31280] <= 8'h00;
            reg_file[31281] <= 8'h00;
            reg_file[31282] <= 8'h00;
            reg_file[31283] <= 8'h00;
            reg_file[31284] <= 8'h00;
            reg_file[31285] <= 8'h00;
            reg_file[31286] <= 8'h00;
            reg_file[31287] <= 8'h00;
            reg_file[31288] <= 8'h00;
            reg_file[31289] <= 8'h00;
            reg_file[31290] <= 8'h00;
            reg_file[31291] <= 8'h00;
            reg_file[31292] <= 8'h00;
            reg_file[31293] <= 8'h00;
            reg_file[31294] <= 8'h00;
            reg_file[31295] <= 8'h00;
            reg_file[31296] <= 8'h00;
            reg_file[31297] <= 8'h00;
            reg_file[31298] <= 8'h00;
            reg_file[31299] <= 8'h00;
            reg_file[31300] <= 8'h00;
            reg_file[31301] <= 8'h00;
            reg_file[31302] <= 8'h00;
            reg_file[31303] <= 8'h00;
            reg_file[31304] <= 8'h00;
            reg_file[31305] <= 8'h00;
            reg_file[31306] <= 8'h00;
            reg_file[31307] <= 8'h00;
            reg_file[31308] <= 8'h00;
            reg_file[31309] <= 8'h00;
            reg_file[31310] <= 8'h00;
            reg_file[31311] <= 8'h00;
            reg_file[31312] <= 8'h00;
            reg_file[31313] <= 8'h00;
            reg_file[31314] <= 8'h00;
            reg_file[31315] <= 8'h00;
            reg_file[31316] <= 8'h00;
            reg_file[31317] <= 8'h00;
            reg_file[31318] <= 8'h00;
            reg_file[31319] <= 8'h00;
            reg_file[31320] <= 8'h00;
            reg_file[31321] <= 8'h00;
            reg_file[31322] <= 8'h00;
            reg_file[31323] <= 8'h00;
            reg_file[31324] <= 8'h00;
            reg_file[31325] <= 8'h00;
            reg_file[31326] <= 8'h00;
            reg_file[31327] <= 8'h00;
            reg_file[31328] <= 8'h00;
            reg_file[31329] <= 8'h00;
            reg_file[31330] <= 8'h00;
            reg_file[31331] <= 8'h00;
            reg_file[31332] <= 8'h00;
            reg_file[31333] <= 8'h00;
            reg_file[31334] <= 8'h00;
            reg_file[31335] <= 8'h00;
            reg_file[31336] <= 8'h00;
            reg_file[31337] <= 8'h00;
            reg_file[31338] <= 8'h00;
            reg_file[31339] <= 8'h00;
            reg_file[31340] <= 8'h00;
            reg_file[31341] <= 8'h00;
            reg_file[31342] <= 8'h00;
            reg_file[31343] <= 8'h00;
            reg_file[31344] <= 8'h00;
            reg_file[31345] <= 8'h00;
            reg_file[31346] <= 8'h00;
            reg_file[31347] <= 8'h00;
            reg_file[31348] <= 8'h00;
            reg_file[31349] <= 8'h00;
            reg_file[31350] <= 8'h00;
            reg_file[31351] <= 8'h00;
            reg_file[31352] <= 8'h00;
            reg_file[31353] <= 8'h00;
            reg_file[31354] <= 8'h00;
            reg_file[31355] <= 8'h00;
            reg_file[31356] <= 8'h00;
            reg_file[31357] <= 8'h00;
            reg_file[31358] <= 8'h00;
            reg_file[31359] <= 8'h00;
            reg_file[31360] <= 8'h00;
            reg_file[31361] <= 8'h00;
            reg_file[31362] <= 8'h00;
            reg_file[31363] <= 8'h00;
            reg_file[31364] <= 8'h00;
            reg_file[31365] <= 8'h00;
            reg_file[31366] <= 8'h00;
            reg_file[31367] <= 8'h00;
            reg_file[31368] <= 8'h00;
            reg_file[31369] <= 8'h00;
            reg_file[31370] <= 8'h00;
            reg_file[31371] <= 8'h00;
            reg_file[31372] <= 8'h00;
            reg_file[31373] <= 8'h00;
            reg_file[31374] <= 8'h00;
            reg_file[31375] <= 8'h00;
            reg_file[31376] <= 8'h00;
            reg_file[31377] <= 8'h00;
            reg_file[31378] <= 8'h00;
            reg_file[31379] <= 8'h00;
            reg_file[31380] <= 8'h00;
            reg_file[31381] <= 8'h00;
            reg_file[31382] <= 8'h00;
            reg_file[31383] <= 8'h00;
            reg_file[31384] <= 8'h00;
            reg_file[31385] <= 8'h00;
            reg_file[31386] <= 8'h00;
            reg_file[31387] <= 8'h00;
            reg_file[31388] <= 8'h00;
            reg_file[31389] <= 8'h00;
            reg_file[31390] <= 8'h00;
            reg_file[31391] <= 8'h00;
            reg_file[31392] <= 8'h00;
            reg_file[31393] <= 8'h00;
            reg_file[31394] <= 8'h00;
            reg_file[31395] <= 8'h00;
            reg_file[31396] <= 8'h00;
            reg_file[31397] <= 8'h00;
            reg_file[31398] <= 8'h00;
            reg_file[31399] <= 8'h00;
            reg_file[31400] <= 8'h00;
            reg_file[31401] <= 8'h00;
            reg_file[31402] <= 8'h00;
            reg_file[31403] <= 8'h00;
            reg_file[31404] <= 8'h00;
            reg_file[31405] <= 8'h00;
            reg_file[31406] <= 8'h00;
            reg_file[31407] <= 8'h00;
            reg_file[31408] <= 8'h00;
            reg_file[31409] <= 8'h00;
            reg_file[31410] <= 8'h00;
            reg_file[31411] <= 8'h00;
            reg_file[31412] <= 8'h00;
            reg_file[31413] <= 8'h00;
            reg_file[31414] <= 8'h00;
            reg_file[31415] <= 8'h00;
            reg_file[31416] <= 8'h00;
            reg_file[31417] <= 8'h00;
            reg_file[31418] <= 8'h00;
            reg_file[31419] <= 8'h00;
            reg_file[31420] <= 8'h00;
            reg_file[31421] <= 8'h00;
            reg_file[31422] <= 8'h00;
            reg_file[31423] <= 8'h00;
            reg_file[31424] <= 8'h00;
            reg_file[31425] <= 8'h00;
            reg_file[31426] <= 8'h00;
            reg_file[31427] <= 8'h00;
            reg_file[31428] <= 8'h00;
            reg_file[31429] <= 8'h00;
            reg_file[31430] <= 8'h00;
            reg_file[31431] <= 8'h00;
            reg_file[31432] <= 8'h00;
            reg_file[31433] <= 8'h00;
            reg_file[31434] <= 8'h00;
            reg_file[31435] <= 8'h00;
            reg_file[31436] <= 8'h00;
            reg_file[31437] <= 8'h00;
            reg_file[31438] <= 8'h00;
            reg_file[31439] <= 8'h00;
            reg_file[31440] <= 8'h00;
            reg_file[31441] <= 8'h00;
            reg_file[31442] <= 8'h00;
            reg_file[31443] <= 8'h00;
            reg_file[31444] <= 8'h00;
            reg_file[31445] <= 8'h00;
            reg_file[31446] <= 8'h00;
            reg_file[31447] <= 8'h00;
            reg_file[31448] <= 8'h00;
            reg_file[31449] <= 8'h00;
            reg_file[31450] <= 8'h00;
            reg_file[31451] <= 8'h00;
            reg_file[31452] <= 8'h00;
            reg_file[31453] <= 8'h00;
            reg_file[31454] <= 8'h00;
            reg_file[31455] <= 8'h00;
            reg_file[31456] <= 8'h00;
            reg_file[31457] <= 8'h00;
            reg_file[31458] <= 8'h00;
            reg_file[31459] <= 8'h00;
            reg_file[31460] <= 8'h00;
            reg_file[31461] <= 8'h00;
            reg_file[31462] <= 8'h00;
            reg_file[31463] <= 8'h00;
            reg_file[31464] <= 8'h00;
            reg_file[31465] <= 8'h00;
            reg_file[31466] <= 8'h00;
            reg_file[31467] <= 8'h00;
            reg_file[31468] <= 8'h00;
            reg_file[31469] <= 8'h00;
            reg_file[31470] <= 8'h00;
            reg_file[31471] <= 8'h00;
            reg_file[31472] <= 8'h00;
            reg_file[31473] <= 8'h00;
            reg_file[31474] <= 8'h00;
            reg_file[31475] <= 8'h00;
            reg_file[31476] <= 8'h00;
            reg_file[31477] <= 8'h00;
            reg_file[31478] <= 8'h00;
            reg_file[31479] <= 8'h00;
            reg_file[31480] <= 8'h00;
            reg_file[31481] <= 8'h00;
            reg_file[31482] <= 8'h00;
            reg_file[31483] <= 8'h00;
            reg_file[31484] <= 8'h00;
            reg_file[31485] <= 8'h00;
            reg_file[31486] <= 8'h00;
            reg_file[31487] <= 8'h00;
            reg_file[31488] <= 8'h00;
            reg_file[31489] <= 8'h00;
            reg_file[31490] <= 8'h00;
            reg_file[31491] <= 8'h00;
            reg_file[31492] <= 8'h00;
            reg_file[31493] <= 8'h00;
            reg_file[31494] <= 8'h00;
            reg_file[31495] <= 8'h00;
            reg_file[31496] <= 8'h00;
            reg_file[31497] <= 8'h00;
            reg_file[31498] <= 8'h00;
            reg_file[31499] <= 8'h00;
            reg_file[31500] <= 8'h00;
            reg_file[31501] <= 8'h00;
            reg_file[31502] <= 8'h00;
            reg_file[31503] <= 8'h00;
            reg_file[31504] <= 8'h00;
            reg_file[31505] <= 8'h00;
            reg_file[31506] <= 8'h00;
            reg_file[31507] <= 8'h00;
            reg_file[31508] <= 8'h00;
            reg_file[31509] <= 8'h00;
            reg_file[31510] <= 8'h00;
            reg_file[31511] <= 8'h00;
            reg_file[31512] <= 8'h00;
            reg_file[31513] <= 8'h00;
            reg_file[31514] <= 8'h00;
            reg_file[31515] <= 8'h00;
            reg_file[31516] <= 8'h00;
            reg_file[31517] <= 8'h00;
            reg_file[31518] <= 8'h00;
            reg_file[31519] <= 8'h00;
            reg_file[31520] <= 8'h00;
            reg_file[31521] <= 8'h00;
            reg_file[31522] <= 8'h00;
            reg_file[31523] <= 8'h00;
            reg_file[31524] <= 8'h00;
            reg_file[31525] <= 8'h00;
            reg_file[31526] <= 8'h00;
            reg_file[31527] <= 8'h00;
            reg_file[31528] <= 8'h00;
            reg_file[31529] <= 8'h00;
            reg_file[31530] <= 8'h00;
            reg_file[31531] <= 8'h00;
            reg_file[31532] <= 8'h00;
            reg_file[31533] <= 8'h00;
            reg_file[31534] <= 8'h00;
            reg_file[31535] <= 8'h00;
            reg_file[31536] <= 8'h00;
            reg_file[31537] <= 8'h00;
            reg_file[31538] <= 8'h00;
            reg_file[31539] <= 8'h00;
            reg_file[31540] <= 8'h00;
            reg_file[31541] <= 8'h00;
            reg_file[31542] <= 8'h00;
            reg_file[31543] <= 8'h00;
            reg_file[31544] <= 8'h00;
            reg_file[31545] <= 8'h00;
            reg_file[31546] <= 8'h00;
            reg_file[31547] <= 8'h00;
            reg_file[31548] <= 8'h00;
            reg_file[31549] <= 8'h00;
            reg_file[31550] <= 8'h00;
            reg_file[31551] <= 8'h00;
            reg_file[31552] <= 8'h00;
            reg_file[31553] <= 8'h00;
            reg_file[31554] <= 8'h00;
            reg_file[31555] <= 8'h00;
            reg_file[31556] <= 8'h00;
            reg_file[31557] <= 8'h00;
            reg_file[31558] <= 8'h00;
            reg_file[31559] <= 8'h00;
            reg_file[31560] <= 8'h00;
            reg_file[31561] <= 8'h00;
            reg_file[31562] <= 8'h00;
            reg_file[31563] <= 8'h00;
            reg_file[31564] <= 8'h00;
            reg_file[31565] <= 8'h00;
            reg_file[31566] <= 8'h00;
            reg_file[31567] <= 8'h00;
            reg_file[31568] <= 8'h00;
            reg_file[31569] <= 8'h00;
            reg_file[31570] <= 8'h00;
            reg_file[31571] <= 8'h00;
            reg_file[31572] <= 8'h00;
            reg_file[31573] <= 8'h00;
            reg_file[31574] <= 8'h00;
            reg_file[31575] <= 8'h00;
            reg_file[31576] <= 8'h00;
            reg_file[31577] <= 8'h00;
            reg_file[31578] <= 8'h00;
            reg_file[31579] <= 8'h00;
            reg_file[31580] <= 8'h00;
            reg_file[31581] <= 8'h00;
            reg_file[31582] <= 8'h00;
            reg_file[31583] <= 8'h00;
            reg_file[31584] <= 8'h00;
            reg_file[31585] <= 8'h00;
            reg_file[31586] <= 8'h00;
            reg_file[31587] <= 8'h00;
            reg_file[31588] <= 8'h00;
            reg_file[31589] <= 8'h00;
            reg_file[31590] <= 8'h00;
            reg_file[31591] <= 8'h00;
            reg_file[31592] <= 8'h00;
            reg_file[31593] <= 8'h00;
            reg_file[31594] <= 8'h00;
            reg_file[31595] <= 8'h00;
            reg_file[31596] <= 8'h00;
            reg_file[31597] <= 8'h00;
            reg_file[31598] <= 8'h00;
            reg_file[31599] <= 8'h00;
            reg_file[31600] <= 8'h00;
            reg_file[31601] <= 8'h00;
            reg_file[31602] <= 8'h00;
            reg_file[31603] <= 8'h00;
            reg_file[31604] <= 8'h00;
            reg_file[31605] <= 8'h00;
            reg_file[31606] <= 8'h00;
            reg_file[31607] <= 8'h00;
            reg_file[31608] <= 8'h00;
            reg_file[31609] <= 8'h00;
            reg_file[31610] <= 8'h00;
            reg_file[31611] <= 8'h00;
            reg_file[31612] <= 8'h00;
            reg_file[31613] <= 8'h00;
            reg_file[31614] <= 8'h00;
            reg_file[31615] <= 8'h00;
            reg_file[31616] <= 8'h00;
            reg_file[31617] <= 8'h00;
            reg_file[31618] <= 8'h00;
            reg_file[31619] <= 8'h00;
            reg_file[31620] <= 8'h00;
            reg_file[31621] <= 8'h00;
            reg_file[31622] <= 8'h00;
            reg_file[31623] <= 8'h00;
            reg_file[31624] <= 8'h00;
            reg_file[31625] <= 8'h00;
            reg_file[31626] <= 8'h00;
            reg_file[31627] <= 8'h00;
            reg_file[31628] <= 8'h00;
            reg_file[31629] <= 8'h00;
            reg_file[31630] <= 8'h00;
            reg_file[31631] <= 8'h00;
            reg_file[31632] <= 8'h00;
            reg_file[31633] <= 8'h00;
            reg_file[31634] <= 8'h00;
            reg_file[31635] <= 8'h00;
            reg_file[31636] <= 8'h00;
            reg_file[31637] <= 8'h00;
            reg_file[31638] <= 8'h00;
            reg_file[31639] <= 8'h00;
            reg_file[31640] <= 8'h00;
            reg_file[31641] <= 8'h00;
            reg_file[31642] <= 8'h00;
            reg_file[31643] <= 8'h00;
            reg_file[31644] <= 8'h00;
            reg_file[31645] <= 8'h00;
            reg_file[31646] <= 8'h00;
            reg_file[31647] <= 8'h00;
            reg_file[31648] <= 8'h00;
            reg_file[31649] <= 8'h00;
            reg_file[31650] <= 8'h00;
            reg_file[31651] <= 8'h00;
            reg_file[31652] <= 8'h00;
            reg_file[31653] <= 8'h00;
            reg_file[31654] <= 8'h00;
            reg_file[31655] <= 8'h00;
            reg_file[31656] <= 8'h00;
            reg_file[31657] <= 8'h00;
            reg_file[31658] <= 8'h00;
            reg_file[31659] <= 8'h00;
            reg_file[31660] <= 8'h00;
            reg_file[31661] <= 8'h00;
            reg_file[31662] <= 8'h00;
            reg_file[31663] <= 8'h00;
            reg_file[31664] <= 8'h00;
            reg_file[31665] <= 8'h00;
            reg_file[31666] <= 8'h00;
            reg_file[31667] <= 8'h00;
            reg_file[31668] <= 8'h00;
            reg_file[31669] <= 8'h00;
            reg_file[31670] <= 8'h00;
            reg_file[31671] <= 8'h00;
            reg_file[31672] <= 8'h00;
            reg_file[31673] <= 8'h00;
            reg_file[31674] <= 8'h00;
            reg_file[31675] <= 8'h00;
            reg_file[31676] <= 8'h00;
            reg_file[31677] <= 8'h00;
            reg_file[31678] <= 8'h00;
            reg_file[31679] <= 8'h00;
            reg_file[31680] <= 8'h00;
            reg_file[31681] <= 8'h00;
            reg_file[31682] <= 8'h00;
            reg_file[31683] <= 8'h00;
            reg_file[31684] <= 8'h00;
            reg_file[31685] <= 8'h00;
            reg_file[31686] <= 8'h00;
            reg_file[31687] <= 8'h00;
            reg_file[31688] <= 8'h00;
            reg_file[31689] <= 8'h00;
            reg_file[31690] <= 8'h00;
            reg_file[31691] <= 8'h00;
            reg_file[31692] <= 8'h00;
            reg_file[31693] <= 8'h00;
            reg_file[31694] <= 8'h00;
            reg_file[31695] <= 8'h00;
            reg_file[31696] <= 8'h00;
            reg_file[31697] <= 8'h00;
            reg_file[31698] <= 8'h00;
            reg_file[31699] <= 8'h00;
            reg_file[31700] <= 8'h00;
            reg_file[31701] <= 8'h00;
            reg_file[31702] <= 8'h00;
            reg_file[31703] <= 8'h00;
            reg_file[31704] <= 8'h00;
            reg_file[31705] <= 8'h00;
            reg_file[31706] <= 8'h00;
            reg_file[31707] <= 8'h00;
            reg_file[31708] <= 8'h00;
            reg_file[31709] <= 8'h00;
            reg_file[31710] <= 8'h00;
            reg_file[31711] <= 8'h00;
            reg_file[31712] <= 8'h00;
            reg_file[31713] <= 8'h00;
            reg_file[31714] <= 8'h00;
            reg_file[31715] <= 8'h00;
            reg_file[31716] <= 8'h00;
            reg_file[31717] <= 8'h00;
            reg_file[31718] <= 8'h00;
            reg_file[31719] <= 8'h00;
            reg_file[31720] <= 8'h00;
            reg_file[31721] <= 8'h00;
            reg_file[31722] <= 8'h00;
            reg_file[31723] <= 8'h00;
            reg_file[31724] <= 8'h00;
            reg_file[31725] <= 8'h00;
            reg_file[31726] <= 8'h00;
            reg_file[31727] <= 8'h00;
            reg_file[31728] <= 8'h00;
            reg_file[31729] <= 8'h00;
            reg_file[31730] <= 8'h00;
            reg_file[31731] <= 8'h00;
            reg_file[31732] <= 8'h00;
            reg_file[31733] <= 8'h00;
            reg_file[31734] <= 8'h00;
            reg_file[31735] <= 8'h00;
            reg_file[31736] <= 8'h00;
            reg_file[31737] <= 8'h00;
            reg_file[31738] <= 8'h00;
            reg_file[31739] <= 8'h00;
            reg_file[31740] <= 8'h00;
            reg_file[31741] <= 8'h00;
            reg_file[31742] <= 8'h00;
            reg_file[31743] <= 8'h00;
            reg_file[31744] <= 8'h00;
            reg_file[31745] <= 8'h00;
            reg_file[31746] <= 8'h00;
            reg_file[31747] <= 8'h00;
            reg_file[31748] <= 8'h00;
            reg_file[31749] <= 8'h00;
            reg_file[31750] <= 8'h00;
            reg_file[31751] <= 8'h00;
            reg_file[31752] <= 8'h00;
            reg_file[31753] <= 8'h00;
            reg_file[31754] <= 8'h00;
            reg_file[31755] <= 8'h00;
            reg_file[31756] <= 8'h00;
            reg_file[31757] <= 8'h00;
            reg_file[31758] <= 8'h00;
            reg_file[31759] <= 8'h00;
            reg_file[31760] <= 8'h00;
            reg_file[31761] <= 8'h00;
            reg_file[31762] <= 8'h00;
            reg_file[31763] <= 8'h00;
            reg_file[31764] <= 8'h00;
            reg_file[31765] <= 8'h00;
            reg_file[31766] <= 8'h00;
            reg_file[31767] <= 8'h00;
            reg_file[31768] <= 8'h00;
            reg_file[31769] <= 8'h00;
            reg_file[31770] <= 8'h00;
            reg_file[31771] <= 8'h00;
            reg_file[31772] <= 8'h00;
            reg_file[31773] <= 8'h00;
            reg_file[31774] <= 8'h00;
            reg_file[31775] <= 8'h00;
            reg_file[31776] <= 8'h00;
            reg_file[31777] <= 8'h00;
            reg_file[31778] <= 8'h00;
            reg_file[31779] <= 8'h00;
            reg_file[31780] <= 8'h00;
            reg_file[31781] <= 8'h00;
            reg_file[31782] <= 8'h00;
            reg_file[31783] <= 8'h00;
            reg_file[31784] <= 8'h00;
            reg_file[31785] <= 8'h00;
            reg_file[31786] <= 8'h00;
            reg_file[31787] <= 8'h00;
            reg_file[31788] <= 8'h00;
            reg_file[31789] <= 8'h00;
            reg_file[31790] <= 8'h00;
            reg_file[31791] <= 8'h00;
            reg_file[31792] <= 8'h00;
            reg_file[31793] <= 8'h00;
            reg_file[31794] <= 8'h00;
            reg_file[31795] <= 8'h00;
            reg_file[31796] <= 8'h00;
            reg_file[31797] <= 8'h00;
            reg_file[31798] <= 8'h00;
            reg_file[31799] <= 8'h00;
            reg_file[31800] <= 8'h00;
            reg_file[31801] <= 8'h00;
            reg_file[31802] <= 8'h00;
            reg_file[31803] <= 8'h00;
            reg_file[31804] <= 8'h00;
            reg_file[31805] <= 8'h00;
            reg_file[31806] <= 8'h00;
            reg_file[31807] <= 8'h00;
            reg_file[31808] <= 8'h00;
            reg_file[31809] <= 8'h00;
            reg_file[31810] <= 8'h00;
            reg_file[31811] <= 8'h00;
            reg_file[31812] <= 8'h00;
            reg_file[31813] <= 8'h00;
            reg_file[31814] <= 8'h00;
            reg_file[31815] <= 8'h00;
            reg_file[31816] <= 8'h00;
            reg_file[31817] <= 8'h00;
            reg_file[31818] <= 8'h00;
            reg_file[31819] <= 8'h00;
            reg_file[31820] <= 8'h00;
            reg_file[31821] <= 8'h00;
            reg_file[31822] <= 8'h00;
            reg_file[31823] <= 8'h00;
            reg_file[31824] <= 8'h00;
            reg_file[31825] <= 8'h00;
            reg_file[31826] <= 8'h00;
            reg_file[31827] <= 8'h00;
            reg_file[31828] <= 8'h00;
            reg_file[31829] <= 8'h00;
            reg_file[31830] <= 8'h00;
            reg_file[31831] <= 8'h00;
            reg_file[31832] <= 8'h00;
            reg_file[31833] <= 8'h00;
            reg_file[31834] <= 8'h00;
            reg_file[31835] <= 8'h00;
            reg_file[31836] <= 8'h00;
            reg_file[31837] <= 8'h00;
            reg_file[31838] <= 8'h00;
            reg_file[31839] <= 8'h00;
            reg_file[31840] <= 8'h00;
            reg_file[31841] <= 8'h00;
            reg_file[31842] <= 8'h00;
            reg_file[31843] <= 8'h00;
            reg_file[31844] <= 8'h00;
            reg_file[31845] <= 8'h00;
            reg_file[31846] <= 8'h00;
            reg_file[31847] <= 8'h00;
            reg_file[31848] <= 8'h00;
            reg_file[31849] <= 8'h00;
            reg_file[31850] <= 8'h00;
            reg_file[31851] <= 8'h00;
            reg_file[31852] <= 8'h00;
            reg_file[31853] <= 8'h00;
            reg_file[31854] <= 8'h00;
            reg_file[31855] <= 8'h00;
            reg_file[31856] <= 8'h00;
            reg_file[31857] <= 8'h00;
            reg_file[31858] <= 8'h00;
            reg_file[31859] <= 8'h00;
            reg_file[31860] <= 8'h00;
            reg_file[31861] <= 8'h00;
            reg_file[31862] <= 8'h00;
            reg_file[31863] <= 8'h00;
            reg_file[31864] <= 8'h00;
            reg_file[31865] <= 8'h00;
            reg_file[31866] <= 8'h00;
            reg_file[31867] <= 8'h00;
            reg_file[31868] <= 8'h00;
            reg_file[31869] <= 8'h00;
            reg_file[31870] <= 8'h00;
            reg_file[31871] <= 8'h00;
            reg_file[31872] <= 8'h00;
            reg_file[31873] <= 8'h00;
            reg_file[31874] <= 8'h00;
            reg_file[31875] <= 8'h00;
            reg_file[31876] <= 8'h00;
            reg_file[31877] <= 8'h00;
            reg_file[31878] <= 8'h00;
            reg_file[31879] <= 8'h00;
            reg_file[31880] <= 8'h00;
            reg_file[31881] <= 8'h00;
            reg_file[31882] <= 8'h00;
            reg_file[31883] <= 8'h00;
            reg_file[31884] <= 8'h00;
            reg_file[31885] <= 8'h00;
            reg_file[31886] <= 8'h00;
            reg_file[31887] <= 8'h00;
            reg_file[31888] <= 8'h00;
            reg_file[31889] <= 8'h00;
            reg_file[31890] <= 8'h00;
            reg_file[31891] <= 8'h00;
            reg_file[31892] <= 8'h00;
            reg_file[31893] <= 8'h00;
            reg_file[31894] <= 8'h00;
            reg_file[31895] <= 8'h00;
            reg_file[31896] <= 8'h00;
            reg_file[31897] <= 8'h00;
            reg_file[31898] <= 8'h00;
            reg_file[31899] <= 8'h00;
            reg_file[31900] <= 8'h00;
            reg_file[31901] <= 8'h00;
            reg_file[31902] <= 8'h00;
            reg_file[31903] <= 8'h00;
            reg_file[31904] <= 8'h00;
            reg_file[31905] <= 8'h00;
            reg_file[31906] <= 8'h00;
            reg_file[31907] <= 8'h00;
            reg_file[31908] <= 8'h00;
            reg_file[31909] <= 8'h00;
            reg_file[31910] <= 8'h00;
            reg_file[31911] <= 8'h00;
            reg_file[31912] <= 8'h00;
            reg_file[31913] <= 8'h00;
            reg_file[31914] <= 8'h00;
            reg_file[31915] <= 8'h00;
            reg_file[31916] <= 8'h00;
            reg_file[31917] <= 8'h00;
            reg_file[31918] <= 8'h00;
            reg_file[31919] <= 8'h00;
            reg_file[31920] <= 8'h00;
            reg_file[31921] <= 8'h00;
            reg_file[31922] <= 8'h00;
            reg_file[31923] <= 8'h00;
            reg_file[31924] <= 8'h00;
            reg_file[31925] <= 8'h00;
            reg_file[31926] <= 8'h00;
            reg_file[31927] <= 8'h00;
            reg_file[31928] <= 8'h00;
            reg_file[31929] <= 8'h00;
            reg_file[31930] <= 8'h00;
            reg_file[31931] <= 8'h00;
            reg_file[31932] <= 8'h00;
            reg_file[31933] <= 8'h00;
            reg_file[31934] <= 8'h00;
            reg_file[31935] <= 8'h00;
            reg_file[31936] <= 8'h00;
            reg_file[31937] <= 8'h00;
            reg_file[31938] <= 8'h00;
            reg_file[31939] <= 8'h00;
            reg_file[31940] <= 8'h00;
            reg_file[31941] <= 8'h00;
            reg_file[31942] <= 8'h00;
            reg_file[31943] <= 8'h00;
            reg_file[31944] <= 8'h00;
            reg_file[31945] <= 8'h00;
            reg_file[31946] <= 8'h00;
            reg_file[31947] <= 8'h00;
            reg_file[31948] <= 8'h00;
            reg_file[31949] <= 8'h00;
            reg_file[31950] <= 8'h00;
            reg_file[31951] <= 8'h00;
            reg_file[31952] <= 8'h00;
            reg_file[31953] <= 8'h00;
            reg_file[31954] <= 8'h00;
            reg_file[31955] <= 8'h00;
            reg_file[31956] <= 8'h00;
            reg_file[31957] <= 8'h00;
            reg_file[31958] <= 8'h00;
            reg_file[31959] <= 8'h00;
            reg_file[31960] <= 8'h00;
            reg_file[31961] <= 8'h00;
            reg_file[31962] <= 8'h00;
            reg_file[31963] <= 8'h00;
            reg_file[31964] <= 8'h00;
            reg_file[31965] <= 8'h00;
            reg_file[31966] <= 8'h00;
            reg_file[31967] <= 8'h00;
            reg_file[31968] <= 8'h00;
            reg_file[31969] <= 8'h00;
            reg_file[31970] <= 8'h00;
            reg_file[31971] <= 8'h00;
            reg_file[31972] <= 8'h00;
            reg_file[31973] <= 8'h00;
            reg_file[31974] <= 8'h00;
            reg_file[31975] <= 8'h00;
            reg_file[31976] <= 8'h00;
            reg_file[31977] <= 8'h00;
            reg_file[31978] <= 8'h00;
            reg_file[31979] <= 8'h00;
            reg_file[31980] <= 8'h00;
            reg_file[31981] <= 8'h00;
            reg_file[31982] <= 8'h00;
            reg_file[31983] <= 8'h00;
            reg_file[31984] <= 8'h00;
            reg_file[31985] <= 8'h00;
            reg_file[31986] <= 8'h00;
            reg_file[31987] <= 8'h00;
            reg_file[31988] <= 8'h00;
            reg_file[31989] <= 8'h00;
            reg_file[31990] <= 8'h00;
            reg_file[31991] <= 8'h00;
            reg_file[31992] <= 8'h00;
            reg_file[31993] <= 8'h00;
            reg_file[31994] <= 8'h00;
            reg_file[31995] <= 8'h00;
            reg_file[31996] <= 8'h00;
            reg_file[31997] <= 8'h00;
            reg_file[31998] <= 8'h00;
            reg_file[31999] <= 8'h00;
            reg_file[32000] <= 8'h00;
            reg_file[32001] <= 8'h00;
            reg_file[32002] <= 8'h00;
            reg_file[32003] <= 8'h00;
            reg_file[32004] <= 8'h00;
            reg_file[32005] <= 8'h00;
            reg_file[32006] <= 8'h00;
            reg_file[32007] <= 8'h00;
            reg_file[32008] <= 8'h00;
            reg_file[32009] <= 8'h00;
            reg_file[32010] <= 8'h00;
            reg_file[32011] <= 8'h00;
            reg_file[32012] <= 8'h00;
            reg_file[32013] <= 8'h00;
            reg_file[32014] <= 8'h00;
            reg_file[32015] <= 8'h00;
            reg_file[32016] <= 8'h00;
            reg_file[32017] <= 8'h00;
            reg_file[32018] <= 8'h00;
            reg_file[32019] <= 8'h00;
            reg_file[32020] <= 8'h00;
            reg_file[32021] <= 8'h00;
            reg_file[32022] <= 8'h00;
            reg_file[32023] <= 8'h00;
            reg_file[32024] <= 8'h00;
            reg_file[32025] <= 8'h00;
            reg_file[32026] <= 8'h00;
            reg_file[32027] <= 8'h00;
            reg_file[32028] <= 8'h00;
            reg_file[32029] <= 8'h00;
            reg_file[32030] <= 8'h00;
            reg_file[32031] <= 8'h00;
            reg_file[32032] <= 8'h00;
            reg_file[32033] <= 8'h00;
            reg_file[32034] <= 8'h00;
            reg_file[32035] <= 8'h00;
            reg_file[32036] <= 8'h00;
            reg_file[32037] <= 8'h00;
            reg_file[32038] <= 8'h00;
            reg_file[32039] <= 8'h00;
            reg_file[32040] <= 8'h00;
            reg_file[32041] <= 8'h00;
            reg_file[32042] <= 8'h00;
            reg_file[32043] <= 8'h00;
            reg_file[32044] <= 8'h00;
            reg_file[32045] <= 8'h00;
            reg_file[32046] <= 8'h00;
            reg_file[32047] <= 8'h00;
            reg_file[32048] <= 8'h00;
            reg_file[32049] <= 8'h00;
            reg_file[32050] <= 8'h00;
            reg_file[32051] <= 8'h00;
            reg_file[32052] <= 8'h00;
            reg_file[32053] <= 8'h00;
            reg_file[32054] <= 8'h00;
            reg_file[32055] <= 8'h00;
            reg_file[32056] <= 8'h00;
            reg_file[32057] <= 8'h00;
            reg_file[32058] <= 8'h00;
            reg_file[32059] <= 8'h00;
            reg_file[32060] <= 8'h00;
            reg_file[32061] <= 8'h00;
            reg_file[32062] <= 8'h00;
            reg_file[32063] <= 8'h00;
            reg_file[32064] <= 8'h00;
            reg_file[32065] <= 8'h00;
            reg_file[32066] <= 8'h00;
            reg_file[32067] <= 8'h00;
            reg_file[32068] <= 8'h00;
            reg_file[32069] <= 8'h00;
            reg_file[32070] <= 8'h00;
            reg_file[32071] <= 8'h00;
            reg_file[32072] <= 8'h00;
            reg_file[32073] <= 8'h00;
            reg_file[32074] <= 8'h00;
            reg_file[32075] <= 8'h00;
            reg_file[32076] <= 8'h00;
            reg_file[32077] <= 8'h00;
            reg_file[32078] <= 8'h00;
            reg_file[32079] <= 8'h00;
            reg_file[32080] <= 8'h00;
            reg_file[32081] <= 8'h00;
            reg_file[32082] <= 8'h00;
            reg_file[32083] <= 8'h00;
            reg_file[32084] <= 8'h00;
            reg_file[32085] <= 8'h00;
            reg_file[32086] <= 8'h00;
            reg_file[32087] <= 8'h00;
            reg_file[32088] <= 8'h00;
            reg_file[32089] <= 8'h00;
            reg_file[32090] <= 8'h00;
            reg_file[32091] <= 8'h00;
            reg_file[32092] <= 8'h00;
            reg_file[32093] <= 8'h00;
            reg_file[32094] <= 8'h00;
            reg_file[32095] <= 8'h00;
            reg_file[32096] <= 8'h00;
            reg_file[32097] <= 8'h00;
            reg_file[32098] <= 8'h00;
            reg_file[32099] <= 8'h00;
            reg_file[32100] <= 8'h00;
            reg_file[32101] <= 8'h00;
            reg_file[32102] <= 8'h00;
            reg_file[32103] <= 8'h00;
            reg_file[32104] <= 8'h00;
            reg_file[32105] <= 8'h00;
            reg_file[32106] <= 8'h00;
            reg_file[32107] <= 8'h00;
            reg_file[32108] <= 8'h00;
            reg_file[32109] <= 8'h00;
            reg_file[32110] <= 8'h00;
            reg_file[32111] <= 8'h00;
            reg_file[32112] <= 8'h00;
            reg_file[32113] <= 8'h00;
            reg_file[32114] <= 8'h00;
            reg_file[32115] <= 8'h00;
            reg_file[32116] <= 8'h00;
            reg_file[32117] <= 8'h00;
            reg_file[32118] <= 8'h00;
            reg_file[32119] <= 8'h00;
            reg_file[32120] <= 8'h00;
            reg_file[32121] <= 8'h00;
            reg_file[32122] <= 8'h00;
            reg_file[32123] <= 8'h00;
            reg_file[32124] <= 8'h00;
            reg_file[32125] <= 8'h00;
            reg_file[32126] <= 8'h00;
            reg_file[32127] <= 8'h00;
            reg_file[32128] <= 8'h00;
            reg_file[32129] <= 8'h00;
            reg_file[32130] <= 8'h00;
            reg_file[32131] <= 8'h00;
            reg_file[32132] <= 8'h00;
            reg_file[32133] <= 8'h00;
            reg_file[32134] <= 8'h00;
            reg_file[32135] <= 8'h00;
            reg_file[32136] <= 8'h00;
            reg_file[32137] <= 8'h00;
            reg_file[32138] <= 8'h00;
            reg_file[32139] <= 8'h00;
            reg_file[32140] <= 8'h00;
            reg_file[32141] <= 8'h00;
            reg_file[32142] <= 8'h00;
            reg_file[32143] <= 8'h00;
            reg_file[32144] <= 8'h00;
            reg_file[32145] <= 8'h00;
            reg_file[32146] <= 8'h00;
            reg_file[32147] <= 8'h00;
            reg_file[32148] <= 8'h00;
            reg_file[32149] <= 8'h00;
            reg_file[32150] <= 8'h00;
            reg_file[32151] <= 8'h00;
            reg_file[32152] <= 8'h00;
            reg_file[32153] <= 8'h00;
            reg_file[32154] <= 8'h00;
            reg_file[32155] <= 8'h00;
            reg_file[32156] <= 8'h00;
            reg_file[32157] <= 8'h00;
            reg_file[32158] <= 8'h00;
            reg_file[32159] <= 8'h00;
            reg_file[32160] <= 8'h00;
            reg_file[32161] <= 8'h00;
            reg_file[32162] <= 8'h00;
            reg_file[32163] <= 8'h00;
            reg_file[32164] <= 8'h00;
            reg_file[32165] <= 8'h00;
            reg_file[32166] <= 8'h00;
            reg_file[32167] <= 8'h00;
            reg_file[32168] <= 8'h00;
            reg_file[32169] <= 8'h00;
            reg_file[32170] <= 8'h00;
            reg_file[32171] <= 8'h00;
            reg_file[32172] <= 8'h00;
            reg_file[32173] <= 8'h00;
            reg_file[32174] <= 8'h00;
            reg_file[32175] <= 8'h00;
            reg_file[32176] <= 8'h00;
            reg_file[32177] <= 8'h00;
            reg_file[32178] <= 8'h00;
            reg_file[32179] <= 8'h00;
            reg_file[32180] <= 8'h00;
            reg_file[32181] <= 8'h00;
            reg_file[32182] <= 8'h00;
            reg_file[32183] <= 8'h00;
            reg_file[32184] <= 8'h00;
            reg_file[32185] <= 8'h00;
            reg_file[32186] <= 8'h00;
            reg_file[32187] <= 8'h00;
            reg_file[32188] <= 8'h00;
            reg_file[32189] <= 8'h00;
            reg_file[32190] <= 8'h00;
            reg_file[32191] <= 8'h00;
            reg_file[32192] <= 8'h00;
            reg_file[32193] <= 8'h00;
            reg_file[32194] <= 8'h00;
            reg_file[32195] <= 8'h00;
            reg_file[32196] <= 8'h00;
            reg_file[32197] <= 8'h00;
            reg_file[32198] <= 8'h00;
            reg_file[32199] <= 8'h00;
            reg_file[32200] <= 8'h00;
            reg_file[32201] <= 8'h00;
            reg_file[32202] <= 8'h00;
            reg_file[32203] <= 8'h00;
            reg_file[32204] <= 8'h00;
            reg_file[32205] <= 8'h00;
            reg_file[32206] <= 8'h00;
            reg_file[32207] <= 8'h00;
            reg_file[32208] <= 8'h00;
            reg_file[32209] <= 8'h00;
            reg_file[32210] <= 8'h00;
            reg_file[32211] <= 8'h00;
            reg_file[32212] <= 8'h00;
            reg_file[32213] <= 8'h00;
            reg_file[32214] <= 8'h00;
            reg_file[32215] <= 8'h00;
            reg_file[32216] <= 8'h00;
            reg_file[32217] <= 8'h00;
            reg_file[32218] <= 8'h00;
            reg_file[32219] <= 8'h00;
            reg_file[32220] <= 8'h00;
            reg_file[32221] <= 8'h00;
            reg_file[32222] <= 8'h00;
            reg_file[32223] <= 8'h00;
            reg_file[32224] <= 8'h00;
            reg_file[32225] <= 8'h00;
            reg_file[32226] <= 8'h00;
            reg_file[32227] <= 8'h00;
            reg_file[32228] <= 8'h00;
            reg_file[32229] <= 8'h00;
            reg_file[32230] <= 8'h00;
            reg_file[32231] <= 8'h00;
            reg_file[32232] <= 8'h00;
            reg_file[32233] <= 8'h00;
            reg_file[32234] <= 8'h00;
            reg_file[32235] <= 8'h00;
            reg_file[32236] <= 8'h00;
            reg_file[32237] <= 8'h00;
            reg_file[32238] <= 8'h00;
            reg_file[32239] <= 8'h00;
            reg_file[32240] <= 8'h00;
            reg_file[32241] <= 8'h00;
            reg_file[32242] <= 8'h00;
            reg_file[32243] <= 8'h00;
            reg_file[32244] <= 8'h00;
            reg_file[32245] <= 8'h00;
            reg_file[32246] <= 8'h00;
            reg_file[32247] <= 8'h00;
            reg_file[32248] <= 8'h00;
            reg_file[32249] <= 8'h00;
            reg_file[32250] <= 8'h00;
            reg_file[32251] <= 8'h00;
            reg_file[32252] <= 8'h00;
            reg_file[32253] <= 8'h00;
            reg_file[32254] <= 8'h00;
            reg_file[32255] <= 8'h00;
            reg_file[32256] <= 8'h00;
            reg_file[32257] <= 8'h00;
            reg_file[32258] <= 8'h00;
            reg_file[32259] <= 8'h00;
            reg_file[32260] <= 8'h00;
            reg_file[32261] <= 8'h00;
            reg_file[32262] <= 8'h00;
            reg_file[32263] <= 8'h00;
            reg_file[32264] <= 8'h00;
            reg_file[32265] <= 8'h00;
            reg_file[32266] <= 8'h00;
            reg_file[32267] <= 8'h00;
            reg_file[32268] <= 8'h00;
            reg_file[32269] <= 8'h00;
            reg_file[32270] <= 8'h00;
            reg_file[32271] <= 8'h00;
            reg_file[32272] <= 8'h00;
            reg_file[32273] <= 8'h00;
            reg_file[32274] <= 8'h00;
            reg_file[32275] <= 8'h00;
            reg_file[32276] <= 8'h00;
            reg_file[32277] <= 8'h00;
            reg_file[32278] <= 8'h00;
            reg_file[32279] <= 8'h00;
            reg_file[32280] <= 8'h00;
            reg_file[32281] <= 8'h00;
            reg_file[32282] <= 8'h00;
            reg_file[32283] <= 8'h00;
            reg_file[32284] <= 8'h00;
            reg_file[32285] <= 8'h00;
            reg_file[32286] <= 8'h00;
            reg_file[32287] <= 8'h00;
            reg_file[32288] <= 8'h00;
            reg_file[32289] <= 8'h00;
            reg_file[32290] <= 8'h00;
            reg_file[32291] <= 8'h00;
            reg_file[32292] <= 8'h00;
            reg_file[32293] <= 8'h00;
            reg_file[32294] <= 8'h00;
            reg_file[32295] <= 8'h00;
            reg_file[32296] <= 8'h00;
            reg_file[32297] <= 8'h00;
            reg_file[32298] <= 8'h00;
            reg_file[32299] <= 8'h00;
            reg_file[32300] <= 8'h00;
            reg_file[32301] <= 8'h00;
            reg_file[32302] <= 8'h00;
            reg_file[32303] <= 8'h00;
            reg_file[32304] <= 8'h00;
            reg_file[32305] <= 8'h00;
            reg_file[32306] <= 8'h00;
            reg_file[32307] <= 8'h00;
            reg_file[32308] <= 8'h00;
            reg_file[32309] <= 8'h00;
            reg_file[32310] <= 8'h00;
            reg_file[32311] <= 8'h00;
            reg_file[32312] <= 8'h00;
            reg_file[32313] <= 8'h00;
            reg_file[32314] <= 8'h00;
            reg_file[32315] <= 8'h00;
            reg_file[32316] <= 8'h00;
            reg_file[32317] <= 8'h00;
            reg_file[32318] <= 8'h00;
            reg_file[32319] <= 8'h00;
            reg_file[32320] <= 8'h00;
            reg_file[32321] <= 8'h00;
            reg_file[32322] <= 8'h00;
            reg_file[32323] <= 8'h00;
            reg_file[32324] <= 8'h00;
            reg_file[32325] <= 8'h00;
            reg_file[32326] <= 8'h00;
            reg_file[32327] <= 8'h00;
            reg_file[32328] <= 8'h00;
            reg_file[32329] <= 8'h00;
            reg_file[32330] <= 8'h00;
            reg_file[32331] <= 8'h00;
            reg_file[32332] <= 8'h00;
            reg_file[32333] <= 8'h00;
            reg_file[32334] <= 8'h00;
            reg_file[32335] <= 8'h00;
            reg_file[32336] <= 8'h00;
            reg_file[32337] <= 8'h00;
            reg_file[32338] <= 8'h00;
            reg_file[32339] <= 8'h00;
            reg_file[32340] <= 8'h00;
            reg_file[32341] <= 8'h00;
            reg_file[32342] <= 8'h00;
            reg_file[32343] <= 8'h00;
            reg_file[32344] <= 8'h00;
            reg_file[32345] <= 8'h00;
            reg_file[32346] <= 8'h00;
            reg_file[32347] <= 8'h00;
            reg_file[32348] <= 8'h00;
            reg_file[32349] <= 8'h00;
            reg_file[32350] <= 8'h00;
            reg_file[32351] <= 8'h00;
            reg_file[32352] <= 8'h00;
            reg_file[32353] <= 8'h00;
            reg_file[32354] <= 8'h00;
            reg_file[32355] <= 8'h00;
            reg_file[32356] <= 8'h00;
            reg_file[32357] <= 8'h00;
            reg_file[32358] <= 8'h00;
            reg_file[32359] <= 8'h00;
            reg_file[32360] <= 8'h00;
            reg_file[32361] <= 8'h00;
            reg_file[32362] <= 8'h00;
            reg_file[32363] <= 8'h00;
            reg_file[32364] <= 8'h00;
            reg_file[32365] <= 8'h00;
            reg_file[32366] <= 8'h00;
            reg_file[32367] <= 8'h00;
            reg_file[32368] <= 8'h00;
            reg_file[32369] <= 8'h00;
            reg_file[32370] <= 8'h00;
            reg_file[32371] <= 8'h00;
            reg_file[32372] <= 8'h00;
            reg_file[32373] <= 8'h00;
            reg_file[32374] <= 8'h00;
            reg_file[32375] <= 8'h00;
            reg_file[32376] <= 8'h00;
            reg_file[32377] <= 8'h00;
            reg_file[32378] <= 8'h00;
            reg_file[32379] <= 8'h00;
            reg_file[32380] <= 8'h00;
            reg_file[32381] <= 8'h00;
            reg_file[32382] <= 8'h00;
            reg_file[32383] <= 8'h00;
            reg_file[32384] <= 8'h00;
            reg_file[32385] <= 8'h00;
            reg_file[32386] <= 8'h00;
            reg_file[32387] <= 8'h00;
            reg_file[32388] <= 8'h00;
            reg_file[32389] <= 8'h00;
            reg_file[32390] <= 8'h00;
            reg_file[32391] <= 8'h00;
            reg_file[32392] <= 8'h00;
            reg_file[32393] <= 8'h00;
            reg_file[32394] <= 8'h00;
            reg_file[32395] <= 8'h00;
            reg_file[32396] <= 8'h00;
            reg_file[32397] <= 8'h00;
            reg_file[32398] <= 8'h00;
            reg_file[32399] <= 8'h00;
            reg_file[32400] <= 8'h00;
            reg_file[32401] <= 8'h00;
            reg_file[32402] <= 8'h00;
            reg_file[32403] <= 8'h00;
            reg_file[32404] <= 8'h00;
            reg_file[32405] <= 8'h00;
            reg_file[32406] <= 8'h00;
            reg_file[32407] <= 8'h00;
            reg_file[32408] <= 8'h00;
            reg_file[32409] <= 8'h00;
            reg_file[32410] <= 8'h00;
            reg_file[32411] <= 8'h00;
            reg_file[32412] <= 8'h00;
            reg_file[32413] <= 8'h00;
            reg_file[32414] <= 8'h00;
            reg_file[32415] <= 8'h00;
            reg_file[32416] <= 8'h00;
            reg_file[32417] <= 8'h00;
            reg_file[32418] <= 8'h00;
            reg_file[32419] <= 8'h00;
            reg_file[32420] <= 8'h00;
            reg_file[32421] <= 8'h00;
            reg_file[32422] <= 8'h00;
            reg_file[32423] <= 8'h00;
            reg_file[32424] <= 8'h00;
            reg_file[32425] <= 8'h00;
            reg_file[32426] <= 8'h00;
            reg_file[32427] <= 8'h00;
            reg_file[32428] <= 8'h00;
            reg_file[32429] <= 8'h00;
            reg_file[32430] <= 8'h00;
            reg_file[32431] <= 8'h00;
            reg_file[32432] <= 8'h00;
            reg_file[32433] <= 8'h00;
            reg_file[32434] <= 8'h00;
            reg_file[32435] <= 8'h00;
            reg_file[32436] <= 8'h00;
            reg_file[32437] <= 8'h00;
            reg_file[32438] <= 8'h00;
            reg_file[32439] <= 8'h00;
            reg_file[32440] <= 8'h00;
            reg_file[32441] <= 8'h00;
            reg_file[32442] <= 8'h00;
            reg_file[32443] <= 8'h00;
            reg_file[32444] <= 8'h00;
            reg_file[32445] <= 8'h00;
            reg_file[32446] <= 8'h00;
            reg_file[32447] <= 8'h00;
            reg_file[32448] <= 8'h00;
            reg_file[32449] <= 8'h00;
            reg_file[32450] <= 8'h00;
            reg_file[32451] <= 8'h00;
            reg_file[32452] <= 8'h00;
            reg_file[32453] <= 8'h00;
            reg_file[32454] <= 8'h00;
            reg_file[32455] <= 8'h00;
            reg_file[32456] <= 8'h00;
            reg_file[32457] <= 8'h00;
            reg_file[32458] <= 8'h00;
            reg_file[32459] <= 8'h00;
            reg_file[32460] <= 8'h00;
            reg_file[32461] <= 8'h00;
            reg_file[32462] <= 8'h00;
            reg_file[32463] <= 8'h00;
            reg_file[32464] <= 8'h00;
            reg_file[32465] <= 8'h00;
            reg_file[32466] <= 8'h00;
            reg_file[32467] <= 8'h00;
            reg_file[32468] <= 8'h00;
            reg_file[32469] <= 8'h00;
            reg_file[32470] <= 8'h00;
            reg_file[32471] <= 8'h00;
            reg_file[32472] <= 8'h00;
            reg_file[32473] <= 8'h00;
            reg_file[32474] <= 8'h00;
            reg_file[32475] <= 8'h00;
            reg_file[32476] <= 8'h00;
            reg_file[32477] <= 8'h00;
            reg_file[32478] <= 8'h00;
            reg_file[32479] <= 8'h00;
            reg_file[32480] <= 8'h00;
            reg_file[32481] <= 8'h00;
            reg_file[32482] <= 8'h00;
            reg_file[32483] <= 8'h00;
            reg_file[32484] <= 8'h00;
            reg_file[32485] <= 8'h00;
            reg_file[32486] <= 8'h00;
            reg_file[32487] <= 8'h00;
            reg_file[32488] <= 8'h00;
            reg_file[32489] <= 8'h00;
            reg_file[32490] <= 8'h00;
            reg_file[32491] <= 8'h00;
            reg_file[32492] <= 8'h00;
            reg_file[32493] <= 8'h00;
            reg_file[32494] <= 8'h00;
            reg_file[32495] <= 8'h00;
            reg_file[32496] <= 8'h00;
            reg_file[32497] <= 8'h00;
            reg_file[32498] <= 8'h00;
            reg_file[32499] <= 8'h00;
            reg_file[32500] <= 8'h00;
            reg_file[32501] <= 8'h00;
            reg_file[32502] <= 8'h00;
            reg_file[32503] <= 8'h00;
            reg_file[32504] <= 8'h00;
            reg_file[32505] <= 8'h00;
            reg_file[32506] <= 8'h00;
            reg_file[32507] <= 8'h00;
            reg_file[32508] <= 8'h00;
            reg_file[32509] <= 8'h00;
            reg_file[32510] <= 8'h00;
            reg_file[32511] <= 8'h00;
            reg_file[32512] <= 8'h00;
            reg_file[32513] <= 8'h00;
            reg_file[32514] <= 8'h00;
            reg_file[32515] <= 8'h00;
            reg_file[32516] <= 8'h00;
            reg_file[32517] <= 8'h00;
            reg_file[32518] <= 8'h00;
            reg_file[32519] <= 8'h00;
            reg_file[32520] <= 8'h00;
            reg_file[32521] <= 8'h00;
            reg_file[32522] <= 8'h00;
            reg_file[32523] <= 8'h00;
            reg_file[32524] <= 8'h00;
            reg_file[32525] <= 8'h00;
            reg_file[32526] <= 8'h00;
            reg_file[32527] <= 8'h00;
            reg_file[32528] <= 8'h00;
            reg_file[32529] <= 8'h00;
            reg_file[32530] <= 8'h00;
            reg_file[32531] <= 8'h00;
            reg_file[32532] <= 8'h00;
            reg_file[32533] <= 8'h00;
            reg_file[32534] <= 8'h00;
            reg_file[32535] <= 8'h00;
            reg_file[32536] <= 8'h00;
            reg_file[32537] <= 8'h00;
            reg_file[32538] <= 8'h00;
            reg_file[32539] <= 8'h00;
            reg_file[32540] <= 8'h00;
            reg_file[32541] <= 8'h00;
            reg_file[32542] <= 8'h00;
            reg_file[32543] <= 8'h00;
            reg_file[32544] <= 8'h00;
            reg_file[32545] <= 8'h00;
            reg_file[32546] <= 8'h00;
            reg_file[32547] <= 8'h00;
            reg_file[32548] <= 8'h00;
            reg_file[32549] <= 8'h00;
            reg_file[32550] <= 8'h00;
            reg_file[32551] <= 8'h00;
            reg_file[32552] <= 8'h00;
            reg_file[32553] <= 8'h00;
            reg_file[32554] <= 8'h00;
            reg_file[32555] <= 8'h00;
            reg_file[32556] <= 8'h00;
            reg_file[32557] <= 8'h00;
            reg_file[32558] <= 8'h00;
            reg_file[32559] <= 8'h00;
            reg_file[32560] <= 8'h00;
            reg_file[32561] <= 8'h00;
            reg_file[32562] <= 8'h00;
            reg_file[32563] <= 8'h00;
            reg_file[32564] <= 8'h00;
            reg_file[32565] <= 8'h00;
            reg_file[32566] <= 8'h00;
            reg_file[32567] <= 8'h00;
            reg_file[32568] <= 8'h00;
            reg_file[32569] <= 8'h00;
            reg_file[32570] <= 8'h00;
            reg_file[32571] <= 8'h00;
            reg_file[32572] <= 8'h00;
            reg_file[32573] <= 8'h00;
            reg_file[32574] <= 8'h00;
            reg_file[32575] <= 8'h00;
            reg_file[32576] <= 8'h00;
            reg_file[32577] <= 8'h00;
            reg_file[32578] <= 8'h00;
            reg_file[32579] <= 8'h00;
            reg_file[32580] <= 8'h00;
            reg_file[32581] <= 8'h00;
            reg_file[32582] <= 8'h00;
            reg_file[32583] <= 8'h00;
            reg_file[32584] <= 8'h00;
            reg_file[32585] <= 8'h00;
            reg_file[32586] <= 8'h00;
            reg_file[32587] <= 8'h00;
            reg_file[32588] <= 8'h00;
            reg_file[32589] <= 8'h00;
            reg_file[32590] <= 8'h00;
            reg_file[32591] <= 8'h00;
            reg_file[32592] <= 8'h00;
            reg_file[32593] <= 8'h00;
            reg_file[32594] <= 8'h00;
            reg_file[32595] <= 8'h00;
            reg_file[32596] <= 8'h00;
            reg_file[32597] <= 8'h00;
            reg_file[32598] <= 8'h00;
            reg_file[32599] <= 8'h00;
            reg_file[32600] <= 8'h00;
            reg_file[32601] <= 8'h00;
            reg_file[32602] <= 8'h00;
            reg_file[32603] <= 8'h00;
            reg_file[32604] <= 8'h00;
            reg_file[32605] <= 8'h00;
            reg_file[32606] <= 8'h00;
            reg_file[32607] <= 8'h00;
            reg_file[32608] <= 8'h00;
            reg_file[32609] <= 8'h00;
            reg_file[32610] <= 8'h00;
            reg_file[32611] <= 8'h00;
            reg_file[32612] <= 8'h00;
            reg_file[32613] <= 8'h00;
            reg_file[32614] <= 8'h00;
            reg_file[32615] <= 8'h00;
            reg_file[32616] <= 8'h00;
            reg_file[32617] <= 8'h00;
            reg_file[32618] <= 8'h00;
            reg_file[32619] <= 8'h00;
            reg_file[32620] <= 8'h00;
            reg_file[32621] <= 8'h00;
            reg_file[32622] <= 8'h00;
            reg_file[32623] <= 8'h00;
            reg_file[32624] <= 8'h00;
            reg_file[32625] <= 8'h00;
            reg_file[32626] <= 8'h00;
            reg_file[32627] <= 8'h00;
            reg_file[32628] <= 8'h00;
            reg_file[32629] <= 8'h00;
            reg_file[32630] <= 8'h00;
            reg_file[32631] <= 8'h00;
            reg_file[32632] <= 8'h00;
            reg_file[32633] <= 8'h00;
            reg_file[32634] <= 8'h00;
            reg_file[32635] <= 8'h00;
            reg_file[32636] <= 8'h00;
            reg_file[32637] <= 8'h00;
            reg_file[32638] <= 8'h00;
            reg_file[32639] <= 8'h00;
            reg_file[32640] <= 8'h00;
            reg_file[32641] <= 8'h00;
            reg_file[32642] <= 8'h00;
            reg_file[32643] <= 8'h00;
            reg_file[32644] <= 8'h00;
            reg_file[32645] <= 8'h00;
            reg_file[32646] <= 8'h00;
            reg_file[32647] <= 8'h00;
            reg_file[32648] <= 8'h00;
            reg_file[32649] <= 8'h00;
            reg_file[32650] <= 8'h00;
            reg_file[32651] <= 8'h00;
            reg_file[32652] <= 8'h00;
            reg_file[32653] <= 8'h00;
            reg_file[32654] <= 8'h00;
            reg_file[32655] <= 8'h00;
            reg_file[32656] <= 8'h00;
            reg_file[32657] <= 8'h00;
            reg_file[32658] <= 8'h00;
            reg_file[32659] <= 8'h00;
            reg_file[32660] <= 8'h00;
            reg_file[32661] <= 8'h00;
            reg_file[32662] <= 8'h00;
            reg_file[32663] <= 8'h00;
            reg_file[32664] <= 8'h00;
            reg_file[32665] <= 8'h00;
            reg_file[32666] <= 8'h00;
            reg_file[32667] <= 8'h00;
            reg_file[32668] <= 8'h00;
            reg_file[32669] <= 8'h00;
            reg_file[32670] <= 8'h00;
            reg_file[32671] <= 8'h00;
            reg_file[32672] <= 8'h00;
            reg_file[32673] <= 8'h00;
            reg_file[32674] <= 8'h00;
            reg_file[32675] <= 8'h00;
            reg_file[32676] <= 8'h00;
            reg_file[32677] <= 8'h00;
            reg_file[32678] <= 8'h00;
            reg_file[32679] <= 8'h00;
            reg_file[32680] <= 8'h00;
            reg_file[32681] <= 8'h00;
            reg_file[32682] <= 8'h00;
            reg_file[32683] <= 8'h00;
            reg_file[32684] <= 8'h00;
            reg_file[32685] <= 8'h00;
            reg_file[32686] <= 8'h00;
            reg_file[32687] <= 8'h00;
            reg_file[32688] <= 8'h00;
            reg_file[32689] <= 8'h00;
            reg_file[32690] <= 8'h00;
            reg_file[32691] <= 8'h00;
            reg_file[32692] <= 8'h00;
            reg_file[32693] <= 8'h00;
            reg_file[32694] <= 8'h00;
            reg_file[32695] <= 8'h00;
            reg_file[32696] <= 8'h00;
            reg_file[32697] <= 8'h00;
            reg_file[32698] <= 8'h00;
            reg_file[32699] <= 8'h00;
            reg_file[32700] <= 8'h00;
            reg_file[32701] <= 8'h00;
            reg_file[32702] <= 8'h00;
            reg_file[32703] <= 8'h00;
            reg_file[32704] <= 8'h00;
            reg_file[32705] <= 8'h00;
            reg_file[32706] <= 8'h00;
            reg_file[32707] <= 8'h00;
            reg_file[32708] <= 8'h00;
            reg_file[32709] <= 8'h00;
            reg_file[32710] <= 8'h00;
            reg_file[32711] <= 8'h00;
            reg_file[32712] <= 8'h00;
            reg_file[32713] <= 8'h00;
            reg_file[32714] <= 8'h00;
            reg_file[32715] <= 8'h00;
            reg_file[32716] <= 8'h00;
            reg_file[32717] <= 8'h00;
            reg_file[32718] <= 8'h00;
            reg_file[32719] <= 8'h00;
            reg_file[32720] <= 8'h00;
            reg_file[32721] <= 8'h00;
            reg_file[32722] <= 8'h00;
            reg_file[32723] <= 8'h00;
            reg_file[32724] <= 8'h00;
            reg_file[32725] <= 8'h00;
            reg_file[32726] <= 8'h00;
            reg_file[32727] <= 8'h00;
            reg_file[32728] <= 8'h00;
            reg_file[32729] <= 8'h00;
            reg_file[32730] <= 8'h00;
            reg_file[32731] <= 8'h00;
            reg_file[32732] <= 8'h00;
            reg_file[32733] <= 8'h00;
            reg_file[32734] <= 8'h00;
            reg_file[32735] <= 8'h00;
            reg_file[32736] <= 8'h00;
            reg_file[32737] <= 8'h00;
            reg_file[32738] <= 8'h00;
            reg_file[32739] <= 8'h00;
            reg_file[32740] <= 8'h00;
            reg_file[32741] <= 8'h00;
            reg_file[32742] <= 8'h00;
            reg_file[32743] <= 8'h00;
            reg_file[32744] <= 8'h00;
            reg_file[32745] <= 8'h00;
            reg_file[32746] <= 8'h00;
            reg_file[32747] <= 8'h00;
            reg_file[32748] <= 8'h00;
            reg_file[32749] <= 8'h00;
            reg_file[32750] <= 8'h00;
            reg_file[32751] <= 8'h00;
            reg_file[32752] <= 8'h00;
            reg_file[32753] <= 8'h00;
            reg_file[32754] <= 8'h00;
            reg_file[32755] <= 8'h00;
            reg_file[32756] <= 8'h00;
            reg_file[32757] <= 8'h00;
            reg_file[32758] <= 8'h00;
            reg_file[32759] <= 8'h00;
            reg_file[32760] <= 8'h00;
            reg_file[32761] <= 8'h00;
            reg_file[32762] <= 8'h00;
            reg_file[32763] <= 8'h00;
            reg_file[32764] <= 8'h00;
            reg_file[32765] <= 8'h00;
            reg_file[32766] <= 8'h00;
            reg_file[32767] <= 8'h00;
        end
        else
        begin
            reg_file <= next_reg_file;
        end
    end

    // combinational logic for memory interface
    always_comb begin : OTHER_MEM_COMB_LOGIC

        //////////////////////
        // default outputs: //
        //////////////////////

        // hold mem
        next_reg_file = reg_file;

        // Vortex outputs
        // mem_rsp_data = 512'd0;   // updated for buffer
        next_mem_rsp_data = 512'd0;

        // AHB outputs
        bpif.error = 1'b0;
        bpif.request_stall = 1'b0;

        //////////////////
        // bad address: //
        //////////////////

        // Vortex bad address
        // if (mem_req_addr[25:8] != 18'b100000000000000000)
        if (mem_req_addr[32-6-1:LOCAL_MEM_SIZE-6] != VORTEX_MEM_SLAVE_AHB_BASE_ADDR[32-1:LOCAL_MEM_SIZE])
        begin
            Vortex_bad_address = 1'b1;
        end
        else
        begin
            Vortex_bad_address = 1'b0;
        end

        // AHB bad address
        // if (gbif.addr[31:14] != 18'b101100000000000000)
        // if (bpif.addr[32-1:LOCAL_MEM_SIZE] != VORTEX_LOCAL_MEM_AHB_BASE_ADDR[32-1:LOCAL_MEM_SIZE])
        // begin
        //     AHB_bad_address = 1'b1;
        //     bpif.error = 1'b1;
        // end
        // else
        // begin
        //     AHB_bad_address = 1'b0;
        //     bpif.error = 1'b0;
        // end

        /////////////////
        // read logic: //
        /////////////////

        // Vortex read logic (this part is automated by load_Vortex_mem_slave.py)
        next_mem_rsp_data[7:0] = reg_file[{mem_req_addr[7:0], 6'd0}];
        next_mem_rsp_data[15:8] = reg_file[{mem_req_addr[7:0], 6'd1}];
        next_mem_rsp_data[23:16] = reg_file[{mem_req_addr[7:0], 6'd2}];
        next_mem_rsp_data[31:24] = reg_file[{mem_req_addr[7:0], 6'd3}];
        next_mem_rsp_data[39:32] = reg_file[{mem_req_addr[7:0], 6'd4}];
        next_mem_rsp_data[47:40] = reg_file[{mem_req_addr[7:0], 6'd5}];
        next_mem_rsp_data[55:48] = reg_file[{mem_req_addr[7:0], 6'd6}];
        next_mem_rsp_data[63:56] = reg_file[{mem_req_addr[7:0], 6'd7}];
        next_mem_rsp_data[71:64] = reg_file[{mem_req_addr[7:0], 6'd8}];
        next_mem_rsp_data[79:72] = reg_file[{mem_req_addr[7:0], 6'd9}];
        next_mem_rsp_data[87:80] = reg_file[{mem_req_addr[7:0], 6'd10}];
        next_mem_rsp_data[95:88] = reg_file[{mem_req_addr[7:0], 6'd11}];
        next_mem_rsp_data[103:96] = reg_file[{mem_req_addr[7:0], 6'd12}];
        next_mem_rsp_data[111:104] = reg_file[{mem_req_addr[7:0], 6'd13}];
        next_mem_rsp_data[119:112] = reg_file[{mem_req_addr[7:0], 6'd14}];
        next_mem_rsp_data[127:120] = reg_file[{mem_req_addr[7:0], 6'd15}];
        next_mem_rsp_data[135:128] = reg_file[{mem_req_addr[7:0], 6'd16}];
        next_mem_rsp_data[143:136] = reg_file[{mem_req_addr[7:0], 6'd17}];
        next_mem_rsp_data[151:144] = reg_file[{mem_req_addr[7:0], 6'd18}];
        next_mem_rsp_data[159:152] = reg_file[{mem_req_addr[7:0], 6'd19}];
        next_mem_rsp_data[167:160] = reg_file[{mem_req_addr[7:0], 6'd20}];
        next_mem_rsp_data[175:168] = reg_file[{mem_req_addr[7:0], 6'd21}];
        next_mem_rsp_data[183:176] = reg_file[{mem_req_addr[7:0], 6'd22}];
        next_mem_rsp_data[191:184] = reg_file[{mem_req_addr[7:0], 6'd23}];
        next_mem_rsp_data[199:192] = reg_file[{mem_req_addr[7:0], 6'd24}];
        next_mem_rsp_data[207:200] = reg_file[{mem_req_addr[7:0], 6'd25}];
        next_mem_rsp_data[215:208] = reg_file[{mem_req_addr[7:0], 6'd26}];
        next_mem_rsp_data[223:216] = reg_file[{mem_req_addr[7:0], 6'd27}];
        next_mem_rsp_data[231:224] = reg_file[{mem_req_addr[7:0], 6'd28}];
        next_mem_rsp_data[239:232] = reg_file[{mem_req_addr[7:0], 6'd29}];
        next_mem_rsp_data[247:240] = reg_file[{mem_req_addr[7:0], 6'd30}];
        next_mem_rsp_data[255:248] = reg_file[{mem_req_addr[7:0], 6'd31}];
        next_mem_rsp_data[263:256] = reg_file[{mem_req_addr[7:0], 6'd32}];
        next_mem_rsp_data[271:264] = reg_file[{mem_req_addr[7:0], 6'd33}];
        next_mem_rsp_data[279:272] = reg_file[{mem_req_addr[7:0], 6'd34}];
        next_mem_rsp_data[287:280] = reg_file[{mem_req_addr[7:0], 6'd35}];
        next_mem_rsp_data[295:288] = reg_file[{mem_req_addr[7:0], 6'd36}];
        next_mem_rsp_data[303:296] = reg_file[{mem_req_addr[7:0], 6'd37}];
        next_mem_rsp_data[311:304] = reg_file[{mem_req_addr[7:0], 6'd38}];
        next_mem_rsp_data[319:312] = reg_file[{mem_req_addr[7:0], 6'd39}];
        next_mem_rsp_data[327:320] = reg_file[{mem_req_addr[7:0], 6'd40}];
        next_mem_rsp_data[335:328] = reg_file[{mem_req_addr[7:0], 6'd41}];
        next_mem_rsp_data[343:336] = reg_file[{mem_req_addr[7:0], 6'd42}];
        next_mem_rsp_data[351:344] = reg_file[{mem_req_addr[7:0], 6'd43}];
        next_mem_rsp_data[359:352] = reg_file[{mem_req_addr[7:0], 6'd44}];
        next_mem_rsp_data[367:360] = reg_file[{mem_req_addr[7:0], 6'd45}];
        next_mem_rsp_data[375:368] = reg_file[{mem_req_addr[7:0], 6'd46}];
        next_mem_rsp_data[383:376] = reg_file[{mem_req_addr[7:0], 6'd47}];
        next_mem_rsp_data[391:384] = reg_file[{mem_req_addr[7:0], 6'd48}];
        next_mem_rsp_data[399:392] = reg_file[{mem_req_addr[7:0], 6'd49}];
        next_mem_rsp_data[407:400] = reg_file[{mem_req_addr[7:0], 6'd50}];
        next_mem_rsp_data[415:408] = reg_file[{mem_req_addr[7:0], 6'd51}];
        next_mem_rsp_data[423:416] = reg_file[{mem_req_addr[7:0], 6'd52}];
        next_mem_rsp_data[431:424] = reg_file[{mem_req_addr[7:0], 6'd53}];
        next_mem_rsp_data[439:432] = reg_file[{mem_req_addr[7:0], 6'd54}];
        next_mem_rsp_data[447:440] = reg_file[{mem_req_addr[7:0], 6'd55}];
        next_mem_rsp_data[455:448] = reg_file[{mem_req_addr[7:0], 6'd56}];
        next_mem_rsp_data[463:456] = reg_file[{mem_req_addr[7:0], 6'd57}];
        next_mem_rsp_data[471:464] = reg_file[{mem_req_addr[7:0], 6'd58}];
        next_mem_rsp_data[479:472] = reg_file[{mem_req_addr[7:0], 6'd59}];
        next_mem_rsp_data[487:480] = reg_file[{mem_req_addr[7:0], 6'd60}];
        next_mem_rsp_data[495:488] = reg_file[{mem_req_addr[7:0], 6'd61}];
        next_mem_rsp_data[503:496] = reg_file[{mem_req_addr[7:0], 6'd62}];
        next_mem_rsp_data[511:504] = reg_file[{mem_req_addr[7:0], 6'd63}];

        // AHB read logic
        bpif.rdata[7:0] = reg_file[{bpif.addr[LOCAL_MEM_SIZE-1:2], 2'd0}];
        bpif.rdata[15:8] = reg_file[{bpif.addr[LOCAL_MEM_SIZE-1:2], 2'd1}];
        bpif.rdata[23:16] = reg_file[{bpif.addr[LOCAL_MEM_SIZE-1:2], 2'd2}];
        bpif.rdata[31:24] = reg_file[{bpif.addr[LOCAL_MEM_SIZE-1:2], 2'd3}];

        //////////////////////////////////////////
        // Vortex write logic (first priority): //
        //////////////////////////////////////////

        // check for valid, write, and address in range
        // if (mem_req_valid & mem_req_rw & ~Vortex_bad_address)
        if (mem_req_valid & mem_req_rw)
        begin
            // this part is automated by load_Vortex_mem_slave.py:
            if (mem_req_byteen[0]) next_reg_file[{mem_req_addr[7:0], 6'd0}] = mem_req_data[7:0];
            if (mem_req_byteen[1]) next_reg_file[{mem_req_addr[7:0], 6'd1}] = mem_req_data[15:8];
            if (mem_req_byteen[2]) next_reg_file[{mem_req_addr[7:0], 6'd2}] = mem_req_data[23:16];
            if (mem_req_byteen[3]) next_reg_file[{mem_req_addr[7:0], 6'd3}] = mem_req_data[31:24];
            if (mem_req_byteen[4]) next_reg_file[{mem_req_addr[7:0], 6'd4}] = mem_req_data[39:32];
            if (mem_req_byteen[5]) next_reg_file[{mem_req_addr[7:0], 6'd5}] = mem_req_data[47:40];
            if (mem_req_byteen[6]) next_reg_file[{mem_req_addr[7:0], 6'd6}] = mem_req_data[55:48];
            if (mem_req_byteen[7]) next_reg_file[{mem_req_addr[7:0], 6'd7}] = mem_req_data[63:56];
            if (mem_req_byteen[8]) next_reg_file[{mem_req_addr[7:0], 6'd8}] = mem_req_data[71:64];
            if (mem_req_byteen[9]) next_reg_file[{mem_req_addr[7:0], 6'd9}] = mem_req_data[79:72];
            if (mem_req_byteen[10]) next_reg_file[{mem_req_addr[7:0], 6'd10}] = mem_req_data[87:80];
            if (mem_req_byteen[11]) next_reg_file[{mem_req_addr[7:0], 6'd11}] = mem_req_data[95:88];
            if (mem_req_byteen[12]) next_reg_file[{mem_req_addr[7:0], 6'd12}] = mem_req_data[103:96];
            if (mem_req_byteen[13]) next_reg_file[{mem_req_addr[7:0], 6'd13}] = mem_req_data[111:104];
            if (mem_req_byteen[14]) next_reg_file[{mem_req_addr[7:0], 6'd14}] = mem_req_data[119:112];
            if (mem_req_byteen[15]) next_reg_file[{mem_req_addr[7:0], 6'd15}] = mem_req_data[127:120];
            if (mem_req_byteen[16]) next_reg_file[{mem_req_addr[7:0], 6'd16}] = mem_req_data[135:128];
            if (mem_req_byteen[17]) next_reg_file[{mem_req_addr[7:0], 6'd17}] = mem_req_data[143:136];
            if (mem_req_byteen[18]) next_reg_file[{mem_req_addr[7:0], 6'd18}] = mem_req_data[151:144];
            if (mem_req_byteen[19]) next_reg_file[{mem_req_addr[7:0], 6'd19}] = mem_req_data[159:152];
            if (mem_req_byteen[20]) next_reg_file[{mem_req_addr[7:0], 6'd20}] = mem_req_data[167:160];
            if (mem_req_byteen[21]) next_reg_file[{mem_req_addr[7:0], 6'd21}] = mem_req_data[175:168];
            if (mem_req_byteen[22]) next_reg_file[{mem_req_addr[7:0], 6'd22}] = mem_req_data[183:176];
            if (mem_req_byteen[23]) next_reg_file[{mem_req_addr[7:0], 6'd23}] = mem_req_data[191:184];
            if (mem_req_byteen[24]) next_reg_file[{mem_req_addr[7:0], 6'd24}] = mem_req_data[199:192];
            if (mem_req_byteen[25]) next_reg_file[{mem_req_addr[7:0], 6'd25}] = mem_req_data[207:200];
            if (mem_req_byteen[26]) next_reg_file[{mem_req_addr[7:0], 6'd26}] = mem_req_data[215:208];
            if (mem_req_byteen[27]) next_reg_file[{mem_req_addr[7:0], 6'd27}] = mem_req_data[223:216];
            if (mem_req_byteen[28]) next_reg_file[{mem_req_addr[7:0], 6'd28}] = mem_req_data[231:224];
            if (mem_req_byteen[29]) next_reg_file[{mem_req_addr[7:0], 6'd29}] = mem_req_data[239:232];
            if (mem_req_byteen[30]) next_reg_file[{mem_req_addr[7:0], 6'd30}] = mem_req_data[247:240];
            if (mem_req_byteen[31]) next_reg_file[{mem_req_addr[7:0], 6'd31}] = mem_req_data[255:248];
            if (mem_req_byteen[32]) next_reg_file[{mem_req_addr[7:0], 6'd32}] = mem_req_data[263:256];
            if (mem_req_byteen[33]) next_reg_file[{mem_req_addr[7:0], 6'd33}] = mem_req_data[271:264];
            if (mem_req_byteen[34]) next_reg_file[{mem_req_addr[7:0], 6'd34}] = mem_req_data[279:272];
            if (mem_req_byteen[35]) next_reg_file[{mem_req_addr[7:0], 6'd35}] = mem_req_data[287:280];
            if (mem_req_byteen[36]) next_reg_file[{mem_req_addr[7:0], 6'd36}] = mem_req_data[295:288];
            if (mem_req_byteen[37]) next_reg_file[{mem_req_addr[7:0], 6'd37}] = mem_req_data[303:296];
            if (mem_req_byteen[38]) next_reg_file[{mem_req_addr[7:0], 6'd38}] = mem_req_data[311:304];
            if (mem_req_byteen[39]) next_reg_file[{mem_req_addr[7:0], 6'd39}] = mem_req_data[319:312];
            if (mem_req_byteen[40]) next_reg_file[{mem_req_addr[7:0], 6'd40}] = mem_req_data[327:320];
            if (mem_req_byteen[41]) next_reg_file[{mem_req_addr[7:0], 6'd41}] = mem_req_data[335:328];
            if (mem_req_byteen[42]) next_reg_file[{mem_req_addr[7:0], 6'd42}] = mem_req_data[343:336];
            if (mem_req_byteen[43]) next_reg_file[{mem_req_addr[7:0], 6'd43}] = mem_req_data[351:344];
            if (mem_req_byteen[44]) next_reg_file[{mem_req_addr[7:0], 6'd44}] = mem_req_data[359:352];
            if (mem_req_byteen[45]) next_reg_file[{mem_req_addr[7:0], 6'd45}] = mem_req_data[367:360];
            if (mem_req_byteen[46]) next_reg_file[{mem_req_addr[7:0], 6'd46}] = mem_req_data[375:368];
            if (mem_req_byteen[47]) next_reg_file[{mem_req_addr[7:0], 6'd47}] = mem_req_data[383:376];
            if (mem_req_byteen[48]) next_reg_file[{mem_req_addr[7:0], 6'd48}] = mem_req_data[391:384];
            if (mem_req_byteen[49]) next_reg_file[{mem_req_addr[7:0], 6'd49}] = mem_req_data[399:392];
            if (mem_req_byteen[50]) next_reg_file[{mem_req_addr[7:0], 6'd50}] = mem_req_data[407:400];
            if (mem_req_byteen[51]) next_reg_file[{mem_req_addr[7:0], 6'd51}] = mem_req_data[415:408];
            if (mem_req_byteen[52]) next_reg_file[{mem_req_addr[7:0], 6'd52}] = mem_req_data[423:416];
            if (mem_req_byteen[53]) next_reg_file[{mem_req_addr[7:0], 6'd53}] = mem_req_data[431:424];
            if (mem_req_byteen[54]) next_reg_file[{mem_req_addr[7:0], 6'd54}] = mem_req_data[439:432];
            if (mem_req_byteen[55]) next_reg_file[{mem_req_addr[7:0], 6'd55}] = mem_req_data[447:440];
            if (mem_req_byteen[56]) next_reg_file[{mem_req_addr[7:0], 6'd56}] = mem_req_data[455:448];
            if (mem_req_byteen[57]) next_reg_file[{mem_req_addr[7:0], 6'd57}] = mem_req_data[463:456];
            if (mem_req_byteen[58]) next_reg_file[{mem_req_addr[7:0], 6'd58}] = mem_req_data[471:464];
            if (mem_req_byteen[59]) next_reg_file[{mem_req_addr[7:0], 6'd59}] = mem_req_data[479:472];
            if (mem_req_byteen[60]) next_reg_file[{mem_req_addr[7:0], 6'd60}] = mem_req_data[487:480];
            if (mem_req_byteen[61]) next_reg_file[{mem_req_addr[7:0], 6'd61}] = mem_req_data[495:488];
            if (mem_req_byteen[62]) next_reg_file[{mem_req_addr[7:0], 6'd62}] = mem_req_data[503:496];
            if (mem_req_byteen[63]) next_reg_file[{mem_req_addr[7:0], 6'd63}] = mem_req_data[511:504];

            // ahb busy
            bpif.request_stall = 1'b1;
        end

        ////////////////////////////////////////
        // AHB write logic (second priority): //
        ////////////////////////////////////////

        // if Vortex not writing, check for write and address in range
        // else if (bpif.wen & ~AHB_bad_address)
        else if (bpif.wen)
        begin
            // assumption: follow word address
            if (bpif.strobe[0]) next_reg_file[{bpif.addr[LOCAL_MEM_SIZE-1:2], 2'd0}] = bpif.wdata[7:0];
            if (bpif.strobe[1]) next_reg_file[{bpif.addr[LOCAL_MEM_SIZE-1:2], 2'd1}] = bpif.wdata[15:8];
            if (bpif.strobe[2]) next_reg_file[{bpif.addr[LOCAL_MEM_SIZE-1:2], 2'd2}] = bpif.wdata[23:16];
            if (bpif.strobe[3]) next_reg_file[{bpif.addr[LOCAL_MEM_SIZE-1:2], 2'd3}] = bpif.wdata[31:24];
        end

        ////////////////////////////////
        // other combinational logic: //
        ////////////////////////////////

        // always ready for request
        mem_req_ready = 1'b1;           

        // read ready immediately
        // mem_rsp_valid = mem_req_valid;   // updated for buffer
        next_mem_rsp_valid = mem_req_valid & ~mem_req_rw;   // only need to respond for reads

        // match req immediately
        // mem_rsp_tag = mem_req_tag;       // updated for buffer
        next_mem_rsp_tag = mem_req_tag;
    end

    // only status registers use Vortex busy

endmodule

