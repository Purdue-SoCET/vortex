/*
    socet115 / zlagpaca@purdue.edu
    Zach Lagpacan

    module for faking memory with basic register file which can interface with Vortex memory interface
*/

// temporary include to have defined vals
// `include "local_mem.vh"
`include "../include/VX_define.vh"
// `include "VX_define.vh"

module local_mem #(
)(
    // seq
    input clk, reset,

    // Memory Request:
    // vortex outputs
    input logic                             mem_req_valid,
    input logic                             mem_req_rw,
    input logic [`VX_MEM_BYTEEN_WIDTH-1:0]  mem_req_byteen, // 64 (512 / 8)
    input logic [`VX_MEM_ADDR_WIDTH-1:0]    mem_req_addr,   // 26
    input logic [`VX_MEM_DATA_WIDTH-1:0]    mem_req_data,   // 512
    input logic [`VX_MEM_TAG_WIDTH-1:0]     mem_req_tag,    // 56 (55 for SM disabled)
    // vortex inputs
    output logic                            mem_req_ready,

    // Memory response:
    // vortex inputs
    output logic                            mem_rsp_valid,        
    output logic [`VX_MEM_DATA_WIDTH-1:0]   mem_rsp_data,   // 512
    output logic [`VX_MEM_TAG_WIDTH-1:0]    mem_rsp_tag,    // 56 (55 for SM disabled)
    // vortex outputs
    input logic                             mem_rsp_ready,

    // Status:
    // vortex outputs
    input logic                             busy,

    // tb:
    output logic                            tb_addr_out_of_bounds
);
    // register file instances
    
    // chunk 0
    logic wen_0_80000000;
    logic [5-1:0] wsel_0_80000000;
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_0_80000000;
    logic [5-1:0] rsel_0_80000000;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_0_80000000;
    
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_0_80000000 [32-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_0_80000000 [32-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_0_80000000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_0_80000000[0][31:0] <= 32'h6F008004;
            reg_val_0_80000000[0][63:32] <= 32'h732F2034;
            reg_val_0_80000000[0][95:64] <= 32'h930F8000;
            reg_val_0_80000000[0][127:96] <= 32'h6308FF03;
            reg_val_0_80000000[0][159:128] <= 32'h930F9000;
            reg_val_0_80000000[0][191:160] <= 32'h6304FF03;
            reg_val_0_80000000[0][223:192] <= 32'h930FB000;
            reg_val_0_80000000[0][255:224] <= 32'h6300FF03;
            reg_val_0_80000000[0][287:256] <= 32'h130F0000;
            reg_val_0_80000000[0][319:288] <= 32'h63040F00;
            reg_val_0_80000000[0][351:320] <= 32'h67000F00;
            reg_val_0_80000000[0][383:352] <= 32'h732F2034;
            reg_val_0_80000000[0][415:384] <= 32'h63540F00;
            reg_val_0_80000000[0][447:416] <= 32'h6F004000;
            reg_val_0_80000000[0][479:448] <= 32'h93E19153;
            reg_val_0_80000000[0][511:480] <= 32'h171F0000;
            reg_val_0_80000000[1][31:0] <= 32'h23223FFC;
            reg_val_0_80000000[1][63:32] <= 32'h6FF09FFF;
            reg_val_0_80000000[1][95:64] <= 32'h93000000;
            reg_val_0_80000000[1][127:96] <= 32'h13010000;
            reg_val_0_80000000[1][159:128] <= 32'h93010000;
            reg_val_0_80000000[1][191:160] <= 32'h13020000;
            reg_val_0_80000000[1][223:192] <= 32'h93020000;
            reg_val_0_80000000[1][255:224] <= 32'h13030000;
            reg_val_0_80000000[1][287:256] <= 32'h93030000;
            reg_val_0_80000000[1][319:288] <= 32'h13040000;
            reg_val_0_80000000[1][351:320] <= 32'h93040000;
            reg_val_0_80000000[1][383:352] <= 32'h13050000;
            reg_val_0_80000000[1][415:384] <= 32'h93050000;
            reg_val_0_80000000[1][447:416] <= 32'h13060000;
            reg_val_0_80000000[1][479:448] <= 32'h93060000;
            reg_val_0_80000000[1][511:480] <= 32'h13070000;
            reg_val_0_80000000[2][31:0] <= 32'h93070000;
            reg_val_0_80000000[2][63:32] <= 32'h13080000;
            reg_val_0_80000000[2][95:64] <= 32'h93080000;
            reg_val_0_80000000[2][127:96] <= 32'h13090000;
            reg_val_0_80000000[2][159:128] <= 32'h93090000;
            reg_val_0_80000000[2][191:160] <= 32'h130A0000;
            reg_val_0_80000000[2][223:192] <= 32'h930A0000;
            reg_val_0_80000000[2][255:224] <= 32'h130B0000;
            reg_val_0_80000000[2][287:256] <= 32'h930B0000;
            reg_val_0_80000000[2][319:288] <= 32'h130C0000;
            reg_val_0_80000000[2][351:320] <= 32'h930C0000;
            reg_val_0_80000000[2][383:352] <= 32'h130D0000;
            reg_val_0_80000000[2][415:384] <= 32'h930D0000;
            reg_val_0_80000000[2][447:416] <= 32'h130E0000;
            reg_val_0_80000000[2][479:448] <= 32'h930E0000;
            reg_val_0_80000000[2][511:480] <= 32'h130F0000;
            reg_val_0_80000000[3][31:0] <= 32'h930F0000;
            reg_val_0_80000000[3][63:32] <= 32'h732540F1;
            reg_val_0_80000000[3][95:64] <= 32'h63100500;
            reg_val_0_80000000[3][127:96] <= 32'h97020000;
            reg_val_0_80000000[3][159:128] <= 32'h93820201;
            reg_val_0_80000000[3][191:160] <= 32'h73905230;
            reg_val_0_80000000[3][223:192] <= 32'h73500018;
            reg_val_0_80000000[3][255:224] <= 32'h97020000;
            reg_val_0_80000000[3][287:256] <= 32'h93820202;
            reg_val_0_80000000[3][319:288] <= 32'h73905230;
            reg_val_0_80000000[3][351:320] <= 32'hB7020080;
            reg_val_0_80000000[3][383:352] <= 32'h9382F2FF;
            reg_val_0_80000000[3][415:384] <= 32'h7390023B;
            reg_val_0_80000000[3][447:416] <= 32'h9302F001;
            reg_val_0_80000000[3][479:448] <= 32'h7390023A;
            reg_val_0_80000000[3][511:480] <= 32'h73504030;
            reg_val_0_80000000[4][31:0] <= 32'h97020000;
            reg_val_0_80000000[4][63:32] <= 32'h93824201;
            reg_val_0_80000000[4][95:64] <= 32'h73905230;
            reg_val_0_80000000[4][127:96] <= 32'h73502030;
            reg_val_0_80000000[4][159:128] <= 32'h73503030;
            reg_val_0_80000000[4][191:160] <= 32'h93010000;
            reg_val_0_80000000[4][223:192] <= 32'h97020000;
            reg_val_0_80000000[4][255:224] <= 32'h9382C2EE;
            reg_val_0_80000000[4][287:256] <= 32'h73905230;
            reg_val_0_80000000[4][319:288] <= 32'h13051000;
            reg_val_0_80000000[4][351:320] <= 32'h1315F501;
            reg_val_0_80000000[4][383:352] <= 32'h634C0500;
            reg_val_0_80000000[4][415:384] <= 32'h0F00F00F;
            reg_val_0_80000000[4][447:416] <= 32'h93011000;
            reg_val_0_80000000[4][479:448] <= 32'h9308D005;
            reg_val_0_80000000[4][511:480] <= 32'h13050000;
            reg_val_0_80000000[5][31:0] <= 32'h73000000;
            reg_val_0_80000000[5][63:32] <= 32'h93020000;
            reg_val_0_80000000[5][95:64] <= 32'h638A0200;
            reg_val_0_80000000[5][127:96] <= 32'h73905210;
            reg_val_0_80000000[5][159:128] <= 32'hB7B20000;
            reg_val_0_80000000[5][191:160] <= 32'h93829210;
            reg_val_0_80000000[5][223:192] <= 32'h73902230;
            reg_val_0_80000000[5][255:224] <= 32'h73500030;
            reg_val_0_80000000[5][287:256] <= 32'h37250000;
            reg_val_0_80000000[5][319:288] <= 32'h73200530;
            reg_val_0_80000000[5][351:320] <= 32'h73503000;
            reg_val_0_80000000[5][383:352] <= 32'h97020000;
            reg_val_0_80000000[5][415:384] <= 32'h93824201;
            reg_val_0_80000000[5][447:416] <= 32'h73901234;
            reg_val_0_80000000[5][479:448] <= 32'h732540F1;
            reg_val_0_80000000[5][511:480] <= 32'h73002030;
            reg_val_0_80000000[6][31:0] <= 32'h93012000;
            reg_val_0_80000000[6][63:32] <= 32'h17250000;
            reg_val_0_80000000[6][95:64] <= 32'h1305C5E7;
            reg_val_0_80000000[6][127:96] <= 32'h07300500;
            reg_val_0_80000000[6][159:128] <= 32'h87308500;
            reg_val_0_80000000[6][191:160] <= 32'h07310501;
            reg_val_0_80000000[6][223:192] <= 32'h83268501;
            reg_val_0_80000000[6][255:224] <= 32'h0323C501;
            reg_val_0_80000000[6][287:256] <= 32'hD3711002;
            reg_val_0_80000000[6][319:288] <= 32'h27303500;
            reg_val_0_80000000[6][351:320] <= 32'h83234500;
            reg_val_0_80000000[6][383:352] <= 32'h03250500;
            reg_val_0_80000000[6][415:384] <= 32'hF3151000;
            reg_val_0_80000000[6][447:416] <= 32'h13060000;
            reg_val_0_80000000[6][479:448] <= 32'h631AD526;
            reg_val_0_80000000[6][511:480] <= 32'h63187326;
            reg_val_0_80000000[7][31:0] <= 32'h6396C526;
            reg_val_0_80000000[7][63:32] <= 32'h93013000;
            reg_val_0_80000000[7][95:64] <= 32'h17250000;
            reg_val_0_80000000[7][127:96] <= 32'h130585E5;
            reg_val_0_80000000[7][159:128] <= 32'h07300500;
            reg_val_0_80000000[7][191:160] <= 32'h87308500;
            reg_val_0_80000000[7][223:192] <= 32'h07310501;
            reg_val_0_80000000[7][255:224] <= 32'h83268501;
            reg_val_0_80000000[7][287:256] <= 32'h0323C501;
            reg_val_0_80000000[7][319:288] <= 32'hD3711002;
            reg_val_0_80000000[7][351:320] <= 32'h27303500;
            reg_val_0_80000000[7][383:352] <= 32'h83234500;
            reg_val_0_80000000[7][415:384] <= 32'h03250500;
            reg_val_0_80000000[7][447:416] <= 32'hF3151000;
            reg_val_0_80000000[7][479:448] <= 32'h13061000;
            reg_val_0_80000000[7][511:480] <= 32'h6318D522;
            reg_val_0_80000000[8][31:0] <= 32'h63167322;
            reg_val_0_80000000[8][63:32] <= 32'h6394C522;
            reg_val_0_80000000[8][95:64] <= 32'h93014000;
            reg_val_0_80000000[8][127:96] <= 32'h17250000;
            reg_val_0_80000000[8][159:128] <= 32'h130545E3;
            reg_val_0_80000000[8][191:160] <= 32'h07300500;
            reg_val_0_80000000[8][223:192] <= 32'h87308500;
            reg_val_0_80000000[8][255:224] <= 32'h07310501;
            reg_val_0_80000000[8][287:256] <= 32'h83268501;
            reg_val_0_80000000[8][319:288] <= 32'h0323C501;
            reg_val_0_80000000[8][351:320] <= 32'hD3711002;
            reg_val_0_80000000[8][383:352] <= 32'h27303500;
            reg_val_0_80000000[8][415:384] <= 32'h83234500;
            reg_val_0_80000000[8][447:416] <= 32'h03250500;
            reg_val_0_80000000[8][479:448] <= 32'hF3151000;
            reg_val_0_80000000[8][511:480] <= 32'h13061000;
            reg_val_0_80000000[9][31:0] <= 32'h6316D51E;
            reg_val_0_80000000[9][63:32] <= 32'h6314731E;
            reg_val_0_80000000[9][95:64] <= 32'h6392C51E;
            reg_val_0_80000000[9][127:96] <= 32'h93015000;
            reg_val_0_80000000[9][159:128] <= 32'h17250000;
            reg_val_0_80000000[9][191:160] <= 32'h130505E1;
            reg_val_0_80000000[9][223:192] <= 32'h07300500;
            reg_val_0_80000000[9][255:224] <= 32'h87308500;
            reg_val_0_80000000[9][287:256] <= 32'h07310501;
            reg_val_0_80000000[9][319:288] <= 32'h83268501;
            reg_val_0_80000000[9][351:320] <= 32'h0323C501;
            reg_val_0_80000000[9][383:352] <= 32'hD371100A;
            reg_val_0_80000000[9][415:384] <= 32'h27303500;
            reg_val_0_80000000[9][447:416] <= 32'h83234500;
            reg_val_0_80000000[9][479:448] <= 32'h03250500;
            reg_val_0_80000000[9][511:480] <= 32'hF3151000;
            reg_val_0_80000000[10][31:0] <= 32'h13060000;
            reg_val_0_80000000[10][63:32] <= 32'h6314D51A;
            reg_val_0_80000000[10][95:64] <= 32'h6312731A;
            reg_val_0_80000000[10][127:96] <= 32'h6390C51A;
            reg_val_0_80000000[10][159:128] <= 32'h93016000;
            reg_val_0_80000000[10][191:160] <= 32'h17250000;
            reg_val_0_80000000[10][223:192] <= 32'h1305C5DE;
            reg_val_0_80000000[10][255:224] <= 32'h07300500;
            reg_val_0_80000000[10][287:256] <= 32'h87308500;
            reg_val_0_80000000[10][319:288] <= 32'h07310501;
            reg_val_0_80000000[10][351:320] <= 32'h83268501;
            reg_val_0_80000000[10][383:352] <= 32'h0323C501;
            reg_val_0_80000000[10][415:384] <= 32'hD371100A;
            reg_val_0_80000000[10][447:416] <= 32'h27303500;
            reg_val_0_80000000[10][479:448] <= 32'h83234500;
            reg_val_0_80000000[10][511:480] <= 32'h03250500;
            reg_val_0_80000000[11][31:0] <= 32'hF3151000;
            reg_val_0_80000000[11][63:32] <= 32'h13061000;
            reg_val_0_80000000[11][95:64] <= 32'h6312D516;
            reg_val_0_80000000[11][127:96] <= 32'h63107316;
            reg_val_0_80000000[11][159:128] <= 32'h639EC514;
            reg_val_0_80000000[11][191:160] <= 32'h93017000;
            reg_val_0_80000000[11][223:192] <= 32'h17250000;
            reg_val_0_80000000[11][255:224] <= 32'h130585DC;
            reg_val_0_80000000[11][287:256] <= 32'h07300500;
            reg_val_0_80000000[11][319:288] <= 32'h87308500;
            reg_val_0_80000000[11][351:320] <= 32'h07310501;
            reg_val_0_80000000[11][383:352] <= 32'h83268501;
            reg_val_0_80000000[11][415:384] <= 32'h0323C501;
            reg_val_0_80000000[11][447:416] <= 32'hD371100A;
            reg_val_0_80000000[11][479:448] <= 32'h27303500;
            reg_val_0_80000000[11][511:480] <= 32'h83234500;
            reg_val_0_80000000[12][31:0] <= 32'h03250500;
            reg_val_0_80000000[12][63:32] <= 32'hF3151000;
            reg_val_0_80000000[12][95:64] <= 32'h13061000;
            reg_val_0_80000000[12][127:96] <= 32'h6310D512;
            reg_val_0_80000000[12][159:128] <= 32'h631E7310;
            reg_val_0_80000000[12][191:160] <= 32'h639CC510;
            reg_val_0_80000000[12][223:192] <= 32'h93018000;
            reg_val_0_80000000[12][255:224] <= 32'h17250000;
            reg_val_0_80000000[12][287:256] <= 32'h130545DA;
            reg_val_0_80000000[12][319:288] <= 32'h07300500;
            reg_val_0_80000000[12][351:320] <= 32'h87308500;
            reg_val_0_80000000[12][383:352] <= 32'h07310501;
            reg_val_0_80000000[12][415:384] <= 32'h83268501;
            reg_val_0_80000000[12][447:416] <= 32'h0323C501;
            reg_val_0_80000000[12][479:448] <= 32'hD3711012;
            reg_val_0_80000000[12][511:480] <= 32'h27303500;
            reg_val_0_80000000[13][31:0] <= 32'h83234500;
            reg_val_0_80000000[13][63:32] <= 32'h03250500;
            reg_val_0_80000000[13][95:64] <= 32'hF3151000;
            reg_val_0_80000000[13][127:96] <= 32'h13060000;
            reg_val_0_80000000[13][159:128] <= 32'h631ED50C;
            reg_val_0_80000000[13][191:160] <= 32'h631C730C;
            reg_val_0_80000000[13][223:192] <= 32'h639AC50C;
            reg_val_0_80000000[13][255:224] <= 32'h93019000;
            reg_val_0_80000000[13][287:256] <= 32'h17250000;
            reg_val_0_80000000[13][319:288] <= 32'h130505D8;
            reg_val_0_80000000[13][351:320] <= 32'h07300500;
            reg_val_0_80000000[13][383:352] <= 32'h87308500;
            reg_val_0_80000000[13][415:384] <= 32'h07310501;
            reg_val_0_80000000[13][447:416] <= 32'h83268501;
            reg_val_0_80000000[13][479:448] <= 32'h0323C501;
            reg_val_0_80000000[13][511:480] <= 32'hD3711012;
            reg_val_0_80000000[14][31:0] <= 32'h27303500;
            reg_val_0_80000000[14][63:32] <= 32'h83234500;
            reg_val_0_80000000[14][95:64] <= 32'h03250500;
            reg_val_0_80000000[14][127:96] <= 32'hF3151000;
            reg_val_0_80000000[14][159:128] <= 32'h13061000;
            reg_val_0_80000000[14][191:160] <= 32'h631CD508;
            reg_val_0_80000000[14][223:192] <= 32'h631A7308;
            reg_val_0_80000000[14][255:224] <= 32'h6398C508;
            reg_val_0_80000000[14][287:256] <= 32'h9301A000;
            reg_val_0_80000000[14][319:288] <= 32'h17250000;
            reg_val_0_80000000[14][351:320] <= 32'h1305C5D5;
            reg_val_0_80000000[14][383:352] <= 32'h07300500;
            reg_val_0_80000000[14][415:384] <= 32'h87308500;
            reg_val_0_80000000[14][447:416] <= 32'h07310501;
            reg_val_0_80000000[14][479:448] <= 32'h83268501;
            reg_val_0_80000000[14][511:480] <= 32'h0323C501;
            reg_val_0_80000000[15][31:0] <= 32'hD3711012;
            reg_val_0_80000000[15][63:32] <= 32'h27303500;
            reg_val_0_80000000[15][95:64] <= 32'h83234500;
            reg_val_0_80000000[15][127:96] <= 32'h03250500;
            reg_val_0_80000000[15][159:128] <= 32'hF3151000;
            reg_val_0_80000000[15][191:160] <= 32'h13061000;
            reg_val_0_80000000[15][223:192] <= 32'h631AD504;
            reg_val_0_80000000[15][255:224] <= 32'h63187304;
            reg_val_0_80000000[15][287:256] <= 32'h6396C504;
            reg_val_0_80000000[15][319:288] <= 32'h9301B000;
            reg_val_0_80000000[15][351:320] <= 32'h17250000;
            reg_val_0_80000000[15][383:352] <= 32'h130585D3;
            reg_val_0_80000000[15][415:384] <= 32'h07300500;
            reg_val_0_80000000[15][447:416] <= 32'h87308500;
            reg_val_0_80000000[15][479:448] <= 32'h07310501;
            reg_val_0_80000000[15][511:480] <= 32'h83268501;
            reg_val_0_80000000[16][31:0] <= 32'h0323C501;
            reg_val_0_80000000[16][63:32] <= 32'hD371100A;
            reg_val_0_80000000[16][95:64] <= 32'h27303500;
            reg_val_0_80000000[16][127:96] <= 32'h83234500;
            reg_val_0_80000000[16][159:128] <= 32'h03250500;
            reg_val_0_80000000[16][191:160] <= 32'hF3151000;
            reg_val_0_80000000[16][223:192] <= 32'h13060001;
            reg_val_0_80000000[16][255:224] <= 32'h6318D500;
            reg_val_0_80000000[16][287:256] <= 32'h63167300;
            reg_val_0_80000000[16][319:288] <= 32'h6394C500;
            reg_val_0_80000000[16][351:320] <= 32'h63103002;
            reg_val_0_80000000[16][383:352] <= 32'h0F00F00F;
            reg_val_0_80000000[16][415:384] <= 32'h63800100;
            reg_val_0_80000000[16][447:416] <= 32'h93911100;
            reg_val_0_80000000[16][479:448] <= 32'h93E11100;
            reg_val_0_80000000[16][511:480] <= 32'h9308D005;
            reg_val_0_80000000[17][31:0] <= 32'h13850100;
            reg_val_0_80000000[17][63:32] <= 32'h73000000;
            reg_val_0_80000000[17][95:64] <= 32'h0F00F00F;
            reg_val_0_80000000[17][127:96] <= 32'h93011000;
            reg_val_0_80000000[17][159:128] <= 32'h9308D005;
            reg_val_0_80000000[17][191:160] <= 32'h13050000;
            reg_val_0_80000000[17][223:192] <= 32'h73000000;
            reg_val_0_80000000[17][255:224] <= 32'h731000C0;
            reg_val_0_80000000[17][287:256] <= 32'h00000000;
            reg_val_0_80000000[17][319:288] <= 32'h00000000;
            reg_val_0_80000000[17][351:320] <= 32'h00000000;
            reg_val_0_80000000[17][383:352] <= 32'h00000000;
            reg_val_0_80000000[17][415:384] <= 32'h00000000;
            reg_val_0_80000000[17][447:416] <= 32'h00000000;
            reg_val_0_80000000[17][479:448] <= 32'h00000000;
            // fill-in reset values:
            reg_val_0_80000000[17][511:480] <= 32'h00000000;
            reg_val_0_80000000[18][31:0] <= 32'h00000000;
            reg_val_0_80000000[18][63:32] <= 32'h00000000;
            reg_val_0_80000000[18][95:64] <= 32'h00000000;
            reg_val_0_80000000[18][127:96] <= 32'h00000000;
            reg_val_0_80000000[18][159:128] <= 32'h00000000;
            reg_val_0_80000000[18][191:160] <= 32'h00000000;
            reg_val_0_80000000[18][223:192] <= 32'h00000000;
            reg_val_0_80000000[18][255:224] <= 32'h00000000;
            reg_val_0_80000000[18][287:256] <= 32'h00000000;
            reg_val_0_80000000[18][319:288] <= 32'h00000000;
            reg_val_0_80000000[18][351:320] <= 32'h00000000;
            reg_val_0_80000000[18][383:352] <= 32'h00000000;
            reg_val_0_80000000[18][415:384] <= 32'h00000000;
            reg_val_0_80000000[18][447:416] <= 32'h00000000;
            reg_val_0_80000000[18][479:448] <= 32'h00000000;
            reg_val_0_80000000[18][511:480] <= 32'h00000000;
            reg_val_0_80000000[19][31:0] <= 32'h00000000;
            reg_val_0_80000000[19][63:32] <= 32'h00000000;
            reg_val_0_80000000[19][95:64] <= 32'h00000000;
            reg_val_0_80000000[19][127:96] <= 32'h00000000;
            reg_val_0_80000000[19][159:128] <= 32'h00000000;
            reg_val_0_80000000[19][191:160] <= 32'h00000000;
            reg_val_0_80000000[19][223:192] <= 32'h00000000;
            reg_val_0_80000000[19][255:224] <= 32'h00000000;
            reg_val_0_80000000[19][287:256] <= 32'h00000000;
            reg_val_0_80000000[19][319:288] <= 32'h00000000;
            reg_val_0_80000000[19][351:320] <= 32'h00000000;
            reg_val_0_80000000[19][383:352] <= 32'h00000000;
            reg_val_0_80000000[19][415:384] <= 32'h00000000;
            reg_val_0_80000000[19][447:416] <= 32'h00000000;
            reg_val_0_80000000[19][479:448] <= 32'h00000000;
            reg_val_0_80000000[19][511:480] <= 32'h00000000;
            reg_val_0_80000000[20][31:0] <= 32'h00000000;
            reg_val_0_80000000[20][63:32] <= 32'h00000000;
            reg_val_0_80000000[20][95:64] <= 32'h00000000;
            reg_val_0_80000000[20][127:96] <= 32'h00000000;
            reg_val_0_80000000[20][159:128] <= 32'h00000000;
            reg_val_0_80000000[20][191:160] <= 32'h00000000;
            reg_val_0_80000000[20][223:192] <= 32'h00000000;
            reg_val_0_80000000[20][255:224] <= 32'h00000000;
            reg_val_0_80000000[20][287:256] <= 32'h00000000;
            reg_val_0_80000000[20][319:288] <= 32'h00000000;
            reg_val_0_80000000[20][351:320] <= 32'h00000000;
            reg_val_0_80000000[20][383:352] <= 32'h00000000;
            reg_val_0_80000000[20][415:384] <= 32'h00000000;
            reg_val_0_80000000[20][447:416] <= 32'h00000000;
            reg_val_0_80000000[20][479:448] <= 32'h00000000;
            reg_val_0_80000000[20][511:480] <= 32'h00000000;
            reg_val_0_80000000[21][31:0] <= 32'h00000000;
            reg_val_0_80000000[21][63:32] <= 32'h00000000;
            reg_val_0_80000000[21][95:64] <= 32'h00000000;
            reg_val_0_80000000[21][127:96] <= 32'h00000000;
            reg_val_0_80000000[21][159:128] <= 32'h00000000;
            reg_val_0_80000000[21][191:160] <= 32'h00000000;
            reg_val_0_80000000[21][223:192] <= 32'h00000000;
            reg_val_0_80000000[21][255:224] <= 32'h00000000;
            reg_val_0_80000000[21][287:256] <= 32'h00000000;
            reg_val_0_80000000[21][319:288] <= 32'h00000000;
            reg_val_0_80000000[21][351:320] <= 32'h00000000;
            reg_val_0_80000000[21][383:352] <= 32'h00000000;
            reg_val_0_80000000[21][415:384] <= 32'h00000000;
            reg_val_0_80000000[21][447:416] <= 32'h00000000;
            reg_val_0_80000000[21][479:448] <= 32'h00000000;
            reg_val_0_80000000[21][511:480] <= 32'h00000000;
            reg_val_0_80000000[22][31:0] <= 32'h00000000;
            reg_val_0_80000000[22][63:32] <= 32'h00000000;
            reg_val_0_80000000[22][95:64] <= 32'h00000000;
            reg_val_0_80000000[22][127:96] <= 32'h00000000;
            reg_val_0_80000000[22][159:128] <= 32'h00000000;
            reg_val_0_80000000[22][191:160] <= 32'h00000000;
            reg_val_0_80000000[22][223:192] <= 32'h00000000;
            reg_val_0_80000000[22][255:224] <= 32'h00000000;
            reg_val_0_80000000[22][287:256] <= 32'h00000000;
            reg_val_0_80000000[22][319:288] <= 32'h00000000;
            reg_val_0_80000000[22][351:320] <= 32'h00000000;
            reg_val_0_80000000[22][383:352] <= 32'h00000000;
            reg_val_0_80000000[22][415:384] <= 32'h00000000;
            reg_val_0_80000000[22][447:416] <= 32'h00000000;
            reg_val_0_80000000[22][479:448] <= 32'h00000000;
            reg_val_0_80000000[22][511:480] <= 32'h00000000;
            reg_val_0_80000000[23][31:0] <= 32'h00000000;
            reg_val_0_80000000[23][63:32] <= 32'h00000000;
            reg_val_0_80000000[23][95:64] <= 32'h00000000;
            reg_val_0_80000000[23][127:96] <= 32'h00000000;
            reg_val_0_80000000[23][159:128] <= 32'h00000000;
            reg_val_0_80000000[23][191:160] <= 32'h00000000;
            reg_val_0_80000000[23][223:192] <= 32'h00000000;
            reg_val_0_80000000[23][255:224] <= 32'h00000000;
            reg_val_0_80000000[23][287:256] <= 32'h00000000;
            reg_val_0_80000000[23][319:288] <= 32'h00000000;
            reg_val_0_80000000[23][351:320] <= 32'h00000000;
            reg_val_0_80000000[23][383:352] <= 32'h00000000;
            reg_val_0_80000000[23][415:384] <= 32'h00000000;
            reg_val_0_80000000[23][447:416] <= 32'h00000000;
            reg_val_0_80000000[23][479:448] <= 32'h00000000;
            reg_val_0_80000000[23][511:480] <= 32'h00000000;
            reg_val_0_80000000[24][31:0] <= 32'h00000000;
            reg_val_0_80000000[24][63:32] <= 32'h00000000;
            reg_val_0_80000000[24][95:64] <= 32'h00000000;
            reg_val_0_80000000[24][127:96] <= 32'h00000000;
            reg_val_0_80000000[24][159:128] <= 32'h00000000;
            reg_val_0_80000000[24][191:160] <= 32'h00000000;
            reg_val_0_80000000[24][223:192] <= 32'h00000000;
            reg_val_0_80000000[24][255:224] <= 32'h00000000;
            reg_val_0_80000000[24][287:256] <= 32'h00000000;
            reg_val_0_80000000[24][319:288] <= 32'h00000000;
            reg_val_0_80000000[24][351:320] <= 32'h00000000;
            reg_val_0_80000000[24][383:352] <= 32'h00000000;
            reg_val_0_80000000[24][415:384] <= 32'h00000000;
            reg_val_0_80000000[24][447:416] <= 32'h00000000;
            reg_val_0_80000000[24][479:448] <= 32'h00000000;
            reg_val_0_80000000[24][511:480] <= 32'h00000000;
            reg_val_0_80000000[25][31:0] <= 32'h00000000;
            reg_val_0_80000000[25][63:32] <= 32'h00000000;
            reg_val_0_80000000[25][95:64] <= 32'h00000000;
            reg_val_0_80000000[25][127:96] <= 32'h00000000;
            reg_val_0_80000000[25][159:128] <= 32'h00000000;
            reg_val_0_80000000[25][191:160] <= 32'h00000000;
            reg_val_0_80000000[25][223:192] <= 32'h00000000;
            reg_val_0_80000000[25][255:224] <= 32'h00000000;
            reg_val_0_80000000[25][287:256] <= 32'h00000000;
            reg_val_0_80000000[25][319:288] <= 32'h00000000;
            reg_val_0_80000000[25][351:320] <= 32'h00000000;
            reg_val_0_80000000[25][383:352] <= 32'h00000000;
            reg_val_0_80000000[25][415:384] <= 32'h00000000;
            reg_val_0_80000000[25][447:416] <= 32'h00000000;
            reg_val_0_80000000[25][479:448] <= 32'h00000000;
            reg_val_0_80000000[25][511:480] <= 32'h00000000;
            reg_val_0_80000000[26][31:0] <= 32'h00000000;
            reg_val_0_80000000[26][63:32] <= 32'h00000000;
            reg_val_0_80000000[26][95:64] <= 32'h00000000;
            reg_val_0_80000000[26][127:96] <= 32'h00000000;
            reg_val_0_80000000[26][159:128] <= 32'h00000000;
            reg_val_0_80000000[26][191:160] <= 32'h00000000;
            reg_val_0_80000000[26][223:192] <= 32'h00000000;
            reg_val_0_80000000[26][255:224] <= 32'h00000000;
            reg_val_0_80000000[26][287:256] <= 32'h00000000;
            reg_val_0_80000000[26][319:288] <= 32'h00000000;
            reg_val_0_80000000[26][351:320] <= 32'h00000000;
            reg_val_0_80000000[26][383:352] <= 32'h00000000;
            reg_val_0_80000000[26][415:384] <= 32'h00000000;
            reg_val_0_80000000[26][447:416] <= 32'h00000000;
            reg_val_0_80000000[26][479:448] <= 32'h00000000;
            reg_val_0_80000000[26][511:480] <= 32'h00000000;
            reg_val_0_80000000[27][31:0] <= 32'h00000000;
            reg_val_0_80000000[27][63:32] <= 32'h00000000;
            reg_val_0_80000000[27][95:64] <= 32'h00000000;
            reg_val_0_80000000[27][127:96] <= 32'h00000000;
            reg_val_0_80000000[27][159:128] <= 32'h00000000;
            reg_val_0_80000000[27][191:160] <= 32'h00000000;
            reg_val_0_80000000[27][223:192] <= 32'h00000000;
            reg_val_0_80000000[27][255:224] <= 32'h00000000;
            reg_val_0_80000000[27][287:256] <= 32'h00000000;
            reg_val_0_80000000[27][319:288] <= 32'h00000000;
            reg_val_0_80000000[27][351:320] <= 32'h00000000;
            reg_val_0_80000000[27][383:352] <= 32'h00000000;
            reg_val_0_80000000[27][415:384] <= 32'h00000000;
            reg_val_0_80000000[27][447:416] <= 32'h00000000;
            reg_val_0_80000000[27][479:448] <= 32'h00000000;
            reg_val_0_80000000[27][511:480] <= 32'h00000000;
            reg_val_0_80000000[28][31:0] <= 32'h00000000;
            reg_val_0_80000000[28][63:32] <= 32'h00000000;
            reg_val_0_80000000[28][95:64] <= 32'h00000000;
            reg_val_0_80000000[28][127:96] <= 32'h00000000;
            reg_val_0_80000000[28][159:128] <= 32'h00000000;
            reg_val_0_80000000[28][191:160] <= 32'h00000000;
            reg_val_0_80000000[28][223:192] <= 32'h00000000;
            reg_val_0_80000000[28][255:224] <= 32'h00000000;
            reg_val_0_80000000[28][287:256] <= 32'h00000000;
            reg_val_0_80000000[28][319:288] <= 32'h00000000;
            reg_val_0_80000000[28][351:320] <= 32'h00000000;
            reg_val_0_80000000[28][383:352] <= 32'h00000000;
            reg_val_0_80000000[28][415:384] <= 32'h00000000;
            reg_val_0_80000000[28][447:416] <= 32'h00000000;
            reg_val_0_80000000[28][479:448] <= 32'h00000000;
            reg_val_0_80000000[28][511:480] <= 32'h00000000;
            reg_val_0_80000000[29][31:0] <= 32'h00000000;
            reg_val_0_80000000[29][63:32] <= 32'h00000000;
            reg_val_0_80000000[29][95:64] <= 32'h00000000;
            reg_val_0_80000000[29][127:96] <= 32'h00000000;
            reg_val_0_80000000[29][159:128] <= 32'h00000000;
            reg_val_0_80000000[29][191:160] <= 32'h00000000;
            reg_val_0_80000000[29][223:192] <= 32'h00000000;
            reg_val_0_80000000[29][255:224] <= 32'h00000000;
            reg_val_0_80000000[29][287:256] <= 32'h00000000;
            reg_val_0_80000000[29][319:288] <= 32'h00000000;
            reg_val_0_80000000[29][351:320] <= 32'h00000000;
            reg_val_0_80000000[29][383:352] <= 32'h00000000;
            reg_val_0_80000000[29][415:384] <= 32'h00000000;
            reg_val_0_80000000[29][447:416] <= 32'h00000000;
            reg_val_0_80000000[29][479:448] <= 32'h00000000;
            reg_val_0_80000000[29][511:480] <= 32'h00000000;
            reg_val_0_80000000[30][31:0] <= 32'h00000000;
            reg_val_0_80000000[30][63:32] <= 32'h00000000;
            reg_val_0_80000000[30][95:64] <= 32'h00000000;
            reg_val_0_80000000[30][127:96] <= 32'h00000000;
            reg_val_0_80000000[30][159:128] <= 32'h00000000;
            reg_val_0_80000000[30][191:160] <= 32'h00000000;
            reg_val_0_80000000[30][223:192] <= 32'h00000000;
            reg_val_0_80000000[30][255:224] <= 32'h00000000;
            reg_val_0_80000000[30][287:256] <= 32'h00000000;
            reg_val_0_80000000[30][319:288] <= 32'h00000000;
            reg_val_0_80000000[30][351:320] <= 32'h00000000;
            reg_val_0_80000000[30][383:352] <= 32'h00000000;
            reg_val_0_80000000[30][415:384] <= 32'h00000000;
            reg_val_0_80000000[30][447:416] <= 32'h00000000;
            reg_val_0_80000000[30][479:448] <= 32'h00000000;
            reg_val_0_80000000[30][511:480] <= 32'h00000000;
            reg_val_0_80000000[31][31:0] <= 32'h00000000;
            reg_val_0_80000000[31][63:32] <= 32'h00000000;
            reg_val_0_80000000[31][95:64] <= 32'h00000000;
            reg_val_0_80000000[31][127:96] <= 32'h00000000;
            reg_val_0_80000000[31][159:128] <= 32'h00000000;
            reg_val_0_80000000[31][191:160] <= 32'h00000000;
            reg_val_0_80000000[31][223:192] <= 32'h00000000;
            reg_val_0_80000000[31][255:224] <= 32'h00000000;
            reg_val_0_80000000[31][287:256] <= 32'h00000000;
            reg_val_0_80000000[31][319:288] <= 32'h00000000;
            reg_val_0_80000000[31][351:320] <= 32'h00000000;
            reg_val_0_80000000[31][383:352] <= 32'h00000000;
            reg_val_0_80000000[31][415:384] <= 32'h00000000;
            reg_val_0_80000000[31][447:416] <= 32'h00000000;
            reg_val_0_80000000[31][479:448] <= 32'h00000000;
            reg_val_0_80000000[31][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_0_80000000 = next_reg_val_0_80000000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_0_80000000
        // hold reg val by default
        for (int i = 0; i < 32; i++)
        begin
            next_reg_val_0_80000000[i] = reg_val_0_80000000[i];
        end
        // update reg val if wen
        if (wen_0_80000000)
        begin
            next_reg_val_0_80000000[wsel_0_80000000] = wdata_0_80000000;
        end
    end
    
    always_comb begin : READ_LOGIC_0_80000000
        // read val at rsel
        rdata_0_80000000 = reg_val_0_80000000[rsel_0_80000000];
    end
    
    // chunk 1
    logic wen_1_80001000;
    logic [1-1:0] wsel_1_80001000;
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_1_80001000;
    logic [1-1:0] rsel_1_80001000;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_1_80001000;
    
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_1_80001000 [2-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_1_80001000 [2-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_1_80001000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_1_80001000[0][31:0] <= 32'h00000000;
            reg_val_1_80001000[0][63:32] <= 32'h00000000;
            reg_val_1_80001000[0][95:64] <= 32'h00000000;
            reg_val_1_80001000[0][127:96] <= 32'h00000000;
            reg_val_1_80001000[0][159:128] <= 32'h00000000;
            reg_val_1_80001000[0][191:160] <= 32'h00000000;
            reg_val_1_80001000[0][223:192] <= 32'h00000000;
            reg_val_1_80001000[0][255:224] <= 32'h00000000;
            reg_val_1_80001000[0][287:256] <= 32'h00000000;
            reg_val_1_80001000[0][319:288] <= 32'h00000000;
            reg_val_1_80001000[0][351:320] <= 32'h00000000;
            reg_val_1_80001000[0][383:352] <= 32'h00000000;
            reg_val_1_80001000[0][415:384] <= 32'h00000000;
            reg_val_1_80001000[0][447:416] <= 32'h00000000;
            reg_val_1_80001000[0][479:448] <= 32'h00000000;
            reg_val_1_80001000[0][511:480] <= 32'h00000000;
            reg_val_1_80001000[1][31:0] <= 32'h00000000;
            reg_val_1_80001000[1][63:32] <= 32'h00000000;
            // fill-in reset values:
            reg_val_1_80001000[1][95:64] <= 32'h00000000;
            reg_val_1_80001000[1][127:96] <= 32'h00000000;
            reg_val_1_80001000[1][159:128] <= 32'h00000000;
            reg_val_1_80001000[1][191:160] <= 32'h00000000;
            reg_val_1_80001000[1][223:192] <= 32'h00000000;
            reg_val_1_80001000[1][255:224] <= 32'h00000000;
            reg_val_1_80001000[1][287:256] <= 32'h00000000;
            reg_val_1_80001000[1][319:288] <= 32'h00000000;
            reg_val_1_80001000[1][351:320] <= 32'h00000000;
            reg_val_1_80001000[1][383:352] <= 32'h00000000;
            reg_val_1_80001000[1][415:384] <= 32'h00000000;
            reg_val_1_80001000[1][447:416] <= 32'h00000000;
            reg_val_1_80001000[1][479:448] <= 32'h00000000;
            reg_val_1_80001000[1][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_1_80001000 = next_reg_val_1_80001000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_1_80001000
        // hold reg val by default
        for (int i = 0; i < 2; i++)
        begin
            next_reg_val_1_80001000[i] = reg_val_1_80001000[i];
        end
        // update reg val if wen
        if (wen_1_80001000)
        begin
            next_reg_val_1_80001000[wsel_1_80001000] = wdata_1_80001000;
        end
    end
    
    always_comb begin : READ_LOGIC_1_80001000
        // read val at rsel
        rdata_1_80001000 = reg_val_1_80001000[rsel_1_80001000];
    end
    
    // chunk 2
    logic wen_2_80002000;
    logic [3-1:0] wsel_2_80002000;
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_2_80002000;
    logic [3-1:0] rsel_2_80002000;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_2_80002000;
    
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_2_80002000 [8-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_2_80002000 [8-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_2_80002000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_2_80002000[0][31:0] <= 32'h00000000;
            reg_val_2_80002000[0][63:32] <= 32'h00000440;
            reg_val_2_80002000[0][95:64] <= 32'h00000000;
            reg_val_2_80002000[0][127:96] <= 32'h0000F03F;
            reg_val_2_80002000[0][159:128] <= 32'h00000000;
            reg_val_2_80002000[0][191:160] <= 32'h00000000;
            reg_val_2_80002000[0][223:192] <= 32'h00000000;
            reg_val_2_80002000[0][255:224] <= 32'h00000C40;
            reg_val_2_80002000[0][287:256] <= 32'h66666666;
            reg_val_2_80002000[0][319:288] <= 32'h664C93C0;
            reg_val_2_80002000[0][351:320] <= 32'h9A999999;
            reg_val_2_80002000[0][383:352] <= 32'h9999F13F;
            reg_val_2_80002000[0][415:384] <= 32'h00000000;
            reg_val_2_80002000[0][447:416] <= 32'h00000000;
            reg_val_2_80002000[0][479:448] <= 32'h00000000;
            reg_val_2_80002000[0][511:480] <= 32'h004893C0;
            reg_val_2_80002000[1][31:0] <= 32'hF1D4C853;
            reg_val_2_80002000[1][63:32] <= 32'hFB210940;
            reg_val_2_80002000[1][95:64] <= 32'h3A8C30E2;
            reg_val_2_80002000[1][127:96] <= 32'h8E79453E;
            reg_val_2_80002000[1][159:128] <= 32'h00000000;
            reg_val_2_80002000[1][191:160] <= 32'h00000000;
            reg_val_2_80002000[1][223:192] <= 32'hDF6D2055;
            reg_val_2_80002000[1][255:224] <= 32'hFB210940;
            reg_val_2_80002000[1][287:256] <= 32'h00000000;
            reg_val_2_80002000[1][319:288] <= 32'h00000440;
            reg_val_2_80002000[1][351:320] <= 32'h00000000;
            reg_val_2_80002000[1][383:352] <= 32'h0000F03F;
            reg_val_2_80002000[1][415:384] <= 32'h00000000;
            reg_val_2_80002000[1][447:416] <= 32'h00000000;
            reg_val_2_80002000[1][479:448] <= 32'h00000000;
            reg_val_2_80002000[1][511:480] <= 32'h0000F83F;
            reg_val_2_80002000[2][31:0] <= 32'h66666666;
            reg_val_2_80002000[2][63:32] <= 32'h664C93C0;
            reg_val_2_80002000[2][95:64] <= 32'h9A999999;
            reg_val_2_80002000[2][127:96] <= 32'h9999F1BF;
            reg_val_2_80002000[2][159:128] <= 32'h00000000;
            reg_val_2_80002000[2][191:160] <= 32'h00000000;
            reg_val_2_80002000[2][223:192] <= 32'h00000000;
            reg_val_2_80002000[2][255:224] <= 32'h004893C0;
            reg_val_2_80002000[2][287:256] <= 32'hF1D4C853;
            reg_val_2_80002000[2][319:288] <= 32'hFB210940;
            reg_val_2_80002000[2][351:320] <= 32'h3A8C30E2;
            reg_val_2_80002000[2][383:352] <= 32'h8E79453E;
            reg_val_2_80002000[2][415:384] <= 32'h00000000;
            reg_val_2_80002000[2][447:416] <= 32'h00000000;
            reg_val_2_80002000[2][479:448] <= 32'h033C7152;
            reg_val_2_80002000[2][511:480] <= 32'hFB210940;
            reg_val_2_80002000[3][31:0] <= 32'h00000000;
            reg_val_2_80002000[3][63:32] <= 32'h00000440;
            reg_val_2_80002000[3][95:64] <= 32'h00000000;
            reg_val_2_80002000[3][127:96] <= 32'h0000F03F;
            reg_val_2_80002000[3][159:128] <= 32'h00000000;
            reg_val_2_80002000[3][191:160] <= 32'h00000000;
            reg_val_2_80002000[3][223:192] <= 32'h00000000;
            reg_val_2_80002000[3][255:224] <= 32'h00000440;
            reg_val_2_80002000[3][287:256] <= 32'h66666666;
            reg_val_2_80002000[3][319:288] <= 32'h664C93C0;
            reg_val_2_80002000[3][351:320] <= 32'h9A999999;
            reg_val_2_80002000[3][383:352] <= 32'h9999F1BF;
            reg_val_2_80002000[3][415:384] <= 32'h00000000;
            reg_val_2_80002000[3][447:416] <= 32'h00000000;
            reg_val_2_80002000[3][479:448] <= 32'h3D0AD7A3;
            reg_val_2_80002000[3][511:480] <= 32'h703A9540;
            reg_val_2_80002000[4][31:0] <= 32'hF1D4C853;
            reg_val_2_80002000[4][63:32] <= 32'hFB210940;
            reg_val_2_80002000[4][95:64] <= 32'h3A8C30E2;
            reg_val_2_80002000[4][127:96] <= 32'h8E79453E;
            reg_val_2_80002000[4][159:128] <= 32'h00000000;
            reg_val_2_80002000[4][191:160] <= 32'h00000000;
            reg_val_2_80002000[4][223:192] <= 32'h09FFC1A5;
            reg_val_2_80002000[4][255:224] <= 32'hC5DD603E;
            reg_val_2_80002000[4][287:256] <= 32'h00000000;
            reg_val_2_80002000[4][319:288] <= 32'h0000F07F;
            reg_val_2_80002000[4][351:320] <= 32'h00000000;
            reg_val_2_80002000[4][383:352] <= 32'h0000F07F;
            reg_val_2_80002000[4][415:384] <= 32'h00000000;
            reg_val_2_80002000[4][447:416] <= 32'h00000000;
            reg_val_2_80002000[4][479:448] <= 32'h00000000;
            reg_val_2_80002000[4][511:480] <= 32'h0000F87F;
            // fill-in reset values:
            reg_val_2_80002000[5][31:0] <= 32'h00000000;
            reg_val_2_80002000[5][63:32] <= 32'h00000000;
            reg_val_2_80002000[5][95:64] <= 32'h00000000;
            reg_val_2_80002000[5][127:96] <= 32'h00000000;
            reg_val_2_80002000[5][159:128] <= 32'h00000000;
            reg_val_2_80002000[5][191:160] <= 32'h00000000;
            reg_val_2_80002000[5][223:192] <= 32'h00000000;
            reg_val_2_80002000[5][255:224] <= 32'h00000000;
            reg_val_2_80002000[5][287:256] <= 32'h00000000;
            reg_val_2_80002000[5][319:288] <= 32'h00000000;
            reg_val_2_80002000[5][351:320] <= 32'h00000000;
            reg_val_2_80002000[5][383:352] <= 32'h00000000;
            reg_val_2_80002000[5][415:384] <= 32'h00000000;
            reg_val_2_80002000[5][447:416] <= 32'h00000000;
            reg_val_2_80002000[5][479:448] <= 32'h00000000;
            reg_val_2_80002000[5][511:480] <= 32'h00000000;
            reg_val_2_80002000[6][31:0] <= 32'h00000000;
            reg_val_2_80002000[6][63:32] <= 32'h00000000;
            reg_val_2_80002000[6][95:64] <= 32'h00000000;
            reg_val_2_80002000[6][127:96] <= 32'h00000000;
            reg_val_2_80002000[6][159:128] <= 32'h00000000;
            reg_val_2_80002000[6][191:160] <= 32'h00000000;
            reg_val_2_80002000[6][223:192] <= 32'h00000000;
            reg_val_2_80002000[6][255:224] <= 32'h00000000;
            reg_val_2_80002000[6][287:256] <= 32'h00000000;
            reg_val_2_80002000[6][319:288] <= 32'h00000000;
            reg_val_2_80002000[6][351:320] <= 32'h00000000;
            reg_val_2_80002000[6][383:352] <= 32'h00000000;
            reg_val_2_80002000[6][415:384] <= 32'h00000000;
            reg_val_2_80002000[6][447:416] <= 32'h00000000;
            reg_val_2_80002000[6][479:448] <= 32'h00000000;
            reg_val_2_80002000[6][511:480] <= 32'h00000000;
            reg_val_2_80002000[7][31:0] <= 32'h00000000;
            reg_val_2_80002000[7][63:32] <= 32'h00000000;
            reg_val_2_80002000[7][95:64] <= 32'h00000000;
            reg_val_2_80002000[7][127:96] <= 32'h00000000;
            reg_val_2_80002000[7][159:128] <= 32'h00000000;
            reg_val_2_80002000[7][191:160] <= 32'h00000000;
            reg_val_2_80002000[7][223:192] <= 32'h00000000;
            reg_val_2_80002000[7][255:224] <= 32'h00000000;
            reg_val_2_80002000[7][287:256] <= 32'h00000000;
            reg_val_2_80002000[7][319:288] <= 32'h00000000;
            reg_val_2_80002000[7][351:320] <= 32'h00000000;
            reg_val_2_80002000[7][383:352] <= 32'h00000000;
            reg_val_2_80002000[7][415:384] <= 32'h00000000;
            reg_val_2_80002000[7][447:416] <= 32'h00000000;
            reg_val_2_80002000[7][479:448] <= 32'h00000000;
            reg_val_2_80002000[7][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_2_80002000 = next_reg_val_2_80002000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_2_80002000
        // hold reg val by default
        for (int i = 0; i < 8; i++)
        begin
            next_reg_val_2_80002000[i] = reg_val_2_80002000[i];
        end
        // update reg val if wen
        if (wen_2_80002000)
        begin
            next_reg_val_2_80002000[wsel_2_80002000] = wdata_2_80002000;
        end
    end
    
    always_comb begin : READ_LOGIC_2_80002000
        // read val at rsel
        rdata_2_80002000 = reg_val_2_80002000[rsel_2_80002000];
    end
    
    // need reg file/chunk selection signal
    logic [2-1:0] chunk_sel;

    // addr hashing logic
    always_comb begin : ADDR_HASHING_LOGIC
        // default as address not out of bounds
        tb_addr_out_of_bounds = 1'b0;
        
        // bad address assertion:
        assert (
            (26'b10000000000000000000000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000000000000 + 32) ||
            (26'b10000000000000000001000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000001000000 + 2) ||
            (26'b10000000000000000010000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000010000000 + 8)
        ) else begin
            $display("mem request at address 0x%h = 0b%b not available in chunks", mem_req_addr, mem_req_addr);
            tb_addr_out_of_bounds = 1'b1;
        end
        
        // bit = 1 branch
        if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 19] == 1'b1)
        begin
            // select chunk @ 0x80002000
            chunk_sel = 2;
        end
        // bit = 0 branch
        else if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 19] == 1'b0)
        begin
            if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 20] == 1'b0)
            begin
                // select chunk @ 0x80000000
                chunk_sel = 0;
            end
            else if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 20] == 1'b1)
            begin
                // select chunk @ 0x80001000
                chunk_sel = 1;
            end
        end
        else
        begin
            $display("error: got to else in high-level branch");
            tb_addr_out_of_bounds = 1'b1;
        end
        
        // hardwired outputs:
        // hardwiring for chunk 0
        wsel_0_80000000 = mem_req_addr[5-1 : 0];
        wdata_0_80000000 = mem_req_data;
        rsel_0_80000000 = mem_req_addr[5-1 : 0];
        // hardwiring for chunk 1
        wsel_1_80001000 = mem_req_addr[1-1 : 0];
        wdata_1_80001000 = mem_req_data;
        rsel_1_80001000 = mem_req_addr[1-1 : 0];
        // hardwiring for chunk 2
        wsel_2_80002000 = mem_req_addr[3-1 : 0];
        wdata_2_80002000 = mem_req_data;
        rsel_2_80002000 = mem_req_addr[3-1 : 0];
        // default outputs:
        mem_rsp_data = '0;
        // chunk wen's:
        wen_0_80000000 = 1'b0;
        wen_1_80001000 = 1'b0;
        wen_2_80002000 = 1'b0;
        
        // case for routing to diff reg file chunks
        casez (chunk_sel)
        
            // select chunk 0 @ 0x80000000
            0:
            begin
                // write routing
                wen_0_80000000 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_0_80000000;
            end
        
            // select chunk 1 @ 0x80001000
            1:
            begin
                // write routing
                wen_1_80001000 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_1_80001000;
            end
        
            // select chunk 2 @ 0x80002000
            2:
            begin
                // write routing
                wen_2_80002000 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_2_80002000;
            end
        
            // shouldn't get here
            default:
            begin
                $display("error: got to default in chunk_sel case");                mem_rsp_data = '0;
                tb_addr_out_of_bounds = 1'b1;
            end
        endcase
    end

    // other combinational logic for memory interface
    always_comb begin : OTHER_MEM_COMB_LOGIC

        mem_req_ready = 1'b1;           // always ready for request
        mem_rsp_valid = mem_req_valid;  // read ready immediately
        mem_rsp_tag = mem_req_tag;      // match req immediately
    end

    // NOTES:
    // don't know what to do with: 
        // mem_req_byteen
        // busy

endmodule
