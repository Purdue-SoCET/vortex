// removed package "fpu_types"
// removed package "gpu_types"
module VX_vortex_to_local_mem (
	clk,
	reset
);
	// Trace: ../../rtl/VX_vortex_local_mem.sv:6:5
	input clk;
	input reset;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:10:5
	wire mem_req_valid;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:11:5
	wire mem_req_rw;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:12:5
	wire [(0 || 0 ? 16 : 64) - 1:0] mem_req_byteen;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:13:5
	wire [(32 - $clog2((0 || 0 ? 16 : 64))) - 1:0] mem_req_addr;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:14:5
	wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_req_data;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:15:5
	wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_req_tag;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:17:5
	wire mem_req_ready;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:21:5
	wire mem_rsp_valid;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:22:5
	wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_rsp_data;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:23:5
	wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_rsp_tag;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:25:5
	wire mem_rsp_ready;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:29:5
	wire busy;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:32:5
	wire tb_addr_out_of_bounds;
	// Trace: ../../rtl/VX_vortex_local_mem.sv:36:5
	Vortex vortex(
		.clk(clk),
		.reset(reset),
		.mem_req_valid(mem_req_valid),
		.mem_req_rw(mem_req_rw),
		.mem_req_byteen(mem_req_byteen),
		.mem_req_addr(mem_req_addr),
		.mem_req_data(mem_req_data),
		.mem_req_tag(mem_req_tag),
		.mem_req_ready(mem_req_ready),
		.mem_rsp_valid(mem_rsp_valid),
		.mem_rsp_data(mem_rsp_data),
		.mem_rsp_tag(mem_rsp_tag),
		.mem_rsp_ready(mem_rsp_ready),
		.busy(busy)
	);
	// Trace: ../../rtl/VX_vortex_local_mem.sv:59:5
	local_mem RAM(
		.clk(clk),
		.reset(reset),
		.mem_req_valid(mem_req_valid),
		.mem_req_rw(mem_req_rw),
		.mem_req_byteen(mem_req_byteen),
		.mem_req_addr(mem_req_addr),
		.mem_req_data(mem_req_data),
		.mem_req_tag(mem_req_tag),
		.mem_req_ready(mem_req_ready),
		.mem_rsp_valid(mem_rsp_valid),
		.mem_rsp_data(mem_rsp_data),
		.mem_rsp_tag(mem_rsp_tag),
		.mem_rsp_ready(mem_rsp_ready),
		.busy(busy),
		.tb_addr_out_of_bounds(tb_addr_out_of_bounds)
	);
endmodule
// removed module with interface ports: VX_alu_unit
module VX_cache_arb (
	clk,
	reset,
	req_valid_in,
	req_rw_in,
	req_byteen_in,
	req_addr_in,
	req_data_in,
	req_tag_in,
	req_ready_in,
	req_valid_out,
	req_rw_out,
	req_byteen_out,
	req_addr_out,
	req_data_out,
	req_tag_out,
	req_ready_out,
	rsp_valid_in,
	rsp_tmask_in,
	rsp_data_in,
	rsp_tag_in,
	rsp_ready_in,
	rsp_valid_out,
	rsp_tmask_out,
	rsp_data_out,
	rsp_tag_out,
	rsp_ready_out
);
	// Trace: ../../rtl/VX_cache_arb.sv:4:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/VX_cache_arb.sv:5:15
	parameter LANES = 1;
	// Trace: ../../rtl/VX_cache_arb.sv:6:15
	parameter DATA_SIZE = 1;
	// Trace: ../../rtl/VX_cache_arb.sv:7:15
	parameter TAG_IN_WIDTH = 1;
	// Trace: ../../rtl/VX_cache_arb.sv:8:15
	parameter TAG_SEL_IDX = 0;
	// Trace: ../../rtl/VX_cache_arb.sv:9:15
	parameter BUFFERED_REQ = 0;
	// Trace: ../../rtl/VX_cache_arb.sv:10:15
	parameter BUFFERED_RSP = 0;
	// Trace: ../../rtl/VX_cache_arb.sv:11:15
	parameter TYPE = "R";
	// Trace: ../../rtl/VX_cache_arb.sv:13:16
	localparam ADDR_WIDTH = 32 - $clog2(DATA_SIZE);
	// Trace: ../../rtl/VX_cache_arb.sv:14:16
	localparam DATA_WIDTH = 8 * DATA_SIZE;
	// Trace: ../../rtl/VX_cache_arb.sv:15:16
	localparam LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: ../../rtl/VX_cache_arb.sv:16:16
	localparam TAG_OUT_WIDTH = TAG_IN_WIDTH + LOG_NUM_REQS;
	// Trace: ../../rtl/VX_cache_arb.sv:18:5
	input wire clk;
	// Trace: ../../rtl/VX_cache_arb.sv:19:5
	input wire reset;
	// Trace: ../../rtl/VX_cache_arb.sv:22:5
	input wire [(NUM_REQS * LANES) - 1:0] req_valid_in;
	// Trace: ../../rtl/VX_cache_arb.sv:23:5
	input wire [(NUM_REQS * LANES) - 1:0] req_rw_in;
	// Trace: ../../rtl/VX_cache_arb.sv:24:5
	input wire [((NUM_REQS * LANES) * DATA_SIZE) - 1:0] req_byteen_in;
	// Trace: ../../rtl/VX_cache_arb.sv:25:5
	input wire [((NUM_REQS * LANES) * ADDR_WIDTH) - 1:0] req_addr_in;
	// Trace: ../../rtl/VX_cache_arb.sv:26:5
	input wire [((NUM_REQS * LANES) * DATA_WIDTH) - 1:0] req_data_in;
	// Trace: ../../rtl/VX_cache_arb.sv:27:5
	input wire [((NUM_REQS * LANES) * TAG_IN_WIDTH) - 1:0] req_tag_in;
	// Trace: ../../rtl/VX_cache_arb.sv:28:5
	output wire [(NUM_REQS * LANES) - 1:0] req_ready_in;
	// Trace: ../../rtl/VX_cache_arb.sv:31:5
	output wire [LANES - 1:0] req_valid_out;
	// Trace: ../../rtl/VX_cache_arb.sv:32:5
	output wire [LANES - 1:0] req_rw_out;
	// Trace: ../../rtl/VX_cache_arb.sv:33:5
	output wire [(LANES * DATA_SIZE) - 1:0] req_byteen_out;
	// Trace: ../../rtl/VX_cache_arb.sv:34:5
	output wire [(LANES * ADDR_WIDTH) - 1:0] req_addr_out;
	// Trace: ../../rtl/VX_cache_arb.sv:35:5
	output wire [(LANES * DATA_WIDTH) - 1:0] req_data_out;
	// Trace: ../../rtl/VX_cache_arb.sv:36:5
	output wire [(LANES * TAG_OUT_WIDTH) - 1:0] req_tag_out;
	// Trace: ../../rtl/VX_cache_arb.sv:37:5
	input wire [LANES - 1:0] req_ready_out;
	// Trace: ../../rtl/VX_cache_arb.sv:40:5
	input wire rsp_valid_in;
	// Trace: ../../rtl/VX_cache_arb.sv:41:5
	input wire [LANES - 1:0] rsp_tmask_in;
	// Trace: ../../rtl/VX_cache_arb.sv:42:5
	input wire [(LANES * DATA_WIDTH) - 1:0] rsp_data_in;
	// Trace: ../../rtl/VX_cache_arb.sv:43:5
	input wire [TAG_OUT_WIDTH - 1:0] rsp_tag_in;
	// Trace: ../../rtl/VX_cache_arb.sv:44:5
	output wire rsp_ready_in;
	// Trace: ../../rtl/VX_cache_arb.sv:47:5
	output wire [NUM_REQS - 1:0] rsp_valid_out;
	// Trace: ../../rtl/VX_cache_arb.sv:48:5
	output wire [(NUM_REQS * LANES) - 1:0] rsp_tmask_out;
	// Trace: ../../rtl/VX_cache_arb.sv:49:5
	output wire [((NUM_REQS * LANES) * DATA_WIDTH) - 1:0] rsp_data_out;
	// Trace: ../../rtl/VX_cache_arb.sv:50:5
	output wire [(NUM_REQS * TAG_IN_WIDTH) - 1:0] rsp_tag_out;
	// Trace: ../../rtl/VX_cache_arb.sv:51:5
	input wire [NUM_REQS - 1:0] rsp_ready_out;
	// Trace: ../../rtl/VX_cache_arb.sv:53:5
	localparam REQ_DATAW = (((TAG_OUT_WIDTH + ADDR_WIDTH) + 1) + DATA_SIZE) + DATA_WIDTH;
	// Trace: ../../rtl/VX_cache_arb.sv:54:5
	localparam RSP_DATAW = (LANES * (1 + DATA_WIDTH)) + TAG_IN_WIDTH;
	// Trace: ../../rtl/VX_cache_arb.sv:56:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_REQS > 1) begin : genblk1
			// Trace: ../../rtl/VX_cache_arb.sv:58:9
			wire [((NUM_REQS * LANES) * REQ_DATAW) - 1:0] req_data_in_merged;
			// Trace: ../../rtl/VX_cache_arb.sv:59:9
			wire [(LANES * REQ_DATAW) - 1:0] req_data_out_merged;
			genvar i;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
				genvar j;
				for (j = 0; j < LANES; j = j + 1) begin : genblk1
					// Trace: ../../rtl/VX_cache_arb.sv:63:17
					wire [TAG_OUT_WIDTH - 1:0] req_tag_in_w;
					// Trace: ../../rtl/VX_cache_arb.sv:65:17
					VX_bits_insert #(
						.N(TAG_IN_WIDTH),
						.S(LOG_NUM_REQS),
						.POS(TAG_SEL_IDX)
					) bits_insert(
						.data_in(req_tag_in[((i * LANES) + j) * TAG_IN_WIDTH+:TAG_IN_WIDTH]),
						.sel_in(sv2v_cast_76B5F_signed(i)),
						.data_out(req_tag_in_w)
					);
					// Trace: ../../rtl/VX_cache_arb.sv:75:17
					assign req_data_in_merged[((i * LANES) + j) * REQ_DATAW+:REQ_DATAW] = {req_tag_in_w, req_addr_in[((i * LANES) + j) * ADDR_WIDTH+:ADDR_WIDTH], req_rw_in[(i * LANES) + j], req_byteen_in[((i * LANES) + j) * DATA_SIZE+:DATA_SIZE], req_data_in[((i * LANES) + j) * DATA_WIDTH+:DATA_WIDTH]};
				end
			end
			// Trace: ../../rtl/VX_cache_arb.sv:79:9
			VX_stream_arbiter #(
				.NUM_REQS(NUM_REQS),
				.LANES(LANES),
				.DATAW(REQ_DATAW),
				.BUFFERED(BUFFERED_REQ),
				.TYPE(TYPE)
			) req_arb(
				.clk(clk),
				.reset(reset),
				.valid_in(req_valid_in),
				.data_in(req_data_in_merged),
				.ready_in(req_ready_in),
				.valid_out(req_valid_out),
				.data_out(req_data_out_merged),
				.ready_out(req_ready_out)
			);
			for (i = 0; i < LANES; i = i + 1) begin : genblk2
				// Trace: ../../rtl/VX_cache_arb.sv:97:13
				assign {req_tag_out[i * TAG_OUT_WIDTH+:TAG_OUT_WIDTH], req_addr_out[i * ADDR_WIDTH+:ADDR_WIDTH], req_rw_out[i], req_byteen_out[i * DATA_SIZE+:DATA_SIZE], req_data_out[i * DATA_WIDTH+:DATA_WIDTH]} = req_data_out_merged[i * REQ_DATAW+:REQ_DATAW];
			end
			// Trace: ../../rtl/VX_cache_arb.sv:102:9
			wire [(NUM_REQS * RSP_DATAW) - 1:0] rsp_data_out_merged;
			// Trace: ../../rtl/VX_cache_arb.sv:104:9
			wire [LOG_NUM_REQS - 1:0] rsp_sel = rsp_tag_in[TAG_SEL_IDX+:LOG_NUM_REQS];
			// Trace: ../../rtl/VX_cache_arb.sv:106:9
			wire [TAG_IN_WIDTH - 1:0] rsp_tag_in_w;
			// Trace: ../../rtl/VX_cache_arb.sv:108:9
			VX_bits_remove #(
				.N(TAG_OUT_WIDTH),
				.S(LOG_NUM_REQS),
				.POS(TAG_SEL_IDX)
			) bits_remove(
				.data_in(rsp_tag_in),
				.data_out(rsp_tag_in_w)
			);
			// Trace: ../../rtl/VX_cache_arb.sv:117:9
			VX_stream_demux #(
				.NUM_REQS(NUM_REQS),
				.LANES(1),
				.DATAW(RSP_DATAW),
				.BUFFERED(BUFFERED_RSP)
			) rsp_demux(
				.clk(clk),
				.reset(reset),
				.sel_in(rsp_sel),
				.valid_in(rsp_valid_in),
				.data_in({rsp_tmask_in, rsp_tag_in_w, rsp_data_in}),
				.ready_in(rsp_ready_in),
				.valid_out(rsp_valid_out),
				.data_out(rsp_data_out_merged),
				.ready_out(rsp_ready_out)
			);
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk3
				// Trace: ../../rtl/VX_cache_arb.sv:135:13
				assign {rsp_tmask_out[i * LANES+:LANES], rsp_tag_out[i * TAG_IN_WIDTH+:TAG_IN_WIDTH], rsp_data_out[DATA_WIDTH * (i * LANES)+:DATA_WIDTH * LANES]} = rsp_data_out_merged[i * RSP_DATAW+:RSP_DATAW];
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/VX_cache_arb.sv:143:9
			assign req_valid_out = req_valid_in;
			// Trace: ../../rtl/VX_cache_arb.sv:144:9
			assign req_tag_out = req_tag_in;
			// Trace: ../../rtl/VX_cache_arb.sv:145:9
			assign req_addr_out = req_addr_in;
			// Trace: ../../rtl/VX_cache_arb.sv:146:9
			assign req_rw_out = req_rw_in;
			// Trace: ../../rtl/VX_cache_arb.sv:147:9
			assign req_byteen_out = req_byteen_in;
			// Trace: ../../rtl/VX_cache_arb.sv:148:9
			assign req_data_out = req_data_in;
			// Trace: ../../rtl/VX_cache_arb.sv:149:9
			assign req_ready_in = req_ready_out;
			// Trace: ../../rtl/VX_cache_arb.sv:151:9
			assign rsp_valid_out = rsp_valid_in;
			// Trace: ../../rtl/VX_cache_arb.sv:152:9
			assign rsp_tmask_out = rsp_tmask_in;
			// Trace: ../../rtl/VX_cache_arb.sv:153:9
			assign rsp_tag_out = rsp_tag_in;
			// Trace: ../../rtl/VX_cache_arb.sv:154:9
			assign rsp_data_out = rsp_data_in;
			// Trace: ../../rtl/VX_cache_arb.sv:155:9
			assign rsp_ready_in = rsp_ready_out;
		end
	endgenerate
endmodule
module VX_cluster (
	clk,
	reset,
	mem_req_valid,
	mem_req_rw,
	mem_req_byteen,
	mem_req_addr,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready,
	busy
);
	// Trace: ../../rtl/VX_cluster.sv:4:15
	parameter CLUSTER_ID = 0;
	// Trace: ../../rtl/VX_cluster.sv:9:5
	input wire clk;
	// Trace: ../../rtl/VX_cluster.sv:10:5
	input wire reset;
	// Trace: ../../rtl/VX_cluster.sv:13:5
	output wire mem_req_valid;
	// Trace: ../../rtl/VX_cluster.sv:14:5
	output wire mem_req_rw;
	// Trace: ../../rtl/VX_cluster.sv:15:5
	output wire [(0 || 0 ? 16 : 64) - 1:0] mem_req_byteen;
	// Trace: ../../rtl/VX_cluster.sv:16:5
	output wire [(32 - $clog2((0 || 0 ? 16 : 64))) - 1:0] mem_req_addr;
	// Trace: ../../rtl/VX_cluster.sv:17:5
	output wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_req_data;
	// Trace: ../../rtl/VX_cluster.sv:18:5
	output wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_req_tag;
	// Trace: ../../rtl/VX_cluster.sv:19:5
	input wire mem_req_ready;
	// Trace: ../../rtl/VX_cluster.sv:22:5
	input wire mem_rsp_valid;
	// Trace: ../../rtl/VX_cluster.sv:23:5
	input wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_rsp_data;
	// Trace: ../../rtl/VX_cluster.sv:24:5
	input wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_rsp_tag;
	// Trace: ../../rtl/VX_cluster.sv:25:5
	output wire mem_rsp_ready;
	// Trace: ../../rtl/VX_cluster.sv:28:5
	output wire busy;
	// Trace: ../../rtl/VX_cluster.sv:32:5
	wire [0:0] per_core_mem_req_valid;
	// Trace: ../../rtl/VX_cluster.sv:33:5
	wire [0:0] per_core_mem_req_rw;
	// Trace: ../../rtl/VX_cluster.sv:34:5
	wire [(0 || 0 ? 16 : 64) - 1:0] per_core_mem_req_byteen;
	// Trace: ../../rtl/VX_cluster.sv:35:5
	wire [(32 - $clog2((0 || 0 ? 16 : 64))) - 1:0] per_core_mem_req_addr;
	// Trace: ../../rtl/VX_cluster.sv:36:5
	wire [((0 || 0 ? 16 : 64) * 8) - 1:0] per_core_mem_req_data;
	// Trace: ../../rtl/VX_cluster.sv:37:5
	wire [(((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0 : (1 - ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0)) + ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) - 1)):(((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? 0 : (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0)] per_core_mem_req_tag;
	// Trace: ../../rtl/VX_cluster.sv:38:5
	wire [0:0] per_core_mem_req_ready;
	// Trace: ../../rtl/VX_cluster.sv:40:5
	wire [0:0] per_core_mem_rsp_valid;
	// Trace: ../../rtl/VX_cluster.sv:41:5
	wire [((0 || 0 ? 16 : 64) * 8) - 1:0] per_core_mem_rsp_data;
	// Trace: ../../rtl/VX_cluster.sv:42:5
	wire [(((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0 : (1 - ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0)) + ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) - 1)):(((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? 0 : (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0)] per_core_mem_rsp_tag;
	// Trace: ../../rtl/VX_cluster.sv:43:5
	wire [0:0] per_core_mem_rsp_ready;
	// Trace: ../../rtl/VX_cluster.sv:45:5
	wire [0:0] per_core_busy;
	// Trace: ../../rtl/VX_cluster.sv:47:5
	genvar i;
	generate
		for (i = 0; i < 1; i = i + 1) begin : genblk1
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_cluster.sv:49:27
			wire core_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_cluster.sv:49:60
			VX_reset_relay __core_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(core_reset)
			);
			// Trace: ../../rtl/VX_cluster.sv:51:9
			VX_core #(.CORE_ID(i + (CLUSTER_ID * 1))) core(
				.clk(clk),
				.reset(core_reset),
				.mem_req_valid(per_core_mem_req_valid[i]),
				.mem_req_rw(per_core_mem_req_rw[i]),
				.mem_req_byteen(per_core_mem_req_byteen[i * (0 || 0 ? 16 : 64)+:(0 || 0 ? 16 : 64)]),
				.mem_req_addr(per_core_mem_req_addr[i * (32 - $clog2((0 || 0 ? 16 : 64)))+:32 - $clog2((0 || 0 ? 16 : 64))]),
				.mem_req_data(per_core_mem_req_data[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8]),
				.mem_req_tag(per_core_mem_req_tag[(((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? 0 : (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) + (i * (((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1 : 1 - ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0)))+:(((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1 : 1 - ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0))]),
				.mem_req_ready(per_core_mem_req_ready[i]),
				.mem_rsp_valid(per_core_mem_rsp_valid[i]),
				.mem_rsp_data(per_core_mem_rsp_data[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8]),
				.mem_rsp_tag(per_core_mem_rsp_tag[(((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? 0 : (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) + (i * (((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1 : 1 - ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0)))+:(((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0) >= 0 ? (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1 : 1 - ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0))]),
				.mem_rsp_ready(per_core_mem_rsp_ready[i]),
				.busy(per_core_busy[i])
			);
		end
	endgenerate
	// Trace: ../../rtl/VX_cluster.sv:76:5
	assign busy = |per_core_busy;
	// Trace: ../../rtl/VX_cluster.sv:78:5
	generate
		if (1) begin : genblk2
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_cluster.sv:147:30
			wire mem_arb_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_cluster.sv:147:63
			VX_reset_relay __mem_arb_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(mem_arb_reset)
			);
			// Trace: ../../rtl/VX_cluster.sv:149:9
			VX_mem_arb #(
				.NUM_REQS(1),
				.DATA_WIDTH((0 || 0 ? 16 : 64) * 8),
				.ADDR_WIDTH(32 - $clog2((0 || 0 ? 16 : 64))),
				.TAG_IN_WIDTH((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1),
				.TYPE("R"),
				.TAG_SEL_IDX(1),
				.BUFFERED_REQ(1),
				.BUFFERED_RSP(1)
			) mem_arb(
				.clk(clk),
				.reset(mem_arb_reset),
				.req_valid_in(per_core_mem_req_valid),
				.req_rw_in(per_core_mem_req_rw),
				.req_byteen_in(per_core_mem_req_byteen),
				.req_addr_in(per_core_mem_req_addr),
				.req_data_in(per_core_mem_req_data),
				.req_tag_in(per_core_mem_req_tag),
				.req_ready_in(per_core_mem_req_ready),
				.req_valid_out(mem_req_valid),
				.req_rw_out(mem_req_rw),
				.req_byteen_out(mem_req_byteen),
				.req_addr_out(mem_req_addr),
				.req_data_out(mem_req_data),
				.req_tag_out(mem_req_tag),
				.req_ready_out(mem_req_ready),
				.rsp_valid_out(per_core_mem_rsp_valid),
				.rsp_data_out(per_core_mem_rsp_data),
				.rsp_tag_out(per_core_mem_rsp_tag),
				.rsp_ready_out(per_core_mem_rsp_ready),
				.rsp_valid_in(mem_rsp_valid),
				.rsp_tag_in(mem_rsp_tag),
				.rsp_data_in(mem_rsp_data),
				.rsp_ready_in(mem_rsp_ready)
			);
		end
	endgenerate
endmodule
// removed module with interface ports: VX_commit
module VX_core (
	clk,
	reset,
	mem_req_valid,
	mem_req_rw,
	mem_req_byteen,
	mem_req_addr,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready,
	busy
);
	// Trace: ../../rtl/VX_core.sv:4:15
	parameter CORE_ID = 0;
	// Trace: ../../rtl/VX_core.sv:9:5
	input wire clk;
	// Trace: ../../rtl/VX_core.sv:10:5
	input wire reset;
	// Trace: ../../rtl/VX_core.sv:13:5
	output wire mem_req_valid;
	// Trace: ../../rtl/VX_core.sv:14:5
	output wire mem_req_rw;
	// Trace: ../../rtl/VX_core.sv:15:5
	output wire [(0 || 0 ? 16 : 64) - 1:0] mem_req_byteen;
	// Trace: ../../rtl/VX_core.sv:16:5
	output wire [(32 - $clog2((0 || 0 ? 16 : 64))) - 1:0] mem_req_addr;
	// Trace: ../../rtl/VX_core.sv:17:5
	output wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_req_data;
	// Trace: ../../rtl/VX_core.sv:18:5
	output wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_req_tag;
	// Trace: ../../rtl/VX_core.sv:19:5
	input wire mem_req_ready;
	// Trace: ../../rtl/VX_core.sv:22:5
	input wire mem_rsp_valid;
	// Trace: ../../rtl/VX_core.sv:23:5
	input wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_rsp_data;
	// Trace: ../../rtl/VX_core.sv:24:5
	input wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_rsp_tag;
	// Trace: ../../rtl/VX_core.sv:25:5
	output wire mem_rsp_ready;
	// Trace: ../../rtl/VX_core.sv:28:5
	output wire busy;
	// Trace: ../../rtl/VX_core.sv:34:5
	// expanded interface instance: mem_req_if
	localparam _param_ABED4_DATA_WIDTH = (0 || 0 ? 16 : 64) * 8;
	localparam _param_ABED4_ADDR_WIDTH = 32 - $clog2((0 || 0 ? 16 : 64));
	localparam _param_ABED4_TAG_WIDTH = (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1;
	generate
		if (1) begin : mem_req_if
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:7:15
			localparam DATA_WIDTH = _param_ABED4_DATA_WIDTH;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:8:15
			localparam ADDR_WIDTH = _param_ABED4_ADDR_WIDTH;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:9:15
			localparam TAG_WIDTH = _param_ABED4_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:10:15
			localparam DATA_SIZE = DATA_WIDTH / 8;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:13:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:14:5
			wire rw;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:15:5
			wire [DATA_SIZE - 1:0] byteen;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:16:5
			wire [ADDR_WIDTH - 1:0] addr;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:17:5
			wire [DATA_WIDTH - 1:0] data;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:18:5
			wire [TAG_WIDTH - 1:0] tag;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:19:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:21:5
			// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:31:5
		end
	endgenerate
	// Trace: ../../rtl/VX_core.sv:40:5
	// expanded interface instance: mem_rsp_if
	localparam _param_F9E76_DATA_WIDTH = (0 || 0 ? 16 : 64) * 8;
	localparam _param_F9E76_TAG_WIDTH = (1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1;
	generate
		if (1) begin : mem_rsp_if
			// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:7:15
			localparam DATA_WIDTH = _param_F9E76_DATA_WIDTH;
			// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:8:15
			localparam TAG_WIDTH = _param_F9E76_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:11:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:12:5
			wire [DATA_WIDTH - 1:0] data;
			// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:13:5
			wire [TAG_WIDTH - 1:0] tag;
			// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:14:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:16:5
			// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:23:5
		end
	endgenerate
	// Trace: ../../rtl/VX_core.sv:45:5
	assign mem_req_valid = mem_req_if.valid;
	// Trace: ../../rtl/VX_core.sv:46:5
	assign mem_req_rw = mem_req_if.rw;
	// Trace: ../../rtl/VX_core.sv:47:5
	assign mem_req_byteen = mem_req_if.byteen;
	// Trace: ../../rtl/VX_core.sv:48:5
	assign mem_req_addr = mem_req_if.addr;
	// Trace: ../../rtl/VX_core.sv:49:5
	assign mem_req_data = mem_req_if.data;
	// Trace: ../../rtl/VX_core.sv:50:5
	assign mem_req_tag = mem_req_if.tag;
	// Trace: ../../rtl/VX_core.sv:51:5
	assign mem_req_if.ready = mem_req_ready;
	// Trace: ../../rtl/VX_core.sv:53:5
	assign mem_rsp_if.valid = mem_rsp_valid;
	// Trace: ../../rtl/VX_core.sv:54:5
	assign mem_rsp_if.data = mem_rsp_data;
	// Trace: ../../rtl/VX_core.sv:55:5
	assign mem_rsp_if.tag = mem_rsp_tag;
	// Trace: ../../rtl/VX_core.sv:56:5
	assign mem_rsp_ready = mem_rsp_if.ready;
	// Trace: ../../rtl/VX_core.sv:60:5
	// expanded interface instance: dcache_req_if
	localparam _param_BD702_NUM_REQS = 2;
	localparam _param_BD702_WORD_SIZE = 4;
	localparam _param_BD702_TAG_WIDTH = 48;
	generate
		if (1) begin : dcache_req_if
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:7:15
			localparam NUM_REQS = _param_BD702_NUM_REQS;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:8:15
			localparam WORD_SIZE = _param_BD702_WORD_SIZE;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:9:15
			localparam TAG_WIDTH = _param_BD702_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:12:5
			wire [1:0] valid;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:13:5
			wire [1:0] rw;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:14:5
			wire [7:0] byteen;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:15:5
			wire [59:0] addr;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:16:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:17:5
			wire [95:0] tag;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:18:5
			wire [1:0] ready;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:20:5
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:30:5
		end
	endgenerate
	// Trace: ../../rtl/VX_core.sv:66:5
	// expanded interface instance: dcache_rsp_if
	localparam _param_2395E_NUM_REQS = 2;
	localparam _param_2395E_WORD_SIZE = 4;
	localparam _param_2395E_TAG_WIDTH = 48;
	generate
		if (1) begin : dcache_rsp_if
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:7:15
			localparam NUM_REQS = _param_2395E_NUM_REQS;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:8:15
			localparam WORD_SIZE = _param_2395E_WORD_SIZE;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:9:15
			localparam TAG_WIDTH = _param_2395E_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:12:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:13:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:14:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:15:5
			wire [47:0] tag;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:16:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:18:5
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:26:5
		end
	endgenerate
	// Trace: ../../rtl/VX_core.sv:72:5
	// expanded interface instance: icache_req_if
	localparam _param_1F99A_WORD_SIZE = 4;
	localparam _param_1F99A_TAG_WIDTH = 45;
	generate
		if (1) begin : icache_req_if
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:7:15
			localparam WORD_SIZE = _param_1F99A_WORD_SIZE;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:8:15
			localparam TAG_WIDTH = _param_1F99A_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:11:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:12:5
			wire [29:0] addr;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:13:5
			wire [44:0] tag;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:14:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:16:5
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:23:5
		end
	endgenerate
	// Trace: ../../rtl/VX_core.sv:77:5
	// expanded interface instance: icache_rsp_if
	localparam _param_396BA_WORD_SIZE = 4;
	localparam _param_396BA_TAG_WIDTH = 45;
	generate
		if (1) begin : icache_rsp_if
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:7:15
			localparam WORD_SIZE = _param_396BA_WORD_SIZE;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:8:15
			localparam TAG_WIDTH = _param_396BA_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:11:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:12:5
			wire [31:0] data;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:13:5
			wire [44:0] tag;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:14:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:16:5
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:23:5
		end
	endgenerate
	// Trace: ../../rtl/VX_core.sv:82:5
	VX_pipeline #(.CORE_ID(CORE_ID)) pipeline(
		.clk(clk),
		.reset(reset),
		.dcache_req_valid(dcache_req_if.valid),
		.dcache_req_rw(dcache_req_if.rw),
		.dcache_req_byteen(dcache_req_if.byteen),
		.dcache_req_addr(dcache_req_if.addr),
		.dcache_req_data(dcache_req_if.data),
		.dcache_req_tag(dcache_req_if.tag),
		.dcache_req_ready(dcache_req_if.ready),
		.dcache_rsp_valid(dcache_rsp_if.valid),
		.dcache_rsp_tmask(dcache_rsp_if.tmask),
		.dcache_rsp_data(dcache_rsp_if.data),
		.dcache_rsp_tag(dcache_rsp_if.tag),
		.dcache_rsp_ready(dcache_rsp_if.ready),
		.icache_req_valid(icache_req_if.valid),
		.icache_req_addr(icache_req_if.addr),
		.icache_req_tag(icache_req_if.tag),
		.icache_req_ready(icache_req_if.ready),
		.icache_rsp_valid(icache_rsp_if.valid),
		.icache_rsp_data(icache_rsp_if.data),
		.icache_rsp_tag(icache_rsp_if.tag),
		.icache_rsp_ready(icache_rsp_if.ready),
		.busy(busy)
	);
	// Trace: ../../rtl/VX_core.sv:127:5
	// expanded module instance: mem_unit
	localparam _param_A06D0_CORE_ID = CORE_ID;
	function automatic [(4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) - 1:0] sv2v_cast_7CD18;
		input reg [(4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) - 1:0] inp;
		sv2v_cast_7CD18 = inp;
	endfunction
	generate
		if (1) begin : mem_unit
			// Trace: ../../rtl/VX_mem_unit.sv:4:15
			localparam CORE_ID = _param_A06D0_CORE_ID;
			// Trace: ../../rtl/VX_mem_unit.sv:8:5
			wire clk;
			// Trace: ../../rtl/VX_mem_unit.sv:9:5
			wire reset;
			// Trace: ../../rtl/VX_mem_unit.sv:16:5
			// removed modport instance dcache_req_if
			// Trace: ../../rtl/VX_mem_unit.sv:17:5
			// removed modport instance dcache_rsp_if
			// Trace: ../../rtl/VX_mem_unit.sv:20:5
			// removed modport instance icache_req_if
			// Trace: ../../rtl/VX_mem_unit.sv:21:5
			// removed modport instance icache_rsp_if
			// Trace: ../../rtl/VX_mem_unit.sv:24:5
			// removed modport instance mem_req_if
			// Trace: ../../rtl/VX_mem_unit.sv:25:5
			// removed modport instance mem_rsp_if
			// Trace: ../../rtl/VX_mem_unit.sv:32:5
			// expanded interface instance: icache_mem_req_if
			localparam _param_03929_DATA_WIDTH = (0 || 0 ? 16 : 64) * 8;
			localparam _param_03929_ADDR_WIDTH = 32 - $clog2((0 || 0 ? 16 : 64));
			localparam _param_03929_TAG_WIDTH = 1;
			if (1) begin : icache_mem_req_if
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:7:15
				localparam DATA_WIDTH = _param_03929_DATA_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:8:15
				localparam ADDR_WIDTH = _param_03929_ADDR_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:9:15
				localparam TAG_WIDTH = _param_03929_TAG_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:10:15
				localparam DATA_SIZE = DATA_WIDTH / 8;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:13:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:14:5
				wire rw;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:15:5
				wire [DATA_SIZE - 1:0] byteen;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:16:5
				wire [ADDR_WIDTH - 1:0] addr;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:17:5
				wire [DATA_WIDTH - 1:0] data;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:18:5
				wire [0:0] tag;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:19:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:21:5
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:31:5
			end
			// Trace: ../../rtl/VX_mem_unit.sv:38:5
			// expanded interface instance: icache_mem_rsp_if
			localparam _param_8D4A5_DATA_WIDTH = (0 || 0 ? 16 : 64) * 8;
			localparam _param_8D4A5_TAG_WIDTH = 1;
			if (1) begin : icache_mem_rsp_if
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:7:15
				localparam DATA_WIDTH = _param_8D4A5_DATA_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:8:15
				localparam TAG_WIDTH = _param_8D4A5_TAG_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:11:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:12:5
				wire [DATA_WIDTH - 1:0] data;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:13:5
				wire [0:0] tag;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:14:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:16:5
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:23:5
			end
			// Trace: ../../rtl/VX_mem_unit.sv:43:5
			// expanded interface instance: dcache_mem_req_if
			localparam _param_B57C2_DATA_WIDTH = (0 || 0 ? 16 : 64) * 8;
			localparam _param_B57C2_ADDR_WIDTH = 32 - $clog2((0 || 0 ? 16 : 64));
			localparam _param_B57C2_TAG_WIDTH = (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48);
			if (1) begin : dcache_mem_req_if
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:7:15
				localparam DATA_WIDTH = _param_B57C2_DATA_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:8:15
				localparam ADDR_WIDTH = _param_B57C2_ADDR_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:9:15
				localparam TAG_WIDTH = _param_B57C2_TAG_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:10:15
				localparam DATA_SIZE = DATA_WIDTH / 8;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:13:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:14:5
				wire rw;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:15:5
				wire [DATA_SIZE - 1:0] byteen;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:16:5
				wire [ADDR_WIDTH - 1:0] addr;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:17:5
				wire [DATA_WIDTH - 1:0] data;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:18:5
				wire [TAG_WIDTH - 1:0] tag;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:19:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:21:5
				// Trace: ../../rtl/interfaces/VX_mem_req_if.sv:31:5
			end
			// Trace: ../../rtl/VX_mem_unit.sv:49:5
			// expanded interface instance: dcache_mem_rsp_if
			localparam _param_79532_DATA_WIDTH = (0 || 0 ? 16 : 64) * 8;
			localparam _param_79532_TAG_WIDTH = (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48);
			if (1) begin : dcache_mem_rsp_if
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:7:15
				localparam DATA_WIDTH = _param_79532_DATA_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:8:15
				localparam TAG_WIDTH = _param_79532_TAG_WIDTH;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:11:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:12:5
				wire [DATA_WIDTH - 1:0] data;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:13:5
				wire [TAG_WIDTH - 1:0] tag;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:14:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:16:5
				// Trace: ../../rtl/interfaces/VX_mem_rsp_if.sv:23:5
			end
			// Trace: ../../rtl/VX_mem_unit.sv:54:5
			// expanded interface instance: dcache_req_tmp_if
			localparam _param_79CA8_NUM_REQS = 2;
			localparam _param_79CA8_WORD_SIZE = 4;
			localparam _param_79CA8_TAG_WIDTH = 47;
			if (1) begin : dcache_req_tmp_if
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:7:15
				localparam NUM_REQS = _param_79CA8_NUM_REQS;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:8:15
				localparam WORD_SIZE = _param_79CA8_WORD_SIZE;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:9:15
				localparam TAG_WIDTH = _param_79CA8_TAG_WIDTH;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:12:5
				wire [1:0] valid;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:13:5
				wire [1:0] rw;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:14:5
				wire [7:0] byteen;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:15:5
				wire [59:0] addr;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:16:5
				wire [63:0] data;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:17:5
				wire [93:0] tag;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:18:5
				wire [1:0] ready;
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:20:5
				// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:30:5
			end
			// Trace: ../../rtl/VX_mem_unit.sv:60:5
			// expanded interface instance: dcache_rsp_tmp_if
			localparam _param_E25F4_NUM_REQS = 2;
			localparam _param_E25F4_WORD_SIZE = 4;
			localparam _param_E25F4_TAG_WIDTH = 47;
			if (1) begin : dcache_rsp_tmp_if
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:7:15
				localparam NUM_REQS = _param_E25F4_NUM_REQS;
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:8:15
				localparam WORD_SIZE = _param_E25F4_WORD_SIZE;
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:9:15
				localparam TAG_WIDTH = _param_E25F4_TAG_WIDTH;
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:12:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:13:5
				wire [1:0] tmask;
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:14:5
				wire [63:0] data;
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:15:5
				wire [46:0] tag;
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:16:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:18:5
				// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:26:5
			end
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:66:25
			wire icache_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:66:58
			VX_reset_relay __icache_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(icache_reset)
			);
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:67:25
			wire dcache_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:67:58
			VX_reset_relay __dcache_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(dcache_reset)
			);
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:68:26
			wire mem_arb_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:68:59
			VX_reset_relay __mem_arb_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(mem_arb_reset)
			);
			// Trace: ../../rtl/VX_mem_unit.sv:70:5
			localparam sv2v_uu_icache_NUM_REQS = 1;
			localparam sv2v_uu_icache_WORD_SIZE = 4;
			// removed localparam type sv2v_uu_icache_core_req_data
			localparam [31:0] sv2v_uu_icache_ext_core_req_data_x = 1'sbx;
			VX_cache #(
				.CACHE_ID((0 + (CORE_ID * 3)) + 0),
				.CACHE_SIZE(16384),
				.CACHE_LINE_SIZE((0 || 0 ? 16 : 64)),
				.NUM_BANKS(1),
				.WORD_SIZE(4),
				.NUM_REQS(1),
				.CREQ_SIZE(0),
				.CRSQ_SIZE(2),
				.MSHR_SIZE(2),
				.MRSQ_SIZE(0),
				.MREQ_SIZE(4),
				.WRITE_ENABLE(0),
				.CORE_TAG_WIDTH(45),
				.CORE_TAG_ID_BITS(1),
				.MEM_TAG_WIDTH(1)
			) icache(
				.clk(clk),
				.reset(icache_reset),
				.core_req_valid(VX_core.icache_req_if.valid),
				.core_req_rw(1'b0),
				.core_req_byteen('b0),
				.core_req_addr(VX_core.icache_req_if.addr),
				.core_req_data(sv2v_uu_icache_ext_core_req_data_x),
				.core_req_tag(VX_core.icache_req_if.tag),
				.core_req_ready(VX_core.icache_req_if.ready),
				.core_rsp_valid(VX_core.icache_rsp_if.valid),
				.core_rsp_data(VX_core.icache_rsp_if.data),
				.core_rsp_tag(VX_core.icache_rsp_if.tag),
				.core_rsp_ready(VX_core.icache_rsp_if.ready),
				.mem_req_valid(icache_mem_req_if.valid),
				.mem_req_rw(icache_mem_req_if.rw),
				.mem_req_byteen(icache_mem_req_if.byteen),
				.mem_req_addr(icache_mem_req_if.addr),
				.mem_req_data(icache_mem_req_if.data),
				.mem_req_tag(icache_mem_req_if.tag),
				.mem_req_ready(icache_mem_req_if.ready),
				.mem_rsp_valid(icache_mem_rsp_if.valid),
				.mem_rsp_data(icache_mem_rsp_if.data),
				.mem_rsp_tag(icache_mem_rsp_if.tag),
				.mem_rsp_ready(icache_mem_rsp_if.ready)
			);
			// Trace: ../../rtl/VX_mem_unit.sv:128:5
			VX_cache #(
				.CACHE_ID((0 + (CORE_ID * 3)) + 1),
				.CACHE_SIZE(16384),
				.CACHE_LINE_SIZE((0 || 0 ? 16 : 64)),
				.NUM_BANKS(2),
				.NUM_PORTS(1),
				.WORD_SIZE(4),
				.NUM_REQS(2),
				.CREQ_SIZE(0),
				.CRSQ_SIZE(2),
				.MSHR_SIZE(4),
				.MRSQ_SIZE(0),
				.MREQ_SIZE(4),
				.WRITE_ENABLE(1),
				.CORE_TAG_WIDTH(47),
				.CORE_TAG_ID_BITS(3),
				.MEM_TAG_WIDTH((4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)),
				.NC_ENABLE(1)
			) dcache(
				.clk(clk),
				.reset(dcache_reset),
				.core_req_valid(dcache_req_tmp_if.valid),
				.core_req_rw(dcache_req_tmp_if.rw),
				.core_req_byteen(dcache_req_tmp_if.byteen),
				.core_req_addr(dcache_req_tmp_if.addr),
				.core_req_data(dcache_req_tmp_if.data),
				.core_req_tag(dcache_req_tmp_if.tag),
				.core_req_ready(dcache_req_tmp_if.ready),
				.core_rsp_valid(dcache_rsp_tmp_if.valid),
				.core_rsp_tmask(dcache_rsp_tmp_if.tmask),
				.core_rsp_data(dcache_rsp_tmp_if.data),
				.core_rsp_tag(dcache_rsp_tmp_if.tag),
				.core_rsp_ready(dcache_rsp_tmp_if.ready),
				.mem_req_valid(dcache_mem_req_if.valid),
				.mem_req_rw(dcache_mem_req_if.rw),
				.mem_req_byteen(dcache_mem_req_if.byteen),
				.mem_req_addr(dcache_mem_req_if.addr),
				.mem_req_data(dcache_mem_req_if.data),
				.mem_req_tag(dcache_mem_req_if.tag),
				.mem_req_ready(dcache_mem_req_if.ready),
				.mem_rsp_valid(dcache_mem_rsp_if.valid),
				.mem_rsp_data(dcache_mem_rsp_if.data),
				.mem_rsp_tag(dcache_mem_rsp_if.tag),
				.mem_rsp_ready(dcache_mem_rsp_if.ready)
			);
			// Trace: ../../rtl/VX_mem_unit.sv:188:5
			if (1) begin : genblk1
				// Trace: ../../rtl/VX_mem_unit.sv:189:9
				// expanded interface instance: smem_req_if
				localparam _param_C3EC4_NUM_REQS = 2;
				localparam _param_C3EC4_WORD_SIZE = 4;
				localparam _param_C3EC4_TAG_WIDTH = 47;
				if (1) begin : smem_req_if
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:7:15
					localparam NUM_REQS = _param_C3EC4_NUM_REQS;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:8:15
					localparam WORD_SIZE = _param_C3EC4_WORD_SIZE;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:9:15
					localparam TAG_WIDTH = _param_C3EC4_TAG_WIDTH;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:12:5
					wire [1:0] valid;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:13:5
					wire [1:0] rw;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:14:5
					wire [7:0] byteen;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:15:5
					wire [59:0] addr;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:16:5
					wire [63:0] data;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:17:5
					wire [93:0] tag;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:18:5
					wire [1:0] ready;
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:20:5
					// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:30:5
				end
				// Trace: ../../rtl/VX_mem_unit.sv:195:9
				// expanded interface instance: smem_rsp_if
				localparam _param_541C4_NUM_REQS = 2;
				localparam _param_541C4_WORD_SIZE = 4;
				localparam _param_541C4_TAG_WIDTH = 47;
				if (1) begin : smem_rsp_if
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:7:15
					localparam NUM_REQS = _param_541C4_NUM_REQS;
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:8:15
					localparam WORD_SIZE = _param_541C4_WORD_SIZE;
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:9:15
					localparam TAG_WIDTH = _param_541C4_TAG_WIDTH;
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:12:5
					wire valid;
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:13:5
					wire [1:0] tmask;
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:14:5
					wire [63:0] data;
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:15:5
					wire [46:0] tag;
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:16:5
					wire ready;
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:18:5
					// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:26:5
				end
				// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:201:31
				wire smem_arb_reset;
				// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:201:64
				VX_reset_relay __smem_arb_reset(
					.clk(clk),
					.reset(reset),
					.reset_o(smem_arb_reset)
				);
				// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:202:27
				wire smem_reset;
				// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_mem_unit.sv:202:60
				VX_reset_relay __smem_reset(
					.clk(clk),
					.reset(reset),
					.reset_o(smem_reset)
				);
				// Trace: ../../rtl/VX_mem_unit.sv:204:9
				VX_smem_arb #(
					.NUM_REQS(2),
					.LANES(2),
					.DATA_SIZE(4),
					.TAG_IN_WIDTH(48),
					.TAG_SEL_IDX(0),
					.TYPE("P"),
					.BUFFERED_REQ(2),
					.BUFFERED_RSP(1)
				) smem_arb(
					.clk(clk),
					.reset(smem_arb_reset),
					.req_valid_in(VX_core.dcache_req_if.valid),
					.req_rw_in(VX_core.dcache_req_if.rw),
					.req_byteen_in(VX_core.dcache_req_if.byteen),
					.req_addr_in(VX_core.dcache_req_if.addr),
					.req_data_in(VX_core.dcache_req_if.data),
					.req_tag_in(VX_core.dcache_req_if.tag),
					.req_ready_in(VX_core.dcache_req_if.ready),
					.req_valid_out({smem_req_if.valid, dcache_req_tmp_if.valid}),
					.req_rw_out({smem_req_if.rw, dcache_req_tmp_if.rw}),
					.req_byteen_out({smem_req_if.byteen, dcache_req_tmp_if.byteen}),
					.req_addr_out({smem_req_if.addr, dcache_req_tmp_if.addr}),
					.req_data_out({smem_req_if.data, dcache_req_tmp_if.data}),
					.req_tag_out({smem_req_if.tag, dcache_req_tmp_if.tag}),
					.req_ready_out({smem_req_if.ready, dcache_req_tmp_if.ready}),
					.rsp_valid_in({smem_rsp_if.valid, dcache_rsp_tmp_if.valid}),
					.rsp_tmask_in({smem_rsp_if.tmask, dcache_rsp_tmp_if.tmask}),
					.rsp_data_in({smem_rsp_if.data, dcache_rsp_tmp_if.data}),
					.rsp_tag_in({smem_rsp_if.tag, dcache_rsp_tmp_if.tag}),
					.rsp_ready_in({smem_rsp_if.ready, dcache_rsp_tmp_if.ready}),
					.rsp_valid_out(VX_core.dcache_rsp_if.valid),
					.rsp_tmask_out(VX_core.dcache_rsp_if.tmask),
					.rsp_tag_out(VX_core.dcache_rsp_if.tag),
					.rsp_data_out(VX_core.dcache_rsp_if.data),
					.rsp_ready_out(VX_core.dcache_rsp_if.ready)
				);
				// Trace: ../../rtl/VX_mem_unit.sv:250:9
				VX_shared_mem #(
					.CACHE_ID((0 + (CORE_ID * 3)) + 2),
					.CACHE_SIZE(4096),
					.NUM_BANKS(2),
					.WORD_SIZE(4),
					.NUM_REQS(2),
					.CREQ_SIZE(2),
					.CRSQ_SIZE(2),
					.CORE_TAG_WIDTH(47),
					.CORE_TAG_ID_BITS(3),
					.BANK_ADDR_OFFSET(8)
				) smem(
					.clk(clk),
					.reset(smem_reset),
					.core_req_valid(smem_req_if.valid),
					.core_req_rw(smem_req_if.rw),
					.core_req_byteen(smem_req_if.byteen),
					.core_req_addr(smem_req_if.addr),
					.core_req_data(smem_req_if.data),
					.core_req_tag(smem_req_if.tag),
					.core_req_ready(smem_req_if.ready),
					.core_rsp_valid(smem_rsp_if.valid),
					.core_rsp_tmask(smem_rsp_if.tmask),
					.core_rsp_data(smem_rsp_if.data),
					.core_rsp_tag(smem_rsp_if.tag),
					.core_rsp_ready(smem_rsp_if.ready)
				);
			end
			// Trace: ../../rtl/VX_mem_unit.sv:310:5
			wire [(4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) - 1:0] icache_mem_req_tag = sv2v_cast_7CD18(icache_mem_req_if.tag);
			// Trace: ../../rtl/VX_mem_unit.sv:311:5
			wire [(4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) - 1:0] icache_mem_rsp_tag;
			// Trace: ../../rtl/VX_mem_unit.sv:312:5
			assign icache_mem_rsp_if.tag = icache_mem_rsp_tag[0:0];
			// Trace: ../../rtl/VX_mem_unit.sv:315:5
			VX_mem_arb #(
				.NUM_REQS(2),
				.DATA_WIDTH((0 || 0 ? 16 : 64) * 8),
				.ADDR_WIDTH(32 - $clog2((0 || 0 ? 16 : 64))),
				.TAG_IN_WIDTH((4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)),
				.TYPE("R"),
				.TAG_SEL_IDX(1),
				.BUFFERED_REQ(1),
				.BUFFERED_RSP(2)
			) mem_arb(
				.clk(clk),
				.reset(mem_arb_reset),
				.req_valid_in({dcache_mem_req_if.valid, icache_mem_req_if.valid}),
				.req_rw_in({dcache_mem_req_if.rw, icache_mem_req_if.rw}),
				.req_byteen_in({dcache_mem_req_if.byteen, icache_mem_req_if.byteen}),
				.req_addr_in({dcache_mem_req_if.addr, icache_mem_req_if.addr}),
				.req_data_in({dcache_mem_req_if.data, icache_mem_req_if.data}),
				.req_tag_in({dcache_mem_req_if.tag, icache_mem_req_tag}),
				.req_ready_in({dcache_mem_req_if.ready, icache_mem_req_if.ready}),
				.req_valid_out(VX_core.mem_req_if.valid),
				.req_rw_out(VX_core.mem_req_if.rw),
				.req_byteen_out(VX_core.mem_req_if.byteen),
				.req_addr_out(VX_core.mem_req_if.addr),
				.req_data_out(VX_core.mem_req_if.data),
				.req_tag_out(VX_core.mem_req_if.tag),
				.req_ready_out(VX_core.mem_req_if.ready),
				.rsp_valid_out({dcache_mem_rsp_if.valid, icache_mem_rsp_if.valid}),
				.rsp_data_out({dcache_mem_rsp_if.data, icache_mem_rsp_if.data}),
				.rsp_tag_out({dcache_mem_rsp_if.tag, icache_mem_rsp_tag}),
				.rsp_ready_out({dcache_mem_rsp_if.ready, icache_mem_rsp_if.ready}),
				.rsp_valid_in(VX_core.mem_rsp_if.valid),
				.rsp_tag_in(VX_core.mem_rsp_if.tag),
				.rsp_data_in(VX_core.mem_rsp_if.data),
				.rsp_ready_in(VX_core.mem_rsp_if.ready)
			);
		end
	endgenerate
	assign mem_unit.clk = clk;
	assign mem_unit.reset = reset;
endmodule
// removed module with interface ports: VX_csr_data
// removed module with interface ports: VX_csr_unit
// removed module with interface ports: VX_decode
// removed module with interface ports: VX_dispatch
// removed module with interface ports: VX_execute
// removed module with interface ports: VX_fetch
// removed module with interface ports: VX_fpu_unit
// removed module with interface ports: VX_gpr_stage
// removed module with interface ports: VX_gpu_unit
// removed module with interface ports: VX_ibuffer
// removed module with interface ports: VX_icache_stage
module VX_ipdom_stack (
	clk,
	reset,
	pair,
	q1,
	q2,
	d,
	push,
	pop,
	index,
	empty,
	full
);
	// Trace: ../../rtl/VX_ipdom_stack.sv:4:15
	parameter WIDTH = 1;
	// Trace: ../../rtl/VX_ipdom_stack.sv:5:15
	parameter DEPTH = 1;
	// Trace: ../../rtl/VX_ipdom_stack.sv:7:5
	input wire clk;
	// Trace: ../../rtl/VX_ipdom_stack.sv:8:5
	input wire reset;
	// Trace: ../../rtl/VX_ipdom_stack.sv:9:5
	input wire pair;
	// Trace: ../../rtl/VX_ipdom_stack.sv:10:5
	input wire [WIDTH - 1:0] q1;
	// Trace: ../../rtl/VX_ipdom_stack.sv:11:5
	input wire [WIDTH - 1:0] q2;
	// Trace: ../../rtl/VX_ipdom_stack.sv:12:5
	output wire [WIDTH - 1:0] d;
	// Trace: ../../rtl/VX_ipdom_stack.sv:13:5
	input wire push;
	// Trace: ../../rtl/VX_ipdom_stack.sv:14:5
	input wire pop;
	// Trace: ../../rtl/VX_ipdom_stack.sv:15:5
	output wire index;
	// Trace: ../../rtl/VX_ipdom_stack.sv:16:5
	output wire empty;
	// Trace: ../../rtl/VX_ipdom_stack.sv:17:5
	output wire full;
	// Trace: ../../rtl/VX_ipdom_stack.sv:19:5
	localparam ADDRW = $clog2(DEPTH);
	// Trace: ../../rtl/VX_ipdom_stack.sv:21:5
	reg is_part [DEPTH - 1:0];
	// Trace: ../../rtl/VX_ipdom_stack.sv:23:5
	reg [ADDRW - 1:0] rd_ptr;
	reg [ADDRW - 1:0] wr_ptr;
	// Trace: ../../rtl/VX_ipdom_stack.sv:25:5
	wire [WIDTH - 1:0] d1;
	wire [WIDTH - 1:0] d2;
	// Trace: ../../rtl/VX_ipdom_stack.sv:27:5
	function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
		input reg signed [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D_signed = inp;
	endfunction
	function automatic [ADDRW - 1:0] sv2v_cast_8BB5D;
		input reg [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D = inp;
	endfunction
	always @(posedge clk)
		// Trace: ../../rtl/VX_ipdom_stack.sv:28:9
		if (reset) begin
			// Trace: ../../rtl/VX_ipdom_stack.sv:29:13
			rd_ptr <= 0;
			// Trace: ../../rtl/VX_ipdom_stack.sv:30:13
			wr_ptr <= 0;
		end
		else
			// Trace: ../../rtl/VX_ipdom_stack.sv:32:13
			if (push) begin
				// Trace: ../../rtl/VX_ipdom_stack.sv:33:17
				rd_ptr <= wr_ptr;
				// Trace: ../../rtl/VX_ipdom_stack.sv:34:17
				wr_ptr <= wr_ptr + sv2v_cast_8BB5D_signed(1);
			end
			else if (pop) begin
				// Trace: ../../rtl/VX_ipdom_stack.sv:36:17
				wr_ptr <= wr_ptr - sv2v_cast_8BB5D(is_part[rd_ptr]);
				// Trace: ../../rtl/VX_ipdom_stack.sv:37:17
				rd_ptr <= rd_ptr - sv2v_cast_8BB5D(is_part[rd_ptr]);
			end
	// Trace: ../../rtl/VX_ipdom_stack.sv:42:5
	VX_dp_ram #(
		.DATAW(WIDTH * 2),
		.SIZE(DEPTH),
		.LUTRAM(1)
	) store(
		.clk(clk),
		.wren(push),
		.waddr(wr_ptr),
		.wdata({q2, q1}),
		.raddr(rd_ptr),
		.rdata({d2, d1})
	);
	// Trace: ../../rtl/VX_ipdom_stack.sv:55:5
	always @(posedge clk)
		// Trace: ../../rtl/VX_ipdom_stack.sv:56:9
		if (push)
			// Trace: ../../rtl/VX_ipdom_stack.sv:57:13
			is_part[wr_ptr] <= ~pair;
		else if (pop)
			// Trace: ../../rtl/VX_ipdom_stack.sv:59:13
			is_part[rd_ptr] <= 1;
	// Trace: ../../rtl/VX_ipdom_stack.sv:63:5
	assign index = is_part[rd_ptr];
	// Trace: ../../rtl/VX_ipdom_stack.sv:64:5
	assign d = (index ? d1 : d2);
	// Trace: ../../rtl/VX_ipdom_stack.sv:65:5
	assign empty = sv2v_cast_8BB5D_signed(0) == wr_ptr;
	// Trace: ../../rtl/VX_ipdom_stack.sv:66:5
	assign full = sv2v_cast_8BB5D_signed(DEPTH - 1) == wr_ptr;
endmodule
// removed module with interface ports: VX_issue
// removed module with interface ports: VX_lsu_unit
module VX_mem_arb (
	clk,
	reset,
	req_valid_in,
	req_tag_in,
	req_addr_in,
	req_rw_in,
	req_byteen_in,
	req_data_in,
	req_ready_in,
	req_valid_out,
	req_tag_out,
	req_addr_out,
	req_rw_out,
	req_byteen_out,
	req_data_out,
	req_ready_out,
	rsp_valid_in,
	rsp_tag_in,
	rsp_data_in,
	rsp_ready_in,
	rsp_valid_out,
	rsp_tag_out,
	rsp_data_out,
	rsp_ready_out
);
	// Trace: ../../rtl/VX_mem_arb.sv:4:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/VX_mem_arb.sv:5:15
	parameter DATA_WIDTH = 1;
	// Trace: ../../rtl/VX_mem_arb.sv:6:15
	parameter ADDR_WIDTH = 1;
	// Trace: ../../rtl/VX_mem_arb.sv:7:15
	parameter TAG_IN_WIDTH = 1;
	// Trace: ../../rtl/VX_mem_arb.sv:8:15
	parameter TAG_SEL_IDX = 0;
	// Trace: ../../rtl/VX_mem_arb.sv:9:15
	parameter BUFFERED_REQ = 0;
	// Trace: ../../rtl/VX_mem_arb.sv:10:15
	parameter BUFFERED_RSP = 0;
	// Trace: ../../rtl/VX_mem_arb.sv:11:15
	parameter TYPE = "P";
	// Trace: ../../rtl/VX_mem_arb.sv:13:15
	parameter DATA_SIZE = DATA_WIDTH / 8;
	// Trace: ../../rtl/VX_mem_arb.sv:14:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: ../../rtl/VX_mem_arb.sv:15:15
	parameter TAG_OUT_WIDTH = TAG_IN_WIDTH + LOG_NUM_REQS;
	// Trace: ../../rtl/VX_mem_arb.sv:17:5
	input wire clk;
	// Trace: ../../rtl/VX_mem_arb.sv:18:5
	input wire reset;
	// Trace: ../../rtl/VX_mem_arb.sv:21:5
	input wire [NUM_REQS - 1:0] req_valid_in;
	// Trace: ../../rtl/VX_mem_arb.sv:22:5
	input wire [(NUM_REQS * TAG_IN_WIDTH) - 1:0] req_tag_in;
	// Trace: ../../rtl/VX_mem_arb.sv:23:5
	input wire [(NUM_REQS * ADDR_WIDTH) - 1:0] req_addr_in;
	// Trace: ../../rtl/VX_mem_arb.sv:24:5
	input wire [NUM_REQS - 1:0] req_rw_in;
	// Trace: ../../rtl/VX_mem_arb.sv:25:5
	input wire [(NUM_REQS * DATA_SIZE) - 1:0] req_byteen_in;
	// Trace: ../../rtl/VX_mem_arb.sv:26:5
	input wire [(NUM_REQS * DATA_WIDTH) - 1:0] req_data_in;
	// Trace: ../../rtl/VX_mem_arb.sv:27:5
	output wire [NUM_REQS - 1:0] req_ready_in;
	// Trace: ../../rtl/VX_mem_arb.sv:30:5
	output wire req_valid_out;
	// Trace: ../../rtl/VX_mem_arb.sv:31:5
	output wire [TAG_OUT_WIDTH - 1:0] req_tag_out;
	// Trace: ../../rtl/VX_mem_arb.sv:32:5
	output wire [ADDR_WIDTH - 1:0] req_addr_out;
	// Trace: ../../rtl/VX_mem_arb.sv:33:5
	output wire req_rw_out;
	// Trace: ../../rtl/VX_mem_arb.sv:34:5
	output wire [DATA_SIZE - 1:0] req_byteen_out;
	// Trace: ../../rtl/VX_mem_arb.sv:35:5
	output wire [DATA_WIDTH - 1:0] req_data_out;
	// Trace: ../../rtl/VX_mem_arb.sv:36:5
	input wire req_ready_out;
	// Trace: ../../rtl/VX_mem_arb.sv:39:5
	input wire rsp_valid_in;
	// Trace: ../../rtl/VX_mem_arb.sv:40:5
	input wire [TAG_OUT_WIDTH - 1:0] rsp_tag_in;
	// Trace: ../../rtl/VX_mem_arb.sv:41:5
	input wire [DATA_WIDTH - 1:0] rsp_data_in;
	// Trace: ../../rtl/VX_mem_arb.sv:42:5
	output wire rsp_ready_in;
	// Trace: ../../rtl/VX_mem_arb.sv:45:5
	output wire [NUM_REQS - 1:0] rsp_valid_out;
	// Trace: ../../rtl/VX_mem_arb.sv:46:5
	output wire [(NUM_REQS * TAG_IN_WIDTH) - 1:0] rsp_tag_out;
	// Trace: ../../rtl/VX_mem_arb.sv:47:5
	output wire [(NUM_REQS * DATA_WIDTH) - 1:0] rsp_data_out;
	// Trace: ../../rtl/VX_mem_arb.sv:48:5
	input wire [NUM_REQS - 1:0] rsp_ready_out;
	// Trace: ../../rtl/VX_mem_arb.sv:50:5
	localparam REQ_DATAW = (((TAG_OUT_WIDTH + ADDR_WIDTH) + 1) + DATA_SIZE) + DATA_WIDTH;
	// Trace: ../../rtl/VX_mem_arb.sv:51:5
	localparam RSP_DATAW = TAG_IN_WIDTH + DATA_WIDTH;
	// Trace: ../../rtl/VX_mem_arb.sv:53:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_REQS > 1) begin : genblk1
			// Trace: ../../rtl/VX_mem_arb.sv:55:9
			wire [(NUM_REQS * REQ_DATAW) - 1:0] req_data_in_merged;
			genvar i;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
				// Trace: ../../rtl/VX_mem_arb.sv:58:13
				wire [TAG_OUT_WIDTH - 1:0] req_tag_in_w;
				// Trace: ../../rtl/VX_mem_arb.sv:60:13
				VX_bits_insert #(
					.N(TAG_IN_WIDTH),
					.S(LOG_NUM_REQS),
					.POS(TAG_SEL_IDX)
				) bits_insert(
					.data_in(req_tag_in[i * TAG_IN_WIDTH+:TAG_IN_WIDTH]),
					.sel_in(sv2v_cast_76B5F_signed(i)),
					.data_out(req_tag_in_w)
				);
				// Trace: ../../rtl/VX_mem_arb.sv:70:13
				assign req_data_in_merged[i * REQ_DATAW+:REQ_DATAW] = {req_tag_in_w, req_addr_in[i * ADDR_WIDTH+:ADDR_WIDTH], req_rw_in[i], req_byteen_in[i * DATA_SIZE+:DATA_SIZE], req_data_in[i * DATA_WIDTH+:DATA_WIDTH]};
			end
			// Trace: ../../rtl/VX_mem_arb.sv:73:9
			VX_stream_arbiter #(
				.NUM_REQS(NUM_REQS),
				.DATAW(REQ_DATAW),
				.BUFFERED(BUFFERED_REQ),
				.TYPE(TYPE)
			) req_arb(
				.clk(clk),
				.reset(reset),
				.valid_in(req_valid_in),
				.data_in(req_data_in_merged),
				.ready_in(req_ready_in),
				.valid_out(req_valid_out),
				.data_out({req_tag_out, req_addr_out, req_rw_out, req_byteen_out, req_data_out}),
				.ready_out(req_ready_out)
			);
			// Trace: ../../rtl/VX_mem_arb.sv:91:9
			wire [(NUM_REQS * RSP_DATAW) - 1:0] rsp_data_out_merged;
			// Trace: ../../rtl/VX_mem_arb.sv:93:9
			wire [LOG_NUM_REQS - 1:0] rsp_sel = rsp_tag_in[TAG_SEL_IDX+:LOG_NUM_REQS];
			// Trace: ../../rtl/VX_mem_arb.sv:95:9
			wire [TAG_IN_WIDTH - 1:0] rsp_tag_in_w;
			// Trace: ../../rtl/VX_mem_arb.sv:97:9
			VX_bits_remove #(
				.N(TAG_OUT_WIDTH),
				.S(LOG_NUM_REQS),
				.POS(TAG_SEL_IDX)
			) bits_remove(
				.data_in(rsp_tag_in),
				.data_out(rsp_tag_in_w)
			);
			// Trace: ../../rtl/VX_mem_arb.sv:106:9
			VX_stream_demux #(
				.NUM_REQS(NUM_REQS),
				.DATAW(RSP_DATAW),
				.BUFFERED(BUFFERED_RSP)
			) rsp_demux(
				.clk(clk),
				.reset(reset),
				.sel_in(rsp_sel),
				.valid_in(rsp_valid_in),
				.data_in({rsp_tag_in_w, rsp_data_in}),
				.ready_in(rsp_ready_in),
				.valid_out(rsp_valid_out),
				.data_out(rsp_data_out_merged),
				.ready_out(rsp_ready_out)
			);
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk2
				// Trace: ../../rtl/VX_mem_arb.sv:123:13
				assign {rsp_tag_out[i * TAG_IN_WIDTH+:TAG_IN_WIDTH], rsp_data_out[i * DATA_WIDTH+:DATA_WIDTH]} = rsp_data_out_merged[i * RSP_DATAW+:RSP_DATAW];
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/VX_mem_arb.sv:131:9
			assign req_valid_out = req_valid_in;
			// Trace: ../../rtl/VX_mem_arb.sv:132:9
			assign req_tag_out = req_tag_in;
			// Trace: ../../rtl/VX_mem_arb.sv:133:9
			assign req_addr_out = req_addr_in;
			// Trace: ../../rtl/VX_mem_arb.sv:134:9
			assign req_rw_out = req_rw_in;
			// Trace: ../../rtl/VX_mem_arb.sv:135:9
			assign req_byteen_out = req_byteen_in;
			// Trace: ../../rtl/VX_mem_arb.sv:136:9
			assign req_data_out = req_data_in;
			// Trace: ../../rtl/VX_mem_arb.sv:137:9
			assign req_ready_in = req_ready_out;
			// Trace: ../../rtl/VX_mem_arb.sv:139:9
			assign rsp_valid_out = rsp_valid_in;
			// Trace: ../../rtl/VX_mem_arb.sv:140:9
			assign rsp_tag_out = rsp_tag_in;
			// Trace: ../../rtl/VX_mem_arb.sv:141:9
			assign rsp_data_out = rsp_data_in;
			// Trace: ../../rtl/VX_mem_arb.sv:142:9
			assign rsp_ready_in = rsp_ready_out;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_mem_unit
module VX_muldiv (
	clk,
	reset,
	alu_op,
	uuid_in,
	wid_in,
	tmask_in,
	PC_in,
	rd_in,
	wb_in,
	alu_in1,
	alu_in2,
	uuid_out,
	wid_out,
	tmask_out,
	PC_out,
	rd_out,
	wb_out,
	data_out,
	valid_in,
	ready_in,
	valid_out,
	ready_out
);
	// Trace: ../../rtl/VX_muldiv.sv:4:5
	input wire clk;
	// Trace: ../../rtl/VX_muldiv.sv:5:5
	input wire reset;
	// Trace: ../../rtl/VX_muldiv.sv:8:5
	input wire [2:0] alu_op;
	// Trace: ../../rtl/VX_muldiv.sv:9:5
	input wire [43:0] uuid_in;
	// Trace: ../../rtl/VX_muldiv.sv:10:5
	input wire [0:0] wid_in;
	// Trace: ../../rtl/VX_muldiv.sv:11:5
	input wire [1:0] tmask_in;
	// Trace: ../../rtl/VX_muldiv.sv:12:5
	input wire [31:0] PC_in;
	// Trace: ../../rtl/VX_muldiv.sv:13:5
	input wire [4:0] rd_in;
	// Trace: ../../rtl/VX_muldiv.sv:14:5
	input wire wb_in;
	// Trace: ../../rtl/VX_muldiv.sv:15:5
	input wire [63:0] alu_in1;
	// Trace: ../../rtl/VX_muldiv.sv:16:5
	input wire [63:0] alu_in2;
	// Trace: ../../rtl/VX_muldiv.sv:19:5
	output wire [43:0] uuid_out;
	// Trace: ../../rtl/VX_muldiv.sv:20:5
	output wire [0:0] wid_out;
	// Trace: ../../rtl/VX_muldiv.sv:21:5
	output wire [1:0] tmask_out;
	// Trace: ../../rtl/VX_muldiv.sv:22:5
	output wire [31:0] PC_out;
	// Trace: ../../rtl/VX_muldiv.sv:23:5
	output wire [4:0] rd_out;
	// Trace: ../../rtl/VX_muldiv.sv:24:5
	output wire wb_out;
	// Trace: ../../rtl/VX_muldiv.sv:25:5
	output wire [63:0] data_out;
	// Trace: ../../rtl/VX_muldiv.sv:28:5
	input wire valid_in;
	// Trace: ../../rtl/VX_muldiv.sv:29:5
	output wire ready_in;
	// Trace: ../../rtl/VX_muldiv.sv:30:5
	output wire valid_out;
	// Trace: ../../rtl/VX_muldiv.sv:31:5
	input wire ready_out;
	// Trace: ../../rtl/VX_muldiv.sv:34:5
	wire is_div_op = alu_op[2];
	// Trace: ../../rtl/VX_muldiv.sv:36:5
	wire [63:0] mul_result;
	// Trace: ../../rtl/VX_muldiv.sv:37:5
	wire [43:0] mul_uuid_out;
	// Trace: ../../rtl/VX_muldiv.sv:38:5
	wire [0:0] mul_wid_out;
	// Trace: ../../rtl/VX_muldiv.sv:39:5
	wire [1:0] mul_tmask_out;
	// Trace: ../../rtl/VX_muldiv.sv:40:5
	wire [31:0] mul_PC_out;
	// Trace: ../../rtl/VX_muldiv.sv:41:5
	wire [4:0] mul_rd_out;
	// Trace: ../../rtl/VX_muldiv.sv:42:5
	wire mul_wb_out;
	// Trace: ../../rtl/VX_muldiv.sv:44:5
	wire stall_out;
	// Trace: ../../rtl/VX_muldiv.sv:46:5
	wire mul_valid_out;
	// Trace: ../../rtl/VX_muldiv.sv:47:5
	wire mul_valid_in = valid_in && !is_div_op;
	// Trace: ../../rtl/VX_muldiv.sv:48:5
	wire mul_ready_in = ~stall_out || ~mul_valid_out;
	// Trace: ../../rtl/VX_muldiv.sv:50:5
	wire is_mulh_in = alu_op != 3'h0;
	// Trace: ../../rtl/VX_muldiv.sv:51:5
	wire is_signed_mul_a = alu_op != 3'h3;
	// Trace: ../../rtl/VX_muldiv.sv:52:5
	wire is_signed_mul_b = (alu_op != 3'h3) && (alu_op != 3'h2);
	// Trace: ../../rtl/VX_muldiv.sv:82:5
	wire is_mulh_out;
	// Trace: ../../rtl/VX_muldiv.sv:84:5
	genvar i;
	generate
		for (i = 0; i < 2; i = i + 1) begin : genblk1
			// Trace: ../../rtl/VX_muldiv.sv:85:9
			wire [32:0] mul_in1 = {is_signed_mul_a & alu_in1[(i * 32) + 31], alu_in1[i * 32+:32]};
			// Trace: ../../rtl/VX_muldiv.sv:86:9
			wire [32:0] mul_in2 = {is_signed_mul_b & alu_in2[(i * 32) + 31], alu_in2[i * 32+:32]};
			// Trace: ../../rtl/VX_muldiv.sv:88:9
			wire [65:0] mul_result_tmp;
			// Trace: ../../rtl/VX_muldiv.sv:91:9
			VX_multiplier #(
				.WIDTHA(33),
				.WIDTHB(33),
				.WIDTHP(66),
				.SIGNED(1),
				.LATENCY(3)
			) multiplier(
				.clk(clk),
				.enable(mul_ready_in),
				.dataa(mul_in1),
				.datab(mul_in2),
				.result(mul_result_tmp)
			);
			// Trace: ../../rtl/VX_muldiv.sv:105:9
			assign mul_result[i * 32+:32] = (is_mulh_out ? mul_result_tmp[63:32] : mul_result_tmp[31:0]);
		end
	endgenerate
	// Trace: ../../rtl/VX_muldiv.sv:108:5
	VX_shift_register #(
		.DATAW(87),
		.DEPTH(3),
		.RESETW(1)
	) mul_shift_reg(
		.clk(clk),
		.reset(reset),
		.enable(mul_ready_in),
		.data_in({mul_valid_in, uuid_in, wid_in, tmask_in, PC_in, rd_in, wb_in, is_mulh_in}),
		.data_out({mul_valid_out, mul_uuid_out, mul_wid_out, mul_tmask_out, mul_PC_out, mul_rd_out, mul_wb_out, is_mulh_out})
	);
	// Trace: ../../rtl/VX_muldiv.sv:124:5
	wire [63:0] div_result;
	// Trace: ../../rtl/VX_muldiv.sv:125:5
	wire [43:0] div_uuid_out;
	// Trace: ../../rtl/VX_muldiv.sv:126:5
	wire [0:0] div_wid_out;
	// Trace: ../../rtl/VX_muldiv.sv:127:5
	wire [1:0] div_tmask_out;
	// Trace: ../../rtl/VX_muldiv.sv:128:5
	wire [31:0] div_PC_out;
	// Trace: ../../rtl/VX_muldiv.sv:129:5
	wire [4:0] div_rd_out;
	// Trace: ../../rtl/VX_muldiv.sv:130:5
	wire div_wb_out;
	// Trace: ../../rtl/VX_muldiv.sv:132:5
	wire is_rem_op_in = (alu_op == 3'h6) || (alu_op == 3'h7);
	// Trace: ../../rtl/VX_muldiv.sv:133:5
	wire is_signed_div = (alu_op == 3'h4) || (alu_op == 3'h6);
	// Trace: ../../rtl/VX_muldiv.sv:134:5
	wire div_valid_in = valid_in && is_div_op;
	// Trace: ../../rtl/VX_muldiv.sv:135:5
	wire div_ready_out = ~stall_out && ~mul_valid_out;
	// Trace: ../../rtl/VX_muldiv.sv:136:5
	wire div_ready_in;
	// Trace: ../../rtl/VX_muldiv.sv:137:5
	wire div_valid_out;
	// Trace: ../../rtl/VX_muldiv.sv:169:5
	wire [63:0] div_result_tmp;
	wire [63:0] rem_result_tmp;
	// Trace: ../../rtl/VX_muldiv.sv:170:5
	wire is_rem_op_out;
	// Trace: ../../rtl/VX_muldiv.sv:172:5
	VX_serial_div #(
		.WIDTHN(32),
		.WIDTHD(32),
		.WIDTHQ(32),
		.WIDTHR(32),
		.LANES(2),
		.TAGW(106)
	) divide(
		.clk(clk),
		.reset(reset),
		.valid_in(div_valid_in),
		.ready_in(div_ready_in),
		.signed_mode(is_signed_div),
		.tag_in({uuid_in, wid_in, tmask_in, PC_in, rd_in, wb_in, is_rem_op_in}),
		.numer(alu_in1),
		.denom(alu_in2),
		.quotient(div_result_tmp),
		.remainder(rem_result_tmp),
		.ready_out(div_ready_out),
		.valid_out(div_valid_out),
		.tag_out({div_uuid_out, div_wid_out, div_tmask_out, div_PC_out, div_rd_out, div_wb_out, is_rem_op_out})
	);
	// Trace: ../../rtl/VX_muldiv.sv:195:5
	assign div_result = (is_rem_op_out ? rem_result_tmp : div_result_tmp);
	// Trace: ../../rtl/VX_muldiv.sv:201:5
	wire rsp_valid = mul_valid_out || div_valid_out;
	// Trace: ../../rtl/VX_muldiv.sv:202:5
	wire [43:0] rsp_uuid = (mul_valid_out ? mul_uuid_out : div_uuid_out);
	// Trace: ../../rtl/VX_muldiv.sv:203:5
	wire [0:0] rsp_wid = (mul_valid_out ? mul_wid_out : div_wid_out);
	// Trace: ../../rtl/VX_muldiv.sv:204:5
	wire [1:0] rsp_tmask = (mul_valid_out ? mul_tmask_out : div_tmask_out);
	// Trace: ../../rtl/VX_muldiv.sv:205:5
	wire [31:0] rsp_PC = (mul_valid_out ? mul_PC_out : div_PC_out);
	// Trace: ../../rtl/VX_muldiv.sv:206:5
	wire [4:0] rsp_rd = (mul_valid_out ? mul_rd_out : div_rd_out);
	// Trace: ../../rtl/VX_muldiv.sv:207:5
	wire rsp_wb = (mul_valid_out ? mul_wb_out : div_wb_out);
	// Trace: ../../rtl/VX_muldiv.sv:208:5
	wire [63:0] rsp_data = (mul_valid_out ? mul_result : div_result);
	// Trace: ../../rtl/VX_muldiv.sv:210:5
	assign stall_out = ~ready_out && valid_out;
	// Trace: ../../rtl/VX_muldiv.sv:212:5
	VX_pipe_register #(
		.DATAW(150),
		.RESETW(1)
	) pipe_reg(
		.clk(clk),
		.reset(reset),
		.enable(~stall_out),
		.data_in({rsp_valid, rsp_uuid, rsp_wid, rsp_tmask, rsp_PC, rsp_rd, rsp_wb, rsp_data}),
		.data_out({valid_out, uuid_out, wid_out, tmask_out, PC_out, rd_out, wb_out, data_out})
	);
	// Trace: ../../rtl/VX_muldiv.sv:224:5
	assign ready_in = (is_div_op ? div_ready_in : mul_ready_in);
endmodule
module VX_pipeline (
	clk,
	reset,
	dcache_req_valid,
	dcache_req_rw,
	dcache_req_byteen,
	dcache_req_addr,
	dcache_req_data,
	dcache_req_tag,
	dcache_req_ready,
	dcache_rsp_valid,
	dcache_rsp_tmask,
	dcache_rsp_data,
	dcache_rsp_tag,
	dcache_rsp_ready,
	icache_req_valid,
	icache_req_addr,
	icache_req_tag,
	icache_req_ready,
	icache_rsp_valid,
	icache_rsp_data,
	icache_rsp_tag,
	icache_rsp_ready,
	busy
);
	// Trace: ../../rtl/VX_pipeline.sv:4:15
	parameter CORE_ID = 0;
	// Trace: ../../rtl/VX_pipeline.sv:9:5
	input wire clk;
	// Trace: ../../rtl/VX_pipeline.sv:10:5
	input wire reset;
	// Trace: ../../rtl/VX_pipeline.sv:13:5
	output wire [1:0] dcache_req_valid;
	// Trace: ../../rtl/VX_pipeline.sv:14:5
	output wire [1:0] dcache_req_rw;
	// Trace: ../../rtl/VX_pipeline.sv:15:5
	output wire [7:0] dcache_req_byteen;
	// Trace: ../../rtl/VX_pipeline.sv:16:5
	output wire [59:0] dcache_req_addr;
	// Trace: ../../rtl/VX_pipeline.sv:17:5
	output wire [63:0] dcache_req_data;
	// Trace: ../../rtl/VX_pipeline.sv:18:5
	output wire [95:0] dcache_req_tag;
	// Trace: ../../rtl/VX_pipeline.sv:19:5
	input wire [1:0] dcache_req_ready;
	// Trace: ../../rtl/VX_pipeline.sv:22:5
	input wire dcache_rsp_valid;
	// Trace: ../../rtl/VX_pipeline.sv:23:5
	input wire [1:0] dcache_rsp_tmask;
	// Trace: ../../rtl/VX_pipeline.sv:24:5
	input wire [63:0] dcache_rsp_data;
	// Trace: ../../rtl/VX_pipeline.sv:25:5
	input wire [47:0] dcache_rsp_tag;
	// Trace: ../../rtl/VX_pipeline.sv:26:5
	output wire dcache_rsp_ready;
	// Trace: ../../rtl/VX_pipeline.sv:29:5
	output wire icache_req_valid;
	// Trace: ../../rtl/VX_pipeline.sv:30:5
	output wire [29:0] icache_req_addr;
	// Trace: ../../rtl/VX_pipeline.sv:31:5
	output wire [44:0] icache_req_tag;
	// Trace: ../../rtl/VX_pipeline.sv:32:5
	input wire icache_req_ready;
	// Trace: ../../rtl/VX_pipeline.sv:35:5
	input wire icache_rsp_valid;
	// Trace: ../../rtl/VX_pipeline.sv:36:5
	input wire [31:0] icache_rsp_data;
	// Trace: ../../rtl/VX_pipeline.sv:37:5
	input wire [44:0] icache_rsp_tag;
	// Trace: ../../rtl/VX_pipeline.sv:38:5
	output wire icache_rsp_ready;
	// Trace: ../../rtl/VX_pipeline.sv:45:5
	output wire busy;
	// Trace: ../../rtl/VX_pipeline.sv:51:5
	// expanded interface instance: dcache_req_if
	localparam _param_BD702_NUM_REQS = 2;
	localparam _param_BD702_WORD_SIZE = 4;
	localparam _param_BD702_TAG_WIDTH = 48;
	generate
		if (1) begin : dcache_req_if
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:7:15
			localparam NUM_REQS = _param_BD702_NUM_REQS;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:8:15
			localparam WORD_SIZE = _param_BD702_WORD_SIZE;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:9:15
			localparam TAG_WIDTH = _param_BD702_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:12:5
			wire [1:0] valid;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:13:5
			wire [1:0] rw;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:14:5
			wire [7:0] byteen;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:15:5
			wire [59:0] addr;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:16:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:17:5
			wire [95:0] tag;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:18:5
			wire [1:0] ready;
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:20:5
			// Trace: ../../rtl/interfaces/VX_dcache_req_if.sv:30:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:57:5
	assign dcache_req_valid = dcache_req_if.valid;
	// Trace: ../../rtl/VX_pipeline.sv:58:5
	assign dcache_req_rw = dcache_req_if.rw;
	// Trace: ../../rtl/VX_pipeline.sv:59:5
	assign dcache_req_byteen = dcache_req_if.byteen;
	// Trace: ../../rtl/VX_pipeline.sv:60:5
	assign dcache_req_addr = dcache_req_if.addr;
	// Trace: ../../rtl/VX_pipeline.sv:61:5
	assign dcache_req_data = dcache_req_if.data;
	// Trace: ../../rtl/VX_pipeline.sv:62:5
	assign dcache_req_tag = dcache_req_if.tag;
	// Trace: ../../rtl/VX_pipeline.sv:63:5
	assign dcache_req_if.ready = dcache_req_ready;
	// Trace: ../../rtl/VX_pipeline.sv:69:5
	// expanded interface instance: dcache_rsp_if
	localparam _param_2395E_NUM_REQS = 2;
	localparam _param_2395E_WORD_SIZE = 4;
	localparam _param_2395E_TAG_WIDTH = 48;
	generate
		if (1) begin : dcache_rsp_if
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:7:15
			localparam NUM_REQS = _param_2395E_NUM_REQS;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:8:15
			localparam WORD_SIZE = _param_2395E_WORD_SIZE;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:9:15
			localparam TAG_WIDTH = _param_2395E_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:12:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:13:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:14:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:15:5
			wire [47:0] tag;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:16:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:18:5
			// Trace: ../../rtl/interfaces/VX_dcache_rsp_if.sv:26:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:75:5
	assign dcache_rsp_if.valid = dcache_rsp_valid;
	// Trace: ../../rtl/VX_pipeline.sv:76:5
	assign dcache_rsp_if.tmask = dcache_rsp_tmask;
	// Trace: ../../rtl/VX_pipeline.sv:77:5
	assign dcache_rsp_if.data = dcache_rsp_data;
	// Trace: ../../rtl/VX_pipeline.sv:78:5
	assign dcache_rsp_if.tag = dcache_rsp_tag;
	// Trace: ../../rtl/VX_pipeline.sv:79:5
	assign dcache_rsp_ready = dcache_rsp_if.ready;
	// Trace: ../../rtl/VX_pipeline.sv:85:5
	// expanded interface instance: icache_req_if
	localparam _param_1F99A_WORD_SIZE = 4;
	localparam _param_1F99A_TAG_WIDTH = 45;
	generate
		if (1) begin : icache_req_if
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:7:15
			localparam WORD_SIZE = _param_1F99A_WORD_SIZE;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:8:15
			localparam TAG_WIDTH = _param_1F99A_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:11:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:12:5
			wire [29:0] addr;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:13:5
			wire [44:0] tag;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:14:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:16:5
			// Trace: ../../rtl/interfaces/VX_icache_req_if.sv:23:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:90:5
	assign icache_req_valid = icache_req_if.valid;
	// Trace: ../../rtl/VX_pipeline.sv:91:5
	assign icache_req_addr = icache_req_if.addr;
	// Trace: ../../rtl/VX_pipeline.sv:92:5
	assign icache_req_tag = icache_req_if.tag;
	// Trace: ../../rtl/VX_pipeline.sv:93:5
	assign icache_req_if.ready = icache_req_ready;
	// Trace: ../../rtl/VX_pipeline.sv:99:5
	// expanded interface instance: icache_rsp_if
	localparam _param_396BA_WORD_SIZE = 4;
	localparam _param_396BA_TAG_WIDTH = 45;
	generate
		if (1) begin : icache_rsp_if
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:7:15
			localparam WORD_SIZE = _param_396BA_WORD_SIZE;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:8:15
			localparam TAG_WIDTH = _param_396BA_TAG_WIDTH;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:11:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:12:5
			wire [31:0] data;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:13:5
			wire [44:0] tag;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:14:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:16:5
			// Trace: ../../rtl/interfaces/VX_icache_rsp_if.sv:23:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:104:5
	assign icache_rsp_if.valid = icache_rsp_valid;
	// Trace: ../../rtl/VX_pipeline.sv:105:5
	assign icache_rsp_if.data = icache_rsp_data;
	// Trace: ../../rtl/VX_pipeline.sv:106:5
	assign icache_rsp_if.tag = icache_rsp_tag;
	// Trace: ../../rtl/VX_pipeline.sv:107:5
	assign icache_rsp_ready = icache_rsp_if.ready;
	// Trace: ../../rtl/VX_pipeline.sv:111:5
	// expanded interface instance: fetch_to_csr_if
	generate
		if (1) begin : fetch_to_csr_if
			// Trace: ../../rtl/interfaces/VX_fetch_to_csr_if.sv:8:5
			wire [3:0] thread_masks;
			// Trace: ../../rtl/interfaces/VX_fetch_to_csr_if.sv:10:5
			// Trace: ../../rtl/interfaces/VX_fetch_to_csr_if.sv:14:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:112:5
	// expanded interface instance: cmt_to_csr_if
	generate
		if (1) begin : cmt_to_csr_if
			// Trace: ../../rtl/interfaces/VX_cmt_to_csr_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_cmt_to_csr_if.sv:12:5
			wire [3:0] commit_size;
			// Trace: ../../rtl/interfaces/VX_cmt_to_csr_if.sv:14:5
			// Trace: ../../rtl/interfaces/VX_cmt_to_csr_if.sv:19:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:113:5
	// expanded interface instance: decode_if
	generate
		if (1) begin : decode_if
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:13:5
			wire [2:0] ex_type;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:14:5
			wire [3:0] op_type;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:15:5
			wire [2:0] op_mod;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:16:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:17:5
			wire use_PC;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:18:5
			wire use_imm;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:19:5
			wire [31:0] imm;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:20:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:21:5
			wire [4:0] rs1;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:22:5
			wire [4:0] rs2;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:23:5
			wire [4:0] rs3;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:24:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:26:5
			// Trace: ../../rtl/interfaces/VX_decode_if.sv:46:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:114:5
	// expanded interface instance: branch_ctl_if
	generate
		if (1) begin : branch_ctl_if
			// Trace: ../../rtl/interfaces/VX_branch_ctl_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_branch_ctl_if.sv:9:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_branch_ctl_if.sv:10:5
			wire taken;
			// Trace: ../../rtl/interfaces/VX_branch_ctl_if.sv:11:5
			wire [31:0] dest;
			// Trace: ../../rtl/interfaces/VX_branch_ctl_if.sv:13:5
			// Trace: ../../rtl/interfaces/VX_branch_ctl_if.sv:20:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:115:5
	// expanded interface instance: warp_ctl_if
	generate
		if (1) begin : warp_ctl_if
			// Trace: ../../rtl/interfaces/VX_warp_ctl_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_warp_ctl_if.sv:9:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_warp_ctl_if.sv:10:5
			// removed localparam type gpu_types_gpu_tmc_t
			wire [2:0] tmc;
			// Trace: ../../rtl/interfaces/VX_warp_ctl_if.sv:11:5
			// removed localparam type gpu_types_gpu_wspawn_t
			wire [34:0] wspawn;
			// Trace: ../../rtl/interfaces/VX_warp_ctl_if.sv:12:5
			// removed localparam type gpu_types_gpu_barrier_t
			wire [3:0] barrier;
			// Trace: ../../rtl/interfaces/VX_warp_ctl_if.sv:13:5
			// removed localparam type gpu_types_gpu_split_t
			wire [37:0] split;
			// Trace: ../../rtl/interfaces/VX_warp_ctl_if.sv:15:5
			// Trace: ../../rtl/interfaces/VX_warp_ctl_if.sv:24:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:116:5
	// expanded interface instance: ifetch_rsp_if
	generate
		if (1) begin : ifetch_rsp_if
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:10:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:11:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:13:5
			wire [31:0] data;
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:14:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:16:5
			// Trace: ../../rtl/interfaces/VX_ifetch_rsp_if.sv:26:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:117:5
	// expanded interface instance: alu_req_if
	generate
		if (1) begin : alu_req_if
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:13:5
			wire [31:0] next_PC;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:14:5
			wire [3:0] op_type;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:15:5
			wire [2:0] op_mod;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:16:5
			wire use_PC;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:17:5
			wire use_imm;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:18:5
			wire [31:0] imm;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:19:5
			wire [0:0] tid;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:20:5
			wire [63:0] rs1_data;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:21:5
			wire [63:0] rs2_data;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:22:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:23:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:24:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:26:5
			// Trace: ../../rtl/interfaces/VX_alu_req_if.sv:46:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:118:5
	// expanded interface instance: lsu_req_if
	generate
		if (1) begin : lsu_req_if
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:13:5
			wire [3:0] op_type;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:14:5
			wire is_fence;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:15:5
			wire [63:0] store_data;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:16:5
			wire [63:0] base_addr;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:17:5
			wire [31:0] offset;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:18:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:19:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:20:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:21:5
			wire is_prefetch;
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:23:5
			// Trace: ../../rtl/interfaces/VX_lsu_req_if.sv:40:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:119:5
	// expanded interface instance: csr_req_if
	generate
		if (1) begin : csr_req_if
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:13:5
			wire [1:0] op_type;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:14:5
			wire [11:0] addr;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:15:5
			wire [31:0] rs1_data;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:16:5
			wire use_imm;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:17:5
			wire [4:0] imm;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:18:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:19:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:20:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:22:5
			// Trace: ../../rtl/interfaces/VX_csr_req_if.sv:38:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:123:5
	// expanded interface instance: gpu_req_if
	generate
		if (1) begin : gpu_req_if
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:13:5
			wire [31:0] next_PC;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:14:5
			wire [3:0] op_type;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:15:5
			wire [2:0] op_mod;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:16:5
			wire [0:0] tid;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:17:5
			wire [63:0] rs1_data;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:18:5
			wire [63:0] rs2_data;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:19:5
			wire [63:0] rs3_data;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:20:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:21:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:22:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:24:5
			// Trace: ../../rtl/interfaces/VX_gpu_req_if.sv:42:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:124:5
	// expanded interface instance: writeback_if
	generate
		if (1) begin : writeback_if
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:10:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:11:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:13:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:14:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:15:5
			wire eop;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:16:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:18:5
			// Trace: ../../rtl/interfaces/VX_writeback_if.sv:30:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:125:5
	// expanded interface instance: wstall_if
	generate
		if (1) begin : wstall_if
			// Trace: ../../rtl/interfaces/VX_wstall_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_wstall_if.sv:9:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_wstall_if.sv:10:5
			wire stalled;
			// Trace: ../../rtl/interfaces/VX_wstall_if.sv:12:5
			// Trace: ../../rtl/interfaces/VX_wstall_if.sv:18:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:126:5
	// expanded interface instance: join_if
	generate
		if (1) begin : join_if
			// Trace: ../../rtl/interfaces/VX_join_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_join_if.sv:9:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_join_if.sv:11:5
			// Trace: ../../rtl/interfaces/VX_join_if.sv:16:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:127:5
	// expanded interface instance: alu_commit_if
	generate
		if (1) begin : alu_commit_if
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:13:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:14:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:15:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:16:5
			wire eop;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:17:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:19:5
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:32:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:128:5
	// expanded interface instance: ld_commit_if
	generate
		if (1) begin : ld_commit_if
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:13:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:14:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:15:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:16:5
			wire eop;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:17:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:19:5
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:32:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:129:5
	// expanded interface instance: st_commit_if
	generate
		if (1) begin : st_commit_if
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:13:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:14:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:15:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:16:5
			wire eop;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:17:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:19:5
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:32:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:130:5
	// expanded interface instance: csr_commit_if
	generate
		if (1) begin : csr_commit_if
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:13:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:14:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:15:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:16:5
			wire eop;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:17:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:19:5
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:32:5
		end
	endgenerate
	// Trace: ../../rtl/VX_pipeline.sv:134:5
	// expanded interface instance: gpu_commit_if
	generate
		if (1) begin : gpu_commit_if
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:8:5
			wire valid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:9:5
			wire [43:0] uuid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:10:5
			wire [0:0] wid;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:11:5
			wire [1:0] tmask;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:12:5
			wire [31:0] PC;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:13:5
			wire [63:0] data;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:14:5
			wire [4:0] rd;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:15:5
			wire wb;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:16:5
			wire eop;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:17:5
			wire ready;
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:19:5
			// Trace: ../../rtl/interfaces/VX_commit_if.sv:32:5
		end
	endgenerate
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:140:24
	wire fetch_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:140:57
	VX_reset_relay __fetch_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(fetch_reset)
	);
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:141:25
	wire decode_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:141:58
	VX_reset_relay __decode_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(decode_reset)
	);
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:142:24
	wire issue_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:142:57
	VX_reset_relay __issue_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(issue_reset)
	);
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:143:26
	wire execute_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:143:59
	VX_reset_relay __execute_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(execute_reset)
	);
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:144:25
	wire commit_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_pipeline.sv:144:58
	VX_reset_relay __commit_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(commit_reset)
	);
	// Trace: ../../rtl/VX_pipeline.sv:146:5
	// expanded module instance: fetch
	localparam _param_852F6_CORE_ID = CORE_ID;
	function automatic signed [43:0] sv2v_cast_44_signed;
		input reg signed [43:0] inp;
		sv2v_cast_44_signed = inp;
	endfunction
	generate
		if (1) begin : fetch
			// Trace: ../../rtl/VX_fetch.sv:4:15
			localparam CORE_ID = _param_852F6_CORE_ID;
			// Trace: ../../rtl/VX_fetch.sv:8:5
			wire clk;
			// Trace: ../../rtl/VX_fetch.sv:9:5
			wire reset;
			// Trace: ../../rtl/VX_fetch.sv:12:5
			// removed modport instance icache_req_if
			// Trace: ../../rtl/VX_fetch.sv:13:5
			// removed modport instance icache_rsp_if
			// Trace: ../../rtl/VX_fetch.sv:16:5
			// removed modport instance wstall_if
			// Trace: ../../rtl/VX_fetch.sv:17:5
			// removed modport instance join_if
			// Trace: ../../rtl/VX_fetch.sv:18:5
			// removed modport instance branch_ctl_if
			// Trace: ../../rtl/VX_fetch.sv:19:5
			// removed modport instance warp_ctl_if
			// Trace: ../../rtl/VX_fetch.sv:22:5
			// removed modport instance ifetch_rsp_if
			// Trace: ../../rtl/VX_fetch.sv:25:5
			// removed modport instance fetch_to_csr_if
			// Trace: ../../rtl/VX_fetch.sv:28:5
			wire busy;
			// Trace: ../../rtl/VX_fetch.sv:31:5
			// expanded interface instance: ifetch_req_if
			if (1) begin : ifetch_req_if
				// Trace: ../../rtl/interfaces/VX_ifetch_req_if.sv:8:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_ifetch_req_if.sv:9:5
				wire [43:0] uuid;
				// Trace: ../../rtl/interfaces/VX_ifetch_req_if.sv:10:5
				wire [1:0] tmask;
				// Trace: ../../rtl/interfaces/VX_ifetch_req_if.sv:11:5
				wire [0:0] wid;
				// Trace: ../../rtl/interfaces/VX_ifetch_req_if.sv:12:5
				wire [31:0] PC;
				// Trace: ../../rtl/interfaces/VX_ifetch_req_if.sv:13:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_ifetch_req_if.sv:15:5
				// Trace: ../../rtl/interfaces/VX_ifetch_req_if.sv:24:5
			end
			// Trace: ../../rtl/VX_fetch.sv:33:5
			// expanded module instance: warp_sched
			localparam _param_4F3BC_CORE_ID = CORE_ID;
			if (1) begin : warp_sched
				// Trace: ../../rtl/VX_warp_sched.sv:4:15
				localparam CORE_ID = _param_4F3BC_CORE_ID;
				// Trace: ../../rtl/VX_warp_sched.sv:8:5
				wire clk;
				// Trace: ../../rtl/VX_warp_sched.sv:9:5
				wire reset;
				// Trace: ../../rtl/VX_warp_sched.sv:11:5
				// removed modport instance warp_ctl_if
				// Trace: ../../rtl/VX_warp_sched.sv:12:5
				// removed modport instance wstall_if
				// Trace: ../../rtl/VX_warp_sched.sv:13:5
				// removed modport instance join_if
				// Trace: ../../rtl/VX_warp_sched.sv:14:5
				// removed modport instance branch_ctl_if
				// Trace: ../../rtl/VX_warp_sched.sv:16:5
				// removed modport instance ifetch_req_if
				// Trace: ../../rtl/VX_warp_sched.sv:18:5
				// removed modport instance fetch_to_csr_if
				// Trace: ../../rtl/VX_warp_sched.sv:20:5
				wire busy;
				// Trace: ../../rtl/VX_warp_sched.sv:25:5
				wire join_else;
				// Trace: ../../rtl/VX_warp_sched.sv:26:5
				wire [31:0] join_pc;
				// Trace: ../../rtl/VX_warp_sched.sv:27:5
				wire [1:0] join_tmask;
				// Trace: ../../rtl/VX_warp_sched.sv:29:5
				reg [1:0] active_warps;
				reg [1:0] active_warps_n;
				// Trace: ../../rtl/VX_warp_sched.sv:30:5
				reg [1:0] stalled_warps;
				// Trace: ../../rtl/VX_warp_sched.sv:32:5
				reg [3:0] thread_masks;
				// Trace: ../../rtl/VX_warp_sched.sv:33:5
				reg [63:0] warp_pcs;
				// Trace: ../../rtl/VX_warp_sched.sv:36:5
				reg [7:0] barrier_masks;
				// Trace: ../../rtl/VX_warp_sched.sv:37:5
				wire reached_barrier_limit;
				// Trace: ../../rtl/VX_warp_sched.sv:40:5
				reg [31:0] wspawn_pc;
				// Trace: ../../rtl/VX_warp_sched.sv:41:5
				reg [1:0] use_wspawn;
				// Trace: ../../rtl/VX_warp_sched.sv:43:5
				wire [0:0] schedule_wid;
				// Trace: ../../rtl/VX_warp_sched.sv:44:5
				wire [1:0] schedule_tmask;
				// Trace: ../../rtl/VX_warp_sched.sv:45:5
				wire [31:0] schedule_pc;
				// Trace: ../../rtl/VX_warp_sched.sv:46:5
				wire schedule_valid;
				// Trace: ../../rtl/VX_warp_sched.sv:47:5
				wire warp_scheduled;
				// Trace: ../../rtl/VX_warp_sched.sv:49:5
				reg [43:0] issued_instrs;
				// Trace: ../../rtl/VX_warp_sched.sv:51:5
				wire ifetch_req_fire = VX_pipeline.fetch.ifetch_req_if.valid && VX_pipeline.fetch.ifetch_req_if.ready;
				// Trace: ../../rtl/VX_warp_sched.sv:53:5
				wire tmc_active = VX_pipeline.warp_ctl_if.tmc[1-:2] != 0;
				// Trace: ../../rtl/VX_warp_sched.sv:55:5
				always @(*) begin
					// Trace: ../../rtl/VX_warp_sched.sv:56:9
					active_warps_n = active_warps;
					// Trace: ../../rtl/VX_warp_sched.sv:57:9
					if (VX_pipeline.warp_ctl_if.valid && VX_pipeline.warp_ctl_if.wspawn[34])
						// Trace: ../../rtl/VX_warp_sched.sv:58:13
						active_warps_n = VX_pipeline.warp_ctl_if.wspawn[33-:2];
					if (VX_pipeline.warp_ctl_if.valid && VX_pipeline.warp_ctl_if.tmc[2])
						// Trace: ../../rtl/VX_warp_sched.sv:61:13
						active_warps_n[VX_pipeline.warp_ctl_if.wid] = tmc_active;
				end
				// Trace: ../../rtl/VX_warp_sched.sv:65:5
				always @(posedge clk)
					// Trace: ../../rtl/VX_warp_sched.sv:66:9
					if (reset) begin
						// Trace: ../../rtl/VX_warp_sched.sv:67:13
						barrier_masks <= 1'sb0;
						// Trace: ../../rtl/VX_warp_sched.sv:68:13
						use_wspawn <= 1'sb0;
						// Trace: ../../rtl/VX_warp_sched.sv:69:13
						stalled_warps <= 1'sb0;
						// Trace: ../../rtl/VX_warp_sched.sv:70:13
						warp_pcs <= 1'sb0;
						// Trace: ../../rtl/VX_warp_sched.sv:71:13
						active_warps <= 1'sb0;
						// Trace: ../../rtl/VX_warp_sched.sv:72:13
						thread_masks <= 1'sb0;
						// Trace: ../../rtl/VX_warp_sched.sv:73:13
						issued_instrs <= 1'sb0;
						// Trace: ../../rtl/VX_warp_sched.sv:76:13
						warp_pcs[0+:32] <= 32'h80000000;
						// Trace: ../../rtl/VX_warp_sched.sv:77:13
						active_warps[0] <= 1;
						// Trace: ../../rtl/VX_warp_sched.sv:78:13
						thread_masks[0+:2] <= 1;
					end
					else begin
						// Trace: ../../rtl/VX_warp_sched.sv:80:13
						if (VX_pipeline.warp_ctl_if.valid && VX_pipeline.warp_ctl_if.wspawn[34]) begin
							// Trace: ../../rtl/VX_warp_sched.sv:81:17
							use_wspawn <= VX_pipeline.warp_ctl_if.wspawn[33-:2] & ~2'sd1;
							// Trace: ../../rtl/VX_warp_sched.sv:82:17
							wspawn_pc <= VX_pipeline.warp_ctl_if.wspawn[31-:32];
						end
						if (VX_pipeline.warp_ctl_if.valid && VX_pipeline.warp_ctl_if.barrier[3]) begin
							// Trace: ../../rtl/VX_warp_sched.sv:86:17
							stalled_warps[VX_pipeline.warp_ctl_if.wid] <= 0;
							// Trace: ../../rtl/VX_warp_sched.sv:87:17
							if (reached_barrier_limit)
								// Trace: ../../rtl/VX_warp_sched.sv:88:21
								barrier_masks[VX_pipeline.warp_ctl_if.barrier[2-:2] * 2+:2] <= 0;
							else
								// Trace: ../../rtl/VX_warp_sched.sv:90:21
								barrier_masks[(VX_pipeline.warp_ctl_if.barrier[2-:2] * 2) + VX_pipeline.warp_ctl_if.wid] <= 1;
						end
						if (VX_pipeline.warp_ctl_if.valid && VX_pipeline.warp_ctl_if.tmc[2]) begin
							// Trace: ../../rtl/VX_warp_sched.sv:95:17
							thread_masks[VX_pipeline.warp_ctl_if.wid * 2+:2] <= VX_pipeline.warp_ctl_if.tmc[1-:2];
							// Trace: ../../rtl/VX_warp_sched.sv:96:17
							stalled_warps[VX_pipeline.warp_ctl_if.wid] <= 0;
						end
						if (VX_pipeline.warp_ctl_if.valid && VX_pipeline.warp_ctl_if.split[37]) begin
							// Trace: ../../rtl/VX_warp_sched.sv:100:17
							stalled_warps[VX_pipeline.warp_ctl_if.wid] <= 0;
							// Trace: ../../rtl/VX_warp_sched.sv:101:17
							if (VX_pipeline.warp_ctl_if.split[36])
								// Trace: ../../rtl/VX_warp_sched.sv:102:21
								thread_masks[VX_pipeline.warp_ctl_if.wid * 2+:2] <= VX_pipeline.warp_ctl_if.split[35-:2];
						end
						if (VX_pipeline.branch_ctl_if.valid) begin
							// Trace: ../../rtl/VX_warp_sched.sv:108:17
							if (VX_pipeline.branch_ctl_if.taken)
								// Trace: ../../rtl/VX_warp_sched.sv:109:21
								warp_pcs[VX_pipeline.branch_ctl_if.wid * 32+:32] <= VX_pipeline.branch_ctl_if.dest;
							// Trace: ../../rtl/VX_warp_sched.sv:111:17
							stalled_warps[VX_pipeline.branch_ctl_if.wid] <= 0;
						end
						if (warp_scheduled) begin
							// Trace: ../../rtl/VX_warp_sched.sv:116:17
							stalled_warps[schedule_wid] <= 1;
							// Trace: ../../rtl/VX_warp_sched.sv:119:17
							use_wspawn[schedule_wid] <= 0;
							// Trace: ../../rtl/VX_warp_sched.sv:120:17
							if (use_wspawn[schedule_wid])
								// Trace: ../../rtl/VX_warp_sched.sv:121:21
								thread_masks[schedule_wid * 2+:2] <= 1;
							// Trace: ../../rtl/VX_warp_sched.sv:124:17
							issued_instrs <= issued_instrs + 1;
						end
						if (ifetch_req_fire)
							// Trace: ../../rtl/VX_warp_sched.sv:128:17
							warp_pcs[VX_pipeline.fetch.ifetch_req_if.wid * 32+:32] <= VX_pipeline.fetch.ifetch_req_if.PC + 4;
						if (VX_pipeline.wstall_if.valid)
							// Trace: ../../rtl/VX_warp_sched.sv:132:17
							stalled_warps[VX_pipeline.wstall_if.wid] <= VX_pipeline.wstall_if.stalled;
						if (VX_pipeline.join_if.valid) begin
							// Trace: ../../rtl/VX_warp_sched.sv:137:17
							if (join_else)
								// Trace: ../../rtl/VX_warp_sched.sv:138:21
								warp_pcs[VX_pipeline.join_if.wid * 32+:32] <= join_pc;
							// Trace: ../../rtl/VX_warp_sched.sv:140:17
							thread_masks[VX_pipeline.join_if.wid * 2+:2] <= join_tmask;
						end
						// Trace: ../../rtl/VX_warp_sched.sv:143:13
						active_warps <= active_warps_n;
					end
				// Trace: ../../rtl/VX_warp_sched.sv:148:5
				assign VX_pipeline.fetch_to_csr_if.thread_masks = thread_masks;
				// Trace: ../../rtl/VX_warp_sched.sv:153:5
				wire [1:0] active_barrier_count;
				// Trace: ../../rtl/VX_warp_sched.sv:155:5
				wire [1:0] barrier_mask = barrier_masks[VX_pipeline.warp_ctl_if.barrier[2-:2] * 2+:2];
				// Trace: macro expansion of POP_COUNT at ../../rtl/VX_warp_sched.sv:156:46
				VX_popcount #(.N(2)) __active_barrier_count(
					.in_i(barrier_mask),
					.cnt_o(active_barrier_count)
				);
				// Trace: ../../rtl/VX_warp_sched.sv:158:5
				assign reached_barrier_limit = active_barrier_count[0:0] == VX_pipeline.warp_ctl_if.barrier[0-:1];
				// Trace: ../../rtl/VX_warp_sched.sv:160:5
				reg [1:0] barrier_stalls;
				// Trace: ../../rtl/VX_warp_sched.sv:161:5
				always @(*) begin
					// Trace: ../../rtl/VX_warp_sched.sv:162:9
					barrier_stalls = barrier_masks[0+:2];
					// Trace: ../../rtl/VX_warp_sched.sv:163:9
					begin : sv2v_autoblock_1
						// Trace: ../../rtl/VX_warp_sched.sv:163:14
						integer i;
						// Trace: ../../rtl/VX_warp_sched.sv:163:14
						for (i = 1; i < 4; i = i + 1)
							begin
								// Trace: ../../rtl/VX_warp_sched.sv:164:13
								barrier_stalls = barrier_stalls | barrier_masks[i * 2+:2];
							end
					end
				end
				// Trace: ../../rtl/VX_warp_sched.sv:170:5
				wire [33:0] ipdom_data [1:0];
				// Trace: ../../rtl/VX_warp_sched.sv:171:5
				wire ipdom_index [1:0];
				// Trace: ../../rtl/VX_warp_sched.sv:173:5
				genvar i;
				for (i = 0; i < 2; i = i + 1) begin : genblk1
					// Trace: ../../rtl/VX_warp_sched.sv:174:9
					wire push = (VX_pipeline.warp_ctl_if.valid && VX_pipeline.warp_ctl_if.split[37]) && (i == VX_pipeline.warp_ctl_if.wid);
					// Trace: ../../rtl/VX_warp_sched.sv:178:9
					wire pop = VX_pipeline.join_if.valid && (i == VX_pipeline.join_if.wid);
					// Trace: ../../rtl/VX_warp_sched.sv:180:9
					wire [1:0] else_tmask = VX_pipeline.warp_ctl_if.split[33-:2];
					// Trace: ../../rtl/VX_warp_sched.sv:181:9
					wire [1:0] orig_tmask = thread_masks[VX_pipeline.warp_ctl_if.wid * 2+:2];
					// Trace: ../../rtl/VX_warp_sched.sv:183:9
					wire [33:0] q_else = {VX_pipeline.warp_ctl_if.split[31-:32], else_tmask};
					// Trace: ../../rtl/VX_warp_sched.sv:184:9
					wire [33:0] q_end = {32'b00000000000000000000000000000000, orig_tmask};
					// Trace: ../../rtl/VX_warp_sched.sv:186:9
					VX_ipdom_stack #(
						.WIDTH(34),
						.DEPTH(4)
					) ipdom_stack(
						.clk(clk),
						.reset(reset),
						.push(push),
						.pop(pop),
						.pair(VX_pipeline.warp_ctl_if.split[36]),
						.q1(q_end),
						.q2(q_else),
						.d(ipdom_data[i]),
						.index(ipdom_index[i])
					);
				end
				// Trace: ../../rtl/VX_warp_sched.sv:204:5
				assign {join_pc, join_tmask} = ipdom_data[VX_pipeline.join_if.wid];
				// Trace: ../../rtl/VX_warp_sched.sv:205:5
				assign join_else = ~ipdom_index[VX_pipeline.join_if.wid];
				// Trace: ../../rtl/VX_warp_sched.sv:209:5
				wire [1:0] ready_warps = active_warps & ~(stalled_warps | barrier_stalls);
				// Trace: ../../rtl/VX_warp_sched.sv:211:5
				VX_lzc #(.N(2)) wid_select(
					.in_i(ready_warps),
					.cnt_o(schedule_wid),
					.valid_o(schedule_valid)
				);
				// Trace: ../../rtl/VX_warp_sched.sv:219:5
				wire [67:0] schedule_data;
				// Trace: ../../rtl/VX_warp_sched.sv:220:5
				for (i = 0; i < 2; i = i + 1) begin : genblk2
					// Trace: ../../rtl/VX_warp_sched.sv:221:9
					assign schedule_data[i * 34+:34] = {(use_wspawn[i] ? 2'sd1 : thread_masks[i * 2+:2]), (use_wspawn[i] ? wspawn_pc : warp_pcs[i * 32+:32])};
				end
				// Trace: ../../rtl/VX_warp_sched.sv:225:5
				assign {schedule_tmask, schedule_pc} = schedule_data[schedule_wid * 34+:34];
				// Trace: ../../rtl/VX_warp_sched.sv:227:5
				wire stall_out = ~VX_pipeline.fetch.ifetch_req_if.ready && VX_pipeline.fetch.ifetch_req_if.valid;
				// Trace: ../../rtl/VX_warp_sched.sv:229:5
				assign warp_scheduled = schedule_valid && ~stall_out;
				// Trace: ../../rtl/VX_warp_sched.sv:231:5
				wire [43:0] instr_uuid = ((issued_instrs * 1) * 1) + sv2v_cast_44_signed(CORE_ID);
				// Trace: ../../rtl/VX_warp_sched.sv:233:5
				VX_pipe_register #(
					.DATAW(80),
					.RESETW(1)
				) pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(!stall_out),
					.data_in({schedule_valid, instr_uuid, schedule_tmask, schedule_pc, schedule_wid}),
					.data_out({VX_pipeline.fetch.ifetch_req_if.valid, VX_pipeline.fetch.ifetch_req_if.uuid, VX_pipeline.fetch.ifetch_req_if.tmask, VX_pipeline.fetch.ifetch_req_if.PC, VX_pipeline.fetch.ifetch_req_if.wid})
				);
				// Trace: ../../rtl/VX_warp_sched.sv:244:5
				assign busy = active_warps != 0;
			end
			assign warp_sched.clk = clk;
			assign warp_sched.reset = reset;
			assign busy = warp_sched.busy;
			// Trace: ../../rtl/VX_fetch.sv:53:5
			// expanded module instance: icache_stage
			localparam _param_8CCB0_CORE_ID = CORE_ID;
			if (1) begin : icache_stage
				// Trace: ../../rtl/VX_icache_stage.sv:4:15
				localparam CORE_ID = _param_8CCB0_CORE_ID;
				// Trace: ../../rtl/VX_icache_stage.sv:8:5
				wire clk;
				// Trace: ../../rtl/VX_icache_stage.sv:9:5
				wire reset;
				// Trace: ../../rtl/VX_icache_stage.sv:12:5
				// removed modport instance icache_req_if
				// Trace: ../../rtl/VX_icache_stage.sv:13:5
				// removed modport instance icache_rsp_if
				// Trace: ../../rtl/VX_icache_stage.sv:16:5
				// removed modport instance ifetch_req_if
				// Trace: ../../rtl/VX_icache_stage.sv:19:5
				// removed modport instance ifetch_rsp_if
				// Trace: ../../rtl/VX_icache_stage.sv:25:5
				localparam OUT_REG = 0;
				// Trace: ../../rtl/VX_icache_stage.sv:27:5
				wire [0:0] req_tag;
				wire [0:0] rsp_tag;
				// Trace: ../../rtl/VX_icache_stage.sv:29:5
				wire icache_req_fire = VX_pipeline.icache_req_if.valid && VX_pipeline.icache_req_if.ready;
				// Trace: ../../rtl/VX_icache_stage.sv:31:5
				assign req_tag = VX_pipeline.fetch.ifetch_req_if.wid;
				// Trace: ../../rtl/VX_icache_stage.sv:32:5
				assign rsp_tag = VX_pipeline.icache_rsp_if.tag[0:0];
				// Trace: ../../rtl/VX_icache_stage.sv:34:5
				wire [43:0] rsp_uuid;
				// Trace: ../../rtl/VX_icache_stage.sv:35:5
				wire [31:0] rsp_PC;
				// Trace: ../../rtl/VX_icache_stage.sv:36:5
				wire [1:0] rsp_tmask;
				// Trace: ../../rtl/VX_icache_stage.sv:38:5
				VX_dp_ram #(
					.DATAW(78),
					.SIZE(2),
					.LUTRAM(1)
				) req_metadata(
					.clk(clk),
					.wren(icache_req_fire),
					.waddr(req_tag),
					.wdata({VX_pipeline.fetch.ifetch_req_if.PC, VX_pipeline.fetch.ifetch_req_if.tmask, VX_pipeline.fetch.ifetch_req_if.uuid}),
					.raddr(rsp_tag),
					.rdata({rsp_PC, rsp_tmask, rsp_uuid})
				);
				// Trace: ../../rtl/VX_icache_stage.sv:55:5
				assign VX_pipeline.icache_req_if.valid = VX_pipeline.fetch.ifetch_req_if.valid;
				// Trace: ../../rtl/VX_icache_stage.sv:56:5
				assign VX_pipeline.icache_req_if.addr = VX_pipeline.fetch.ifetch_req_if.PC[31:2];
				// Trace: ../../rtl/VX_icache_stage.sv:57:5
				assign VX_pipeline.icache_req_if.tag = {VX_pipeline.fetch.ifetch_req_if.uuid, req_tag};
				// Trace: ../../rtl/VX_icache_stage.sv:60:5
				assign VX_pipeline.fetch.ifetch_req_if.ready = VX_pipeline.icache_req_if.ready;
				// Trace: ../../rtl/VX_icache_stage.sv:62:5
				wire [0:0] rsp_wid = rsp_tag;
				// Trace: ../../rtl/VX_icache_stage.sv:64:5
				wire stall_out = ~VX_pipeline.ifetch_rsp_if.ready && (1'd1 && VX_pipeline.ifetch_rsp_if.valid);
				// Trace: ../../rtl/VX_icache_stage.sv:66:5
				VX_pipe_register #(
					.DATAW(112),
					.RESETW(1),
					.DEPTH(OUT_REG)
				) pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(!stall_out),
					.data_in({VX_pipeline.icache_rsp_if.valid, rsp_wid, rsp_tmask, rsp_PC, VX_pipeline.icache_rsp_if.data, rsp_uuid}),
					.data_out({VX_pipeline.ifetch_rsp_if.valid, VX_pipeline.ifetch_rsp_if.wid, VX_pipeline.ifetch_rsp_if.tmask, VX_pipeline.ifetch_rsp_if.PC, VX_pipeline.ifetch_rsp_if.data, VX_pipeline.ifetch_rsp_if.uuid})
				);
				// Trace: ../../rtl/VX_icache_stage.sv:79:5
				assign VX_pipeline.icache_rsp_if.ready = ~stall_out;
			end
			assign icache_stage.clk = clk;
			assign icache_stage.reset = reset;
		end
	endgenerate
	assign fetch.clk = clk;
	assign fetch.reset = fetch_reset;
	assign busy = fetch.busy;
	// Trace: ../../rtl/VX_pipeline.sv:163:5
	// expanded module instance: decode
	localparam _param_21B54_CORE_ID = CORE_ID;
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	generate
		if (1) begin : decode
			// Trace: ../../rtl/VX_decode.sv:18:15
			localparam CORE_ID = _param_21B54_CORE_ID;
			// Trace: ../../rtl/VX_decode.sv:20:5
			wire clk;
			// Trace: ../../rtl/VX_decode.sv:21:5
			wire reset;
			// Trace: ../../rtl/VX_decode.sv:28:5
			// removed modport instance ifetch_rsp_if
			// Trace: ../../rtl/VX_decode.sv:31:5
			// removed modport instance decode_if
			// Trace: ../../rtl/VX_decode.sv:32:5
			// removed modport instance wstall_if
			// Trace: ../../rtl/VX_decode.sv:33:5
			// removed modport instance join_if
			// Trace: ../../rtl/VX_decode.sv:39:5
			reg [2:0] ex_type;
			// Trace: ../../rtl/VX_decode.sv:40:5
			reg [3:0] op_type;
			// Trace: ../../rtl/VX_decode.sv:41:5
			reg [2:0] op_mod;
			// Trace: ../../rtl/VX_decode.sv:42:5
			reg [4:0] rd_r;
			reg [4:0] rs1_r;
			reg [4:0] rs2_r;
			reg [4:0] rs3_r;
			// Trace: ../../rtl/VX_decode.sv:43:5
			reg [31:0] imm;
			// Trace: ../../rtl/VX_decode.sv:44:5
			reg use_rd;
			reg use_PC;
			reg use_imm;
			// Trace: ../../rtl/VX_decode.sv:45:5
			reg is_join;
			reg is_wstall;
			// Trace: ../../rtl/VX_decode.sv:47:5
			wire [31:0] instr = VX_pipeline.ifetch_rsp_if.data;
			// Trace: ../../rtl/VX_decode.sv:48:5
			wire [6:0] opcode = instr[6:0];
			// Trace: ../../rtl/VX_decode.sv:49:5
			wire [1:0] func2 = instr[26:25];
			// Trace: ../../rtl/VX_decode.sv:50:5
			wire [2:0] func3 = instr[14:12];
			// Trace: ../../rtl/VX_decode.sv:51:5
			wire [6:0] func7 = instr[31:25];
			// Trace: ../../rtl/VX_decode.sv:52:5
			wire [11:0] u_12 = instr[31:20];
			// Trace: ../../rtl/VX_decode.sv:54:5
			wire [4:0] rd = instr[11:7];
			// Trace: ../../rtl/VX_decode.sv:55:5
			wire [4:0] rs1 = instr[19:15];
			// Trace: ../../rtl/VX_decode.sv:56:5
			wire [4:0] rs2 = instr[24:20];
			// Trace: ../../rtl/VX_decode.sv:57:5
			wire [4:0] rs3 = instr[31:27];
			// Trace: ../../rtl/VX_decode.sv:59:5
			wire [19:0] upper_imm = {func7, rs2, rs1, func3};
			// Trace: ../../rtl/VX_decode.sv:60:5
			wire [11:0] alu_imm = (func3[0] && ~func3[1] ? {{7 {1'b0}}, rs2} : u_12);
			// Trace: ../../rtl/VX_decode.sv:61:5
			wire [11:0] s_imm = {func7, rd};
			// Trace: ../../rtl/VX_decode.sv:62:5
			wire [12:0] b_imm = {instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
			// Trace: ../../rtl/VX_decode.sv:63:5
			wire [20:0] jal_imm = {instr[31], instr[19:12], instr[20], instr[30:21], 1'b0};
			// Trace: ../../rtl/VX_decode.sv:67:5
			always @(*) begin
				// Trace: ../../rtl/VX_decode.sv:69:9
				ex_type = 0;
				// Trace: ../../rtl/VX_decode.sv:70:9
				op_type = 1'sbx;
				// Trace: ../../rtl/VX_decode.sv:71:9
				op_mod = 0;
				// Trace: ../../rtl/VX_decode.sv:72:9
				rd_r = 0;
				// Trace: ../../rtl/VX_decode.sv:73:9
				rs1_r = 0;
				// Trace: ../../rtl/VX_decode.sv:74:9
				rs2_r = 0;
				// Trace: ../../rtl/VX_decode.sv:75:9
				rs3_r = 0;
				// Trace: ../../rtl/VX_decode.sv:76:9
				imm = 1'sbx;
				// Trace: ../../rtl/VX_decode.sv:77:9
				use_imm = 0;
				// Trace: ../../rtl/VX_decode.sv:78:9
				use_PC = 0;
				// Trace: ../../rtl/VX_decode.sv:79:9
				use_rd = 0;
				// Trace: ../../rtl/VX_decode.sv:80:9
				is_join = 0;
				// Trace: ../../rtl/VX_decode.sv:81:9
				is_wstall = 0;
				// Trace: ../../rtl/VX_decode.sv:83:9
				case (opcode)
					7'b0010011: begin
						// Trace: ../../rtl/VX_decode.sv:85:17
						ex_type = 3'h1;
						// Trace: ../../rtl/VX_decode.sv:86:17
						case (func3)
							3'h0:
								// Trace: ../../rtl/VX_decode.sv:87:27
								op_type = 4'b0000;
							3'h1:
								// Trace: ../../rtl/VX_decode.sv:88:27
								op_type = 4'b1111;
							3'h2:
								// Trace: ../../rtl/VX_decode.sv:89:27
								op_type = 4'b0101;
							3'h3:
								// Trace: ../../rtl/VX_decode.sv:90:27
								op_type = 4'b0100;
							3'h4:
								// Trace: ../../rtl/VX_decode.sv:91:27
								op_type = 4'b1110;
							3'h5:
								// Trace: ../../rtl/VX_decode.sv:92:27
								op_type = (func7[5] ? 4'b1001 : 4'b1000);
							3'h6:
								// Trace: ../../rtl/VX_decode.sv:93:27
								op_type = 4'b1101;
							3'h7:
								// Trace: ../../rtl/VX_decode.sv:94:27
								op_type = 4'b1100;
							default:
								;
						endcase
						// Trace: ../../rtl/VX_decode.sv:97:17
						use_rd = 1;
						// Trace: ../../rtl/VX_decode.sv:98:17
						use_imm = 1;
						// Trace: ../../rtl/VX_decode.sv:99:17
						imm = {{20 {alu_imm[11]}}, alu_imm};
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:100:31
						rd_r = rd;
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:101:32
						rs1_r = rs1;
					end
					7'b0110011: begin
						// Trace: ../../rtl/VX_decode.sv:104:17
						ex_type = 3'h1;
						// Trace: ../../rtl/VX_decode.sv:121:17
						// Trace: ../../rtl/VX_decode.sv:122:21
						case (func3)
							3'h0:
								// Trace: ../../rtl/VX_decode.sv:123:31
								op_type = (func7[5] ? 4'b1011 : 4'b0000);
							3'h1:
								// Trace: ../../rtl/VX_decode.sv:124:31
								op_type = 4'b1111;
							3'h2:
								// Trace: ../../rtl/VX_decode.sv:125:31
								op_type = 4'b0101;
							3'h3:
								// Trace: ../../rtl/VX_decode.sv:126:31
								op_type = 4'b0100;
							3'h4:
								// Trace: ../../rtl/VX_decode.sv:127:31
								op_type = 4'b1110;
							3'h5:
								// Trace: ../../rtl/VX_decode.sv:128:31
								op_type = (func7[5] ? 4'b1001 : 4'b1000);
							3'h6:
								// Trace: ../../rtl/VX_decode.sv:129:31
								op_type = 4'b1101;
							3'h7:
								// Trace: ../../rtl/VX_decode.sv:130:31
								op_type = 4'b1100;
							default:
								;
						endcase
						// Trace: ../../rtl/VX_decode.sv:134:17
						use_rd = 1;
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:135:31
						rd_r = rd;
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:136:32
						rs1_r = rs1;
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:137:32
						rs2_r = rs2;
					end
					7'b0110111: begin
						// Trace: ../../rtl/VX_decode.sv:140:17
						ex_type = 3'h1;
						// Trace: ../../rtl/VX_decode.sv:141:17
						op_type = 4'b0010;
						// Trace: ../../rtl/VX_decode.sv:142:17
						use_rd = 1;
						// Trace: ../../rtl/VX_decode.sv:143:17
						use_imm = 1;
						// Trace: ../../rtl/VX_decode.sv:144:17
						imm = {upper_imm, 12'sd0};
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:145:31
						rd_r = rd;
						// Trace: ../../rtl/VX_decode.sv:146:17
						rs1_r = 0;
					end
					7'b0010111: begin
						// Trace: ../../rtl/VX_decode.sv:149:17
						ex_type = 3'h1;
						// Trace: ../../rtl/VX_decode.sv:150:17
						op_type = 4'b0011;
						// Trace: ../../rtl/VX_decode.sv:151:17
						use_rd = 1;
						// Trace: ../../rtl/VX_decode.sv:152:17
						use_imm = 1;
						// Trace: ../../rtl/VX_decode.sv:153:17
						use_PC = 1;
						// Trace: ../../rtl/VX_decode.sv:154:17
						imm = {upper_imm, 12'sd0};
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:155:31
						rd_r = rd;
					end
					7'b1101111: begin
						// Trace: ../../rtl/VX_decode.sv:158:17
						ex_type = 3'h1;
						// Trace: ../../rtl/VX_decode.sv:159:17
						op_type = 4'b1000;
						// Trace: ../../rtl/VX_decode.sv:160:17
						op_mod = 1;
						// Trace: ../../rtl/VX_decode.sv:161:17
						use_rd = 1;
						// Trace: ../../rtl/VX_decode.sv:162:17
						use_imm = 1;
						// Trace: ../../rtl/VX_decode.sv:163:17
						use_PC = 1;
						// Trace: ../../rtl/VX_decode.sv:164:17
						is_wstall = 1;
						// Trace: ../../rtl/VX_decode.sv:165:17
						imm = {{11 {jal_imm[20]}}, jal_imm};
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:166:31
						rd_r = rd;
					end
					7'b1100111: begin
						// Trace: ../../rtl/VX_decode.sv:169:17
						ex_type = 3'h1;
						// Trace: ../../rtl/VX_decode.sv:170:17
						op_type = 4'b1001;
						// Trace: ../../rtl/VX_decode.sv:171:17
						op_mod = 1;
						// Trace: ../../rtl/VX_decode.sv:172:17
						use_rd = 1;
						// Trace: ../../rtl/VX_decode.sv:173:17
						use_imm = 1;
						// Trace: ../../rtl/VX_decode.sv:174:17
						is_wstall = 1;
						// Trace: ../../rtl/VX_decode.sv:175:17
						imm = {{20 {u_12[11]}}, u_12};
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:176:31
						rd_r = rd;
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:177:32
						rs1_r = rs1;
					end
					7'b1100011: begin
						// Trace: ../../rtl/VX_decode.sv:180:17
						ex_type = 3'h1;
						// Trace: ../../rtl/VX_decode.sv:181:17
						case (func3)
							3'h0:
								// Trace: ../../rtl/VX_decode.sv:182:27
								op_type = 4'b0000;
							3'h1:
								// Trace: ../../rtl/VX_decode.sv:183:27
								op_type = 4'b0010;
							3'h4:
								// Trace: ../../rtl/VX_decode.sv:184:27
								op_type = 4'b0101;
							3'h5:
								// Trace: ../../rtl/VX_decode.sv:185:27
								op_type = 4'b0111;
							3'h6:
								// Trace: ../../rtl/VX_decode.sv:186:27
								op_type = 4'b0100;
							3'h7:
								// Trace: ../../rtl/VX_decode.sv:187:27
								op_type = 4'b0110;
							default:
								;
						endcase
						// Trace: ../../rtl/VX_decode.sv:190:17
						op_mod = 1;
						// Trace: ../../rtl/VX_decode.sv:191:17
						use_imm = 1;
						// Trace: ../../rtl/VX_decode.sv:192:17
						use_PC = 1;
						// Trace: ../../rtl/VX_decode.sv:193:17
						is_wstall = 1;
						// Trace: ../../rtl/VX_decode.sv:194:17
						imm = {{19 {b_imm[12]}}, b_imm};
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:195:32
						rs1_r = rs1;
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:196:32
						rs2_r = rs2;
					end
					7'b0001111: begin
						// Trace: ../../rtl/VX_decode.sv:199:17
						ex_type = 3'h2;
						// Trace: ../../rtl/VX_decode.sv:200:17
						op_mod = 3'sd1;
					end
					7'b1110011:
						// Trace: ../../rtl/VX_decode.sv:203:17
						if (func3[1:0] != 0) begin
							// Trace: ../../rtl/VX_decode.sv:204:21
							ex_type = 3'h3;
							// Trace: ../../rtl/VX_decode.sv:205:21
							op_type = sv2v_cast_4(func3[1:0]);
							// Trace: ../../rtl/VX_decode.sv:206:21
							use_rd = 1;
							// Trace: ../../rtl/VX_decode.sv:207:21
							use_imm = func3[2];
							// Trace: ../../rtl/VX_decode.sv:208:21
							imm[11:0] = u_12;
							// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:209:35
							rd_r = rd;
							// Trace: ../../rtl/VX_decode.sv:210:21
							if (func3[2])
								// Trace: ../../rtl/VX_decode.sv:211:25
								imm[12+:5] = rs1;
							else
								// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:213:40
								rs1_r = rs1;
						end
						else begin
							// Trace: ../../rtl/VX_decode.sv:216:21
							ex_type = 3'h1;
							// Trace: ../../rtl/VX_decode.sv:217:21
							case (u_12)
								12'h000:
									// Trace: ../../rtl/VX_decode.sv:218:34
									op_type = 4'b1010;
								12'h001:
									// Trace: ../../rtl/VX_decode.sv:219:34
									op_type = 4'b1011;
								12'h002:
									// Trace: ../../rtl/VX_decode.sv:220:34
									op_type = 4'b1100;
								12'h102:
									// Trace: ../../rtl/VX_decode.sv:221:34
									op_type = 4'b1101;
								12'h302:
									// Trace: ../../rtl/VX_decode.sv:222:34
									op_type = 4'b1110;
								default:
									;
							endcase
							// Trace: ../../rtl/VX_decode.sv:225:21
							op_mod = 1;
							// Trace: ../../rtl/VX_decode.sv:226:21
							use_rd = 1;
							// Trace: ../../rtl/VX_decode.sv:227:21
							use_imm = 1;
							// Trace: ../../rtl/VX_decode.sv:228:21
							use_PC = 1;
							// Trace: ../../rtl/VX_decode.sv:229:21
							is_wstall = 1;
							// Trace: ../../rtl/VX_decode.sv:230:21
							imm = 32'd4;
							// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:231:35
							rd_r = rd;
						end
					7'b0000011: begin
						// Trace: ../../rtl/VX_decode.sv:238:17
						ex_type = 3'h2;
						// Trace: ../../rtl/VX_decode.sv:239:17
						op_type = sv2v_cast_4({1'b0, func3});
						// Trace: ../../rtl/VX_decode.sv:240:17
						use_rd = 1;
						// Trace: ../../rtl/VX_decode.sv:241:17
						imm = {{20 {u_12[11]}}, u_12};
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:247:31
						rd_r = rd;
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:248:32
						rs1_r = rs1;
					end
					7'b0100011: begin
						// Trace: ../../rtl/VX_decode.sv:254:17
						ex_type = 3'h2;
						// Trace: ../../rtl/VX_decode.sv:255:17
						op_type = sv2v_cast_4({1'b1, func3});
						// Trace: ../../rtl/VX_decode.sv:256:17
						imm = {{20 {s_imm[11]}}, s_imm};
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:257:32
						rs1_r = rs1;
						// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:263:32
						rs2_r = rs2;
					end
					7'b1101011: begin
						// Trace: ../../rtl/VX_decode.sv:354:17
						ex_type = 3'h5;
						// Trace: ../../rtl/VX_decode.sv:355:17
						case (func3)
							3'h0: begin
								// Trace: ../../rtl/VX_decode.sv:357:25
								op_type = (rs2[0] ? 4'h5 : 4'h0);
								// Trace: ../../rtl/VX_decode.sv:358:25
								is_wstall = 1;
								// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:359:40
								rs1_r = rs1;
							end
							3'h1: begin
								// Trace: ../../rtl/VX_decode.sv:362:25
								op_type = 4'h1;
								// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:363:40
								rs1_r = rs1;
								// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:364:40
								rs2_r = rs2;
							end
							3'h2: begin
								// Trace: ../../rtl/VX_decode.sv:367:25
								op_type = 4'h2;
								// Trace: ../../rtl/VX_decode.sv:368:25
								is_wstall = 1;
								// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:369:40
								rs1_r = rs1;
							end
							3'h3: begin
								// Trace: ../../rtl/VX_decode.sv:372:25
								op_type = 4'h3;
								// Trace: ../../rtl/VX_decode.sv:373:25
								is_join = 1;
							end
							3'h4: begin
								// Trace: ../../rtl/VX_decode.sv:376:25
								op_type = 4'h4;
								// Trace: ../../rtl/VX_decode.sv:377:25
								is_wstall = 1;
								// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:378:40
								rs1_r = rs1;
								// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:379:40
								rs2_r = rs2;
							end
							3'h5: begin
								// Trace: ../../rtl/VX_decode.sv:382:25
								ex_type = 3'h2;
								// Trace: ../../rtl/VX_decode.sv:383:25
								op_type = 4'b0010;
								// Trace: ../../rtl/VX_decode.sv:384:25
								op_mod = 3'sd2;
								// Trace: macro expansion of USED_IREG at ../../rtl/VX_decode.sv:385:40
								rs1_r = rs1;
							end
							default:
								;
						endcase
					end
					7'b1011011:
						// Trace: ../../rtl/VX_decode.sv:391:17
						case (func3)
							default:
								;
						endcase
					default:
						;
				endcase
			end
			// Trace: ../../rtl/VX_decode.sv:414:5
			wire wb = use_rd && |rd_r;
			// Trace: ../../rtl/VX_decode.sv:416:5
			assign VX_pipeline.decode_if.valid = VX_pipeline.ifetch_rsp_if.valid;
			// Trace: ../../rtl/VX_decode.sv:417:5
			assign VX_pipeline.decode_if.uuid = VX_pipeline.ifetch_rsp_if.uuid;
			// Trace: ../../rtl/VX_decode.sv:418:5
			assign VX_pipeline.decode_if.wid = VX_pipeline.ifetch_rsp_if.wid;
			// Trace: ../../rtl/VX_decode.sv:419:5
			assign VX_pipeline.decode_if.tmask = VX_pipeline.ifetch_rsp_if.tmask;
			// Trace: ../../rtl/VX_decode.sv:420:5
			assign VX_pipeline.decode_if.PC = VX_pipeline.ifetch_rsp_if.PC;
			// Trace: ../../rtl/VX_decode.sv:421:5
			assign VX_pipeline.decode_if.ex_type = ex_type;
			// Trace: ../../rtl/VX_decode.sv:422:5
			assign VX_pipeline.decode_if.op_type = op_type;
			// Trace: ../../rtl/VX_decode.sv:423:5
			assign VX_pipeline.decode_if.op_mod = op_mod;
			// Trace: ../../rtl/VX_decode.sv:424:5
			assign VX_pipeline.decode_if.wb = wb;
			// Trace: ../../rtl/VX_decode.sv:425:5
			assign VX_pipeline.decode_if.rd = rd_r;
			// Trace: ../../rtl/VX_decode.sv:426:5
			assign VX_pipeline.decode_if.rs1 = rs1_r;
			// Trace: ../../rtl/VX_decode.sv:427:5
			assign VX_pipeline.decode_if.rs2 = rs2_r;
			// Trace: ../../rtl/VX_decode.sv:428:5
			assign VX_pipeline.decode_if.rs3 = rs3_r;
			// Trace: ../../rtl/VX_decode.sv:429:5
			assign VX_pipeline.decode_if.imm = imm;
			// Trace: ../../rtl/VX_decode.sv:430:5
			assign VX_pipeline.decode_if.use_PC = use_PC;
			// Trace: ../../rtl/VX_decode.sv:431:5
			assign VX_pipeline.decode_if.use_imm = use_imm;
			// Trace: ../../rtl/VX_decode.sv:435:5
			wire ifetch_rsp_fire = VX_pipeline.ifetch_rsp_if.valid && VX_pipeline.ifetch_rsp_if.ready;
			// Trace: ../../rtl/VX_decode.sv:437:5
			assign VX_pipeline.join_if.valid = ifetch_rsp_fire && is_join;
			// Trace: ../../rtl/VX_decode.sv:438:5
			assign VX_pipeline.join_if.wid = VX_pipeline.ifetch_rsp_if.wid;
			// Trace: ../../rtl/VX_decode.sv:440:5
			assign VX_pipeline.wstall_if.valid = ifetch_rsp_fire;
			// Trace: ../../rtl/VX_decode.sv:441:5
			assign VX_pipeline.wstall_if.wid = VX_pipeline.ifetch_rsp_if.wid;
			// Trace: ../../rtl/VX_decode.sv:442:5
			assign VX_pipeline.wstall_if.stalled = is_wstall;
			// Trace: ../../rtl/VX_decode.sv:444:5
			assign VX_pipeline.ifetch_rsp_if.ready = VX_pipeline.decode_if.ready;
		end
	endgenerate
	assign decode.clk = clk;
	assign decode.reset = decode_reset;
	// Trace: ../../rtl/VX_pipeline.sv:177:5
	// expanded module instance: issue
	localparam _param_CF65A_CORE_ID = CORE_ID;
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	function automatic signed [1:0] sv2v_cast_2_signed;
		input reg signed [1:0] inp;
		sv2v_cast_2_signed = inp;
	endfunction
	generate
		if (1) begin : issue
			// Trace: ../../rtl/VX_issue.sv:4:15
			localparam CORE_ID = _param_CF65A_CORE_ID;
			// Trace: ../../rtl/VX_issue.sv:8:5
			wire clk;
			// Trace: ../../rtl/VX_issue.sv:9:5
			wire reset;
			// Trace: ../../rtl/VX_issue.sv:15:5
			// removed modport instance decode_if
			// Trace: ../../rtl/VX_issue.sv:16:5
			// removed modport instance writeback_if
			// Trace: ../../rtl/VX_issue.sv:18:5
			// removed modport instance alu_req_if
			// Trace: ../../rtl/VX_issue.sv:19:5
			// removed modport instance lsu_req_if
			// Trace: ../../rtl/VX_issue.sv:20:5
			// removed modport instance csr_req_if
			// Trace: ../../rtl/VX_issue.sv:24:5
			// removed modport instance gpu_req_if
			// Trace: ../../rtl/VX_issue.sv:26:5
			// expanded interface instance: ibuffer_if
			if (1) begin : ibuffer_if
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:8:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:9:5
				wire [43:0] uuid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:10:5
				wire [0:0] wid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:11:5
				wire [1:0] tmask;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:12:5
				wire [31:0] PC;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:13:5
				wire [2:0] ex_type;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:14:5
				wire [3:0] op_type;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:15:5
				wire [2:0] op_mod;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:16:5
				wire wb;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:17:5
				wire use_PC;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:18:5
				wire use_imm;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:19:5
				wire [31:0] imm;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:20:5
				wire [4:0] rd;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:21:5
				wire [4:0] rs1;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:22:5
				wire [4:0] rs2;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:23:5
				wire [4:0] rs3;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:25:5
				wire [4:0] rd_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:26:5
				wire [4:0] rs1_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:27:5
				wire [4:0] rs2_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:28:5
				wire [4:0] rs3_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:29:5
				wire [0:0] wid_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:31:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:33:5
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:58:5
			end
			// Trace: ../../rtl/VX_issue.sv:27:5
			// expanded interface instance: gpr_req_if
			if (1) begin : gpr_req_if
				// Trace: ../../rtl/interfaces/VX_gpr_req_if.sv:8:5
				wire [0:0] wid;
				// Trace: ../../rtl/interfaces/VX_gpr_req_if.sv:9:5
				wire [4:0] rs1;
				// Trace: ../../rtl/interfaces/VX_gpr_req_if.sv:10:5
				wire [4:0] rs2;
				// Trace: ../../rtl/interfaces/VX_gpr_req_if.sv:11:5
				wire [4:0] rs3;
				// Trace: ../../rtl/interfaces/VX_gpr_req_if.sv:13:5
				// Trace: ../../rtl/interfaces/VX_gpr_req_if.sv:20:5
			end
			// Trace: ../../rtl/VX_issue.sv:28:5
			// expanded interface instance: gpr_rsp_if
			if (1) begin : gpr_rsp_if
				// Trace: ../../rtl/interfaces/VX_gpr_rsp_if.sv:8:5
				wire [63:0] rs1_data;
				// Trace: ../../rtl/interfaces/VX_gpr_rsp_if.sv:9:5
				wire [63:0] rs2_data;
				// Trace: ../../rtl/interfaces/VX_gpr_rsp_if.sv:10:5
				wire [63:0] rs3_data;
				// Trace: ../../rtl/interfaces/VX_gpr_rsp_if.sv:12:5
				// Trace: ../../rtl/interfaces/VX_gpr_rsp_if.sv:18:5
			end
			// Trace: ../../rtl/VX_issue.sv:29:5
			// expanded interface instance: sboard_wb_if
			if (1) begin : sboard_wb_if
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:8:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:9:5
				wire [43:0] uuid;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:10:5
				wire [1:0] tmask;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:11:5
				wire [0:0] wid;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:12:5
				wire [31:0] PC;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:13:5
				wire [4:0] rd;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:14:5
				wire [63:0] data;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:15:5
				wire eop;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:16:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:18:5
				// Trace: ../../rtl/interfaces/VX_writeback_if.sv:30:5
			end
			// Trace: ../../rtl/VX_issue.sv:30:5
			// expanded interface instance: scoreboard_if
			if (1) begin : scoreboard_if
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:8:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:9:5
				wire [43:0] uuid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:10:5
				wire [0:0] wid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:11:5
				wire [1:0] tmask;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:12:5
				wire [31:0] PC;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:13:5
				wire [2:0] ex_type;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:14:5
				wire [3:0] op_type;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:15:5
				wire [2:0] op_mod;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:16:5
				wire wb;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:17:5
				wire use_PC;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:18:5
				wire use_imm;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:19:5
				wire [31:0] imm;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:20:5
				wire [4:0] rd;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:21:5
				wire [4:0] rs1;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:22:5
				wire [4:0] rs2;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:23:5
				wire [4:0] rs3;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:25:5
				wire [4:0] rd_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:26:5
				wire [4:0] rs1_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:27:5
				wire [4:0] rs2_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:28:5
				wire [4:0] rs3_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:29:5
				wire [0:0] wid_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:31:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:33:5
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:58:5
			end
			// Trace: ../../rtl/VX_issue.sv:31:5
			// expanded interface instance: dispatch_if
			if (1) begin : dispatch_if
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:8:5
				wire valid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:9:5
				wire [43:0] uuid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:10:5
				wire [0:0] wid;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:11:5
				wire [1:0] tmask;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:12:5
				wire [31:0] PC;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:13:5
				wire [2:0] ex_type;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:14:5
				wire [3:0] op_type;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:15:5
				wire [2:0] op_mod;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:16:5
				wire wb;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:17:5
				wire use_PC;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:18:5
				wire use_imm;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:19:5
				wire [31:0] imm;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:20:5
				wire [4:0] rd;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:21:5
				wire [4:0] rs1;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:22:5
				wire [4:0] rs2;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:23:5
				wire [4:0] rs3;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:25:5
				wire [4:0] rd_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:26:5
				wire [4:0] rs1_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:27:5
				wire [4:0] rs2_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:28:5
				wire [4:0] rs3_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:29:5
				wire [0:0] wid_n;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:31:5
				wire ready;
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:33:5
				// Trace: ../../rtl/interfaces/VX_ibuffer_if.sv:58:5
			end
			// Trace: ../../rtl/VX_issue.sv:34:5
			assign gpr_req_if.wid = ibuffer_if.wid;
			// Trace: ../../rtl/VX_issue.sv:35:5
			assign gpr_req_if.rs1 = ibuffer_if.rs1;
			// Trace: ../../rtl/VX_issue.sv:36:5
			assign gpr_req_if.rs2 = ibuffer_if.rs2;
			// Trace: ../../rtl/VX_issue.sv:37:5
			assign gpr_req_if.rs3 = ibuffer_if.rs3;
			// Trace: ../../rtl/VX_issue.sv:40:5
			assign sboard_wb_if.valid = VX_pipeline.writeback_if.valid;
			// Trace: ../../rtl/VX_issue.sv:41:5
			assign sboard_wb_if.uuid = VX_pipeline.writeback_if.uuid;
			// Trace: ../../rtl/VX_issue.sv:42:5
			assign sboard_wb_if.wid = VX_pipeline.writeback_if.wid;
			// Trace: ../../rtl/VX_issue.sv:43:5
			assign sboard_wb_if.PC = VX_pipeline.writeback_if.PC;
			// Trace: ../../rtl/VX_issue.sv:44:5
			assign sboard_wb_if.rd = VX_pipeline.writeback_if.rd;
			// Trace: ../../rtl/VX_issue.sv:45:5
			assign sboard_wb_if.eop = VX_pipeline.writeback_if.eop;
			// Trace: ../../rtl/VX_issue.sv:48:5
			assign scoreboard_if.valid = ibuffer_if.valid && dispatch_if.ready;
			// Trace: ../../rtl/VX_issue.sv:49:5
			assign scoreboard_if.uuid = ibuffer_if.uuid;
			// Trace: ../../rtl/VX_issue.sv:50:5
			assign scoreboard_if.wid = ibuffer_if.wid;
			// Trace: ../../rtl/VX_issue.sv:51:5
			assign scoreboard_if.PC = ibuffer_if.PC;
			// Trace: ../../rtl/VX_issue.sv:52:5
			assign scoreboard_if.wb = ibuffer_if.wb;
			// Trace: ../../rtl/VX_issue.sv:53:5
			assign scoreboard_if.rd = ibuffer_if.rd;
			// Trace: ../../rtl/VX_issue.sv:54:5
			assign scoreboard_if.rd_n = ibuffer_if.rd_n;
			// Trace: ../../rtl/VX_issue.sv:55:5
			assign scoreboard_if.rs1_n = ibuffer_if.rs1_n;
			// Trace: ../../rtl/VX_issue.sv:56:5
			assign scoreboard_if.rs2_n = ibuffer_if.rs2_n;
			// Trace: ../../rtl/VX_issue.sv:57:5
			assign scoreboard_if.rs3_n = ibuffer_if.rs3_n;
			// Trace: ../../rtl/VX_issue.sv:58:5
			assign scoreboard_if.wid_n = ibuffer_if.wid_n;
			// Trace: ../../rtl/VX_issue.sv:61:5
			assign dispatch_if.valid = ibuffer_if.valid && scoreboard_if.ready;
			// Trace: ../../rtl/VX_issue.sv:62:5
			assign dispatch_if.uuid = ibuffer_if.uuid;
			// Trace: ../../rtl/VX_issue.sv:63:5
			assign dispatch_if.wid = ibuffer_if.wid;
			// Trace: ../../rtl/VX_issue.sv:64:5
			assign dispatch_if.tmask = ibuffer_if.tmask;
			// Trace: ../../rtl/VX_issue.sv:65:5
			assign dispatch_if.PC = ibuffer_if.PC;
			// Trace: ../../rtl/VX_issue.sv:66:5
			assign dispatch_if.ex_type = ibuffer_if.ex_type;
			// Trace: ../../rtl/VX_issue.sv:67:5
			assign dispatch_if.op_type = ibuffer_if.op_type;
			// Trace: ../../rtl/VX_issue.sv:68:5
			assign dispatch_if.op_mod = ibuffer_if.op_mod;
			// Trace: ../../rtl/VX_issue.sv:69:5
			assign dispatch_if.wb = ibuffer_if.wb;
			// Trace: ../../rtl/VX_issue.sv:70:5
			assign dispatch_if.rd = ibuffer_if.rd;
			// Trace: ../../rtl/VX_issue.sv:71:5
			assign dispatch_if.rs1 = ibuffer_if.rs1;
			// Trace: ../../rtl/VX_issue.sv:72:5
			assign dispatch_if.imm = ibuffer_if.imm;
			// Trace: ../../rtl/VX_issue.sv:73:5
			assign dispatch_if.use_PC = ibuffer_if.use_PC;
			// Trace: ../../rtl/VX_issue.sv:74:5
			assign dispatch_if.use_imm = ibuffer_if.use_imm;
			// Trace: ../../rtl/VX_issue.sv:77:5
			assign ibuffer_if.ready = scoreboard_if.ready && dispatch_if.ready;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_issue.sv:79:23
			wire ibuf_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_issue.sv:79:56
			VX_reset_relay __ibuf_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(ibuf_reset)
			);
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_issue.sv:80:29
			wire scoreboard_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_issue.sv:80:62
			VX_reset_relay __scoreboard_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(scoreboard_reset)
			);
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_issue.sv:81:22
			wire gpr_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_issue.sv:81:55
			VX_reset_relay __gpr_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(gpr_reset)
			);
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_issue.sv:82:27
			wire dispatch_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_issue.sv:82:60
			VX_reset_relay __dispatch_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(dispatch_reset)
			);
			// Trace: ../../rtl/VX_issue.sv:84:5
			// expanded module instance: ibuffer
			localparam _param_D579A_CORE_ID = CORE_ID;
			if (1) begin : ibuffer
				// Trace: ../../rtl/VX_ibuffer.sv:4:15
				localparam CORE_ID = _param_D579A_CORE_ID;
				// Trace: ../../rtl/VX_ibuffer.sv:6:5
				wire clk;
				// Trace: ../../rtl/VX_ibuffer.sv:7:5
				wire reset;
				// Trace: ../../rtl/VX_ibuffer.sv:10:5
				// removed modport instance decode_if
				// Trace: ../../rtl/VX_ibuffer.sv:13:5
				// removed modport instance ibuffer_if
				// Trace: ../../rtl/VX_ibuffer.sv:18:5
				localparam DATAW = 143;
				// Trace: ../../rtl/VX_ibuffer.sv:19:5
				localparam ADDRW = 2;
				// Trace: ../../rtl/VX_ibuffer.sv:20:5
				localparam NWARPSW = 2;
				// Trace: ../../rtl/VX_ibuffer.sv:22:5
				reg [3:0] used_r;
				// Trace: ../../rtl/VX_ibuffer.sv:23:5
				reg [1:0] full_r;
				reg [1:0] empty_r;
				reg [1:0] alm_empty_r;
				// Trace: ../../rtl/VX_ibuffer.sv:25:5
				wire [1:0] q_full;
				wire [1:0] q_empty;
				wire [1:0] q_alm_empty;
				// Trace: ../../rtl/VX_ibuffer.sv:26:5
				wire [142:0] q_data_in;
				// Trace: ../../rtl/VX_ibuffer.sv:27:5
				wire [285:0] q_data_prev;
				// Trace: ../../rtl/VX_ibuffer.sv:28:5
				reg [285:0] q_data_out;
				// Trace: ../../rtl/VX_ibuffer.sv:30:5
				wire enq_fire = VX_pipeline.decode_if.valid && VX_pipeline.decode_if.ready;
				// Trace: ../../rtl/VX_ibuffer.sv:31:5
				wire deq_fire = VX_pipeline.issue.ibuffer_if.valid && VX_pipeline.issue.ibuffer_if.ready;
				// Trace: ../../rtl/VX_ibuffer.sv:33:5
				genvar i;
				for (i = 0; i < 2; i = i + 1) begin : genblk1
					// Trace: ../../rtl/VX_ibuffer.sv:35:9
					wire writing = enq_fire && (i == VX_pipeline.decode_if.wid);
					// Trace: ../../rtl/VX_ibuffer.sv:36:9
					wire reading = deq_fire && (i == VX_pipeline.issue.ibuffer_if.wid);
					// Trace: ../../rtl/VX_ibuffer.sv:38:9
					wire going_empty = empty_r[i] || (alm_empty_r[i] && reading);
					// Trace: ../../rtl/VX_ibuffer.sv:40:9
					VX_elastic_buffer #(
						.DATAW(DATAW),
						.SIZE(2),
						.OUT_REG(1)
					) queue(
						.clk(clk),
						.reset(reset),
						.valid_in(writing && !going_empty),
						.data_in(q_data_in),
						.ready_out(reading),
						.data_out(q_data_prev[i * 143+:143])
					);
					// Trace: ../../rtl/VX_ibuffer.sv:55:9
					always @(posedge clk) begin
						// Trace: ../../rtl/VX_ibuffer.sv:56:13
						if (reset) begin
							// Trace: ../../rtl/VX_ibuffer.sv:57:17
							used_r[i * 2+:2] <= 0;
							// Trace: ../../rtl/VX_ibuffer.sv:58:17
							full_r[i] <= 0;
							// Trace: ../../rtl/VX_ibuffer.sv:59:17
							empty_r[i] <= 1;
							// Trace: ../../rtl/VX_ibuffer.sv:60:17
							alm_empty_r[i] <= 1;
						end
						else begin
							// Trace: ../../rtl/VX_ibuffer.sv:62:17
							if (writing) begin
								begin
									// Trace: ../../rtl/VX_ibuffer.sv:63:21
									if (!reading) begin
										// Trace: ../../rtl/VX_ibuffer.sv:64:25
										empty_r[i] <= 0;
										// Trace: ../../rtl/VX_ibuffer.sv:65:25
										if (used_r[i * 2+:2] == 1)
											// Trace: ../../rtl/VX_ibuffer.sv:66:29
											alm_empty_r[i] <= 0;
										if (used_r[i * 2+:2] == 2'sd2)
											// Trace: ../../rtl/VX_ibuffer.sv:68:29
											full_r[i] <= 1;
									end
								end
							end
							else if (reading) begin
								// Trace: ../../rtl/VX_ibuffer.sv:71:21
								full_r[i] <= 0;
								// Trace: ../../rtl/VX_ibuffer.sv:72:21
								if (used_r[i * 2+:2] == 2'sd1)
									// Trace: ../../rtl/VX_ibuffer.sv:73:25
									empty_r[i] <= 1;
								if (used_r[i * 2+:2] == 2'sd2)
									// Trace: ../../rtl/VX_ibuffer.sv:75:25
									alm_empty_r[i] <= 1;
							end
							// Trace: ../../rtl/VX_ibuffer.sv:77:17
							used_r[i * 2+:2] <= used_r[i * 2+:2] + sv2v_cast_2_signed($signed(sv2v_cast_2(writing) - sv2v_cast_2(reading)));
						end
						if (writing && going_empty)
							// Trace: ../../rtl/VX_ibuffer.sv:81:17
							q_data_out[i * 143+:143] <= q_data_in;
						else if (reading)
							// Trace: ../../rtl/VX_ibuffer.sv:83:17
							q_data_out[i * 143+:143] <= q_data_prev[i * 143+:143];
					end
					// Trace: ../../rtl/VX_ibuffer.sv:87:9
					assign q_full[i] = full_r[i];
					// Trace: ../../rtl/VX_ibuffer.sv:88:9
					assign q_empty[i] = empty_r[i];
					// Trace: ../../rtl/VX_ibuffer.sv:89:9
					assign q_alm_empty[i] = alm_empty_r[i];
				end
				// Trace: ../../rtl/VX_ibuffer.sv:94:5
				reg [1:0] valid_table;
				reg [1:0] valid_table_n;
				// Trace: ../../rtl/VX_ibuffer.sv:95:5
				reg [0:0] deq_wid;
				reg [0:0] deq_wid_n;
				// Trace: ../../rtl/VX_ibuffer.sv:96:5
				reg [0:0] deq_wid_rr;
				reg [0:0] deq_wid_rr_n;
				// Trace: ../../rtl/VX_ibuffer.sv:97:5
				reg deq_valid;
				reg deq_valid_n;
				// Trace: ../../rtl/VX_ibuffer.sv:98:5
				reg [142:0] deq_instr;
				reg [142:0] deq_instr_n;
				// Trace: ../../rtl/VX_ibuffer.sv:99:5
				reg [1:0] num_warps;
				// Trace: ../../rtl/VX_ibuffer.sv:104:5
				always @(*) begin
					// Trace: ../../rtl/VX_ibuffer.sv:105:9
					valid_table_n = valid_table;
					// Trace: ../../rtl/VX_ibuffer.sv:106:9
					if (deq_fire)
						// Trace: ../../rtl/VX_ibuffer.sv:107:13
						valid_table_n[deq_wid] = !q_alm_empty[deq_wid];
					if (enq_fire)
						// Trace: ../../rtl/VX_ibuffer.sv:110:13
						valid_table_n[VX_pipeline.decode_if.wid] = 1;
				end
				// Trace: ../../rtl/VX_ibuffer.sv:115:5
				// rewrote reg-to-output bindings
				wire [1:1] sv2v_tmp_rr_arbiter_grant_index;
				always @(*) deq_wid_rr_n = sv2v_tmp_rr_arbiter_grant_index;
				VX_rr_arbiter #(.NUM_REQS(2)) rr_arbiter(
					.clk(clk),
					.reset(reset),
					.requests(valid_table_n),
					.grant_index(sv2v_tmp_rr_arbiter_grant_index)
				);
				// Trace: ../../rtl/VX_ibuffer.sv:128:5
				always @(*)
					// Trace: ../../rtl/VX_ibuffer.sv:129:9
					if (num_warps > 1) begin
						// Trace: ../../rtl/VX_ibuffer.sv:130:13
						deq_valid_n = 1;
						// Trace: ../../rtl/VX_ibuffer.sv:131:13
						deq_wid_n = deq_wid_rr;
						// Trace: ../../rtl/VX_ibuffer.sv:132:13
						deq_instr_n = q_data_out[deq_wid_rr * 143+:143];
					end
					else if ((1 == num_warps) && !(deq_fire && q_alm_empty[deq_wid])) begin
						// Trace: ../../rtl/VX_ibuffer.sv:134:13
						deq_valid_n = 1;
						// Trace: ../../rtl/VX_ibuffer.sv:135:13
						deq_wid_n = deq_wid;
						// Trace: ../../rtl/VX_ibuffer.sv:136:13
						deq_instr_n = (deq_fire ? q_data_prev[deq_wid * 143+:143] : q_data_out[deq_wid * 143+:143]);
					end
					else begin
						// Trace: ../../rtl/VX_ibuffer.sv:138:13
						deq_valid_n = enq_fire;
						// Trace: ../../rtl/VX_ibuffer.sv:139:13
						deq_wid_n = VX_pipeline.decode_if.wid;
						// Trace: ../../rtl/VX_ibuffer.sv:140:13
						deq_instr_n = q_data_in;
					end
				// Trace: ../../rtl/VX_ibuffer.sv:144:5
				wire warp_added = enq_fire && q_empty[VX_pipeline.decode_if.wid];
				// Trace: ../../rtl/VX_ibuffer.sv:145:5
				wire warp_removed = (deq_fire && ~(enq_fire && (VX_pipeline.decode_if.wid == deq_wid))) && q_alm_empty[deq_wid];
				// Trace: ../../rtl/VX_ibuffer.sv:147:5
				always @(posedge clk) begin
					// Trace: ../../rtl/VX_ibuffer.sv:148:9
					if (reset) begin
						// Trace: ../../rtl/VX_ibuffer.sv:149:13
						valid_table <= 0;
						// Trace: ../../rtl/VX_ibuffer.sv:150:13
						deq_valid <= 0;
						// Trace: ../../rtl/VX_ibuffer.sv:151:13
						num_warps <= 0;
					end
					else begin
						// Trace: ../../rtl/VX_ibuffer.sv:153:13
						valid_table <= valid_table_n;
						// Trace: ../../rtl/VX_ibuffer.sv:154:13
						deq_valid <= deq_valid_n;
						// Trace: ../../rtl/VX_ibuffer.sv:157:13
						if (warp_added && !warp_removed)
							// Trace: ../../rtl/VX_ibuffer.sv:158:17
							num_warps <= num_warps + 2'sd1;
						else if (warp_removed && !warp_added)
							// Trace: ../../rtl/VX_ibuffer.sv:160:17
							num_warps <= num_warps - 2'sd1;
					end
					// Trace: ../../rtl/VX_ibuffer.sv:164:9
					deq_wid <= deq_wid_n;
					// Trace: ../../rtl/VX_ibuffer.sv:165:9
					deq_wid_rr <= deq_wid_rr_n;
					// Trace: ../../rtl/VX_ibuffer.sv:166:9
					deq_instr <= deq_instr_n;
				end
				// Trace: ../../rtl/VX_ibuffer.sv:169:5
				assign VX_pipeline.decode_if.ready = ~q_full[VX_pipeline.decode_if.wid];
				// Trace: ../../rtl/VX_ibuffer.sv:171:5
				assign q_data_in = {VX_pipeline.decode_if.uuid, VX_pipeline.decode_if.tmask, VX_pipeline.decode_if.PC, VX_pipeline.decode_if.ex_type, VX_pipeline.decode_if.op_type, VX_pipeline.decode_if.op_mod, VX_pipeline.decode_if.wb, VX_pipeline.decode_if.use_PC, VX_pipeline.decode_if.use_imm, VX_pipeline.decode_if.imm, VX_pipeline.decode_if.rd, VX_pipeline.decode_if.rs1, VX_pipeline.decode_if.rs2, VX_pipeline.decode_if.rs3};
				// Trace: ../../rtl/VX_ibuffer.sv:186:5
				assign VX_pipeline.issue.ibuffer_if.valid = deq_valid;
				// Trace: ../../rtl/VX_ibuffer.sv:187:5
				assign VX_pipeline.issue.ibuffer_if.wid = deq_wid;
				// Trace: ../../rtl/VX_ibuffer.sv:188:5
				assign {VX_pipeline.issue.ibuffer_if.uuid, VX_pipeline.issue.ibuffer_if.tmask, VX_pipeline.issue.ibuffer_if.PC, VX_pipeline.issue.ibuffer_if.ex_type, VX_pipeline.issue.ibuffer_if.op_type, VX_pipeline.issue.ibuffer_if.op_mod, VX_pipeline.issue.ibuffer_if.wb, VX_pipeline.issue.ibuffer_if.use_PC, VX_pipeline.issue.ibuffer_if.use_imm, VX_pipeline.issue.ibuffer_if.imm, VX_pipeline.issue.ibuffer_if.rd, VX_pipeline.issue.ibuffer_if.rs1, VX_pipeline.issue.ibuffer_if.rs2, VX_pipeline.issue.ibuffer_if.rs3} = deq_instr;
				// Trace: ../../rtl/VX_ibuffer.sv:204:5
				assign VX_pipeline.issue.ibuffer_if.wid_n = deq_wid_n;
				// Trace: ../../rtl/VX_ibuffer.sv:205:5
				assign VX_pipeline.issue.ibuffer_if.rd_n = deq_instr_n[15+:5];
				// Trace: ../../rtl/VX_ibuffer.sv:206:5
				assign VX_pipeline.issue.ibuffer_if.rs1_n = deq_instr_n[10+:5];
				// Trace: ../../rtl/VX_ibuffer.sv:207:5
				assign VX_pipeline.issue.ibuffer_if.rs2_n = deq_instr_n[5+:5];
				// Trace: ../../rtl/VX_ibuffer.sv:208:5
				assign VX_pipeline.issue.ibuffer_if.rs3_n = deq_instr_n[0+:5];
			end
			assign ibuffer.clk = clk;
			assign ibuffer.reset = ibuf_reset;
			// Trace: ../../rtl/VX_issue.sv:93:5
			// expanded module instance: scoreboard
			localparam _param_85D2C_CORE_ID = CORE_ID;
			if (1) begin : scoreboard
				// Trace: ../../rtl/VX_scoreboard.sv:4:15
				localparam CORE_ID = _param_85D2C_CORE_ID;
				// Trace: ../../rtl/VX_scoreboard.sv:6:5
				wire clk;
				// Trace: ../../rtl/VX_scoreboard.sv:7:5
				wire reset;
				// Trace: ../../rtl/VX_scoreboard.sv:9:5
				// removed modport instance ibuffer_if
				// Trace: ../../rtl/VX_scoreboard.sv:10:5
				// removed modport instance writeback_if
				// Trace: ../../rtl/VX_scoreboard.sv:12:5
				reg [63:0] inuse_regs;
				reg [63:0] inuse_regs_n;
				// Trace: ../../rtl/VX_scoreboard.sv:14:5
				wire reserve_reg = (VX_pipeline.issue.scoreboard_if.valid && VX_pipeline.issue.scoreboard_if.ready) && VX_pipeline.issue.scoreboard_if.wb;
				// Trace: ../../rtl/VX_scoreboard.sv:16:5
				wire release_reg = (VX_pipeline.issue.sboard_wb_if.valid && VX_pipeline.issue.sboard_wb_if.ready) && VX_pipeline.issue.sboard_wb_if.eop;
				// Trace: ../../rtl/VX_scoreboard.sv:18:5
				always @(*) begin
					// Trace: ../../rtl/VX_scoreboard.sv:19:9
					inuse_regs_n = inuse_regs;
					// Trace: ../../rtl/VX_scoreboard.sv:20:9
					if (reserve_reg)
						// Trace: ../../rtl/VX_scoreboard.sv:21:13
						inuse_regs_n[(VX_pipeline.issue.scoreboard_if.wid * 32) + VX_pipeline.issue.scoreboard_if.rd] = 1;
					if (release_reg)
						// Trace: ../../rtl/VX_scoreboard.sv:24:13
						inuse_regs_n[(VX_pipeline.issue.sboard_wb_if.wid * 32) + VX_pipeline.issue.sboard_wb_if.rd] = 0;
				end
				// Trace: ../../rtl/VX_scoreboard.sv:28:5
				always @(posedge clk)
					// Trace: ../../rtl/VX_scoreboard.sv:29:9
					if (reset)
						// Trace: ../../rtl/VX_scoreboard.sv:30:13
						inuse_regs <= 1'sb0;
					else
						// Trace: ../../rtl/VX_scoreboard.sv:32:13
						inuse_regs <= inuse_regs_n;
				// Trace: ../../rtl/VX_scoreboard.sv:36:5
				reg deq_inuse_rd;
				reg deq_inuse_rs1;
				reg deq_inuse_rs2;
				reg deq_inuse_rs3;
				// Trace: ../../rtl/VX_scoreboard.sv:38:5
				always @(posedge clk) begin
					// Trace: ../../rtl/VX_scoreboard.sv:39:9
					deq_inuse_rd <= inuse_regs_n[(VX_pipeline.issue.scoreboard_if.wid_n * 32) + VX_pipeline.issue.scoreboard_if.rd_n];
					// Trace: ../../rtl/VX_scoreboard.sv:40:9
					deq_inuse_rs1 <= inuse_regs_n[(VX_pipeline.issue.scoreboard_if.wid_n * 32) + VX_pipeline.issue.scoreboard_if.rs1_n];
					// Trace: ../../rtl/VX_scoreboard.sv:41:9
					deq_inuse_rs2 <= inuse_regs_n[(VX_pipeline.issue.scoreboard_if.wid_n * 32) + VX_pipeline.issue.scoreboard_if.rs2_n];
					// Trace: ../../rtl/VX_scoreboard.sv:42:9
					deq_inuse_rs3 <= inuse_regs_n[(VX_pipeline.issue.scoreboard_if.wid_n * 32) + VX_pipeline.issue.scoreboard_if.rs3_n];
				end
				// Trace: ../../rtl/VX_scoreboard.sv:45:5
				assign VX_pipeline.issue.sboard_wb_if.ready = 1'b1;
				// Trace: ../../rtl/VX_scoreboard.sv:47:5
				assign VX_pipeline.issue.scoreboard_if.ready = ~(((deq_inuse_rd | deq_inuse_rs1) | deq_inuse_rs2) | deq_inuse_rs3);
				// Trace: ../../rtl/VX_scoreboard.sv:54:5
				reg [31:0] deadlock_ctr;
				// Trace: ../../rtl/VX_scoreboard.sv:55:5
				wire [31:0] deadlock_timeout = 10000;
				// Trace: ../../rtl/VX_scoreboard.sv:57:5
				always @(posedge clk)
					// Trace: ../../rtl/VX_scoreboard.sv:58:9
					if (reset)
						// Trace: ../../rtl/VX_scoreboard.sv:59:13
						deadlock_ctr <= 0;
					else begin
						// Trace: ../../rtl/VX_scoreboard.sv:68:13
						if (release_reg)
							// Trace: macro expansion of ASSERT at ../../rtl/VX_scoreboard.sv:71:112
							if (inuse_regs[(VX_pipeline.issue.sboard_wb_if.wid * 32) + VX_pipeline.issue.sboard_wb_if.rd] != 0)
								;
						if (VX_pipeline.issue.scoreboard_if.valid && ~VX_pipeline.issue.scoreboard_if.ready) begin
							// Trace: ../../rtl/VX_scoreboard.sv:74:17
							deadlock_ctr <= deadlock_ctr + 1;
							// Trace: macro expansion of ASSERT at ../../rtl/VX_scoreboard.sv:78:94
							if (deadlock_ctr < deadlock_timeout)
								;
						end
						else if (VX_pipeline.issue.scoreboard_if.valid && VX_pipeline.issue.scoreboard_if.ready)
							// Trace: ../../rtl/VX_scoreboard.sv:80:17
							deadlock_ctr <= 0;
					end
			end
			assign scoreboard.clk = clk;
			assign scoreboard.reset = scoreboard_reset;
			// Trace: ../../rtl/VX_issue.sv:102:5
			// expanded module instance: gpr_stage
			localparam _param_E2C9E_CORE_ID = CORE_ID;
			if (1) begin : gpr_stage
				// Trace: ../../rtl/VX_gpr_stage.sv:4:15
				localparam CORE_ID = _param_E2C9E_CORE_ID;
				// Trace: ../../rtl/VX_gpr_stage.sv:6:5
				wire clk;
				// Trace: ../../rtl/VX_gpr_stage.sv:7:5
				wire reset;
				// Trace: ../../rtl/VX_gpr_stage.sv:10:5
				// removed modport instance writeback_if
				// Trace: ../../rtl/VX_gpr_stage.sv:11:5
				// removed modport instance gpr_req_if
				// Trace: ../../rtl/VX_gpr_stage.sv:14:5
				// removed modport instance gpr_rsp_if
				// Trace: ../../rtl/VX_gpr_stage.sv:20:5
				localparam RAM_SIZE = 64;
				// Trace: ../../rtl/VX_gpr_stage.sv:23:5
				wire write_enable = VX_pipeline.writeback_if.valid && (VX_pipeline.writeback_if.rd != 0);
				// Trace: ../../rtl/VX_gpr_stage.sv:25:5
				wire [1:0] wren;
				// Trace: ../../rtl/VX_gpr_stage.sv:26:5
				genvar i;
				for (i = 0; i < 2; i = i + 1) begin : genblk1
					// Trace: ../../rtl/VX_gpr_stage.sv:27:9
					assign wren[i] = write_enable && VX_pipeline.writeback_if.tmask[i];
				end
				// Trace: ../../rtl/VX_gpr_stage.sv:30:5
				wire [5:0] waddr;
				wire [5:0] raddr1;
				wire [5:0] raddr2;
				// Trace: ../../rtl/VX_gpr_stage.sv:31:5
				assign waddr = {VX_pipeline.writeback_if.wid, VX_pipeline.writeback_if.rd};
				// Trace: ../../rtl/VX_gpr_stage.sv:32:5
				assign raddr1 = {VX_pipeline.issue.gpr_req_if.wid, VX_pipeline.issue.gpr_req_if.rs1};
				// Trace: ../../rtl/VX_gpr_stage.sv:33:5
				assign raddr2 = {VX_pipeline.issue.gpr_req_if.wid, VX_pipeline.issue.gpr_req_if.rs2};
				// Trace: ../../rtl/VX_gpr_stage.sv:35:5
				for (i = 0; i < 2; i = i + 1) begin : genblk2
					// Trace: ../../rtl/VX_gpr_stage.sv:36:9
					VX_dp_ram #(
						.DATAW(32),
						.SIZE(RAM_SIZE),
						.INIT_ENABLE(1),
						.INIT_VALUE(0)
					) dp_ram1(
						.clk(clk),
						.wren(wren[i]),
						.waddr(waddr),
						.wdata(VX_pipeline.writeback_if.data[i * 32+:32]),
						.raddr(raddr1),
						.rdata(VX_pipeline.issue.gpr_rsp_if.rs1_data[i * 32+:32])
					);
					// Trace: ../../rtl/VX_gpr_stage.sv:50:9
					VX_dp_ram #(
						.DATAW(32),
						.SIZE(RAM_SIZE),
						.INIT_ENABLE(1),
						.INIT_VALUE(0)
					) dp_ram2(
						.clk(clk),
						.wren(wren[i]),
						.waddr(waddr),
						.wdata(VX_pipeline.writeback_if.data[i * 32+:32]),
						.raddr(raddr2),
						.rdata(VX_pipeline.issue.gpr_rsp_if.rs2_data[i * 32+:32])
					);
				end
				// Trace: ../../rtl/VX_gpr_stage.sv:86:5
				assign VX_pipeline.issue.gpr_rsp_if.rs3_data = 1'sbx;
				// Trace: ../../rtl/VX_gpr_stage.sv:89:5
				assign VX_pipeline.writeback_if.ready = 1'b1;
			end
			assign gpr_stage.clk = clk;
			assign gpr_stage.reset = gpr_reset;
			// Trace: ../../rtl/VX_issue.sv:112:5
			// expanded module instance: dispatch
			if (1) begin : dispatch
				// Trace: ../../rtl/VX_dispatch.sv:4:5
				wire clk;
				// Trace: ../../rtl/VX_dispatch.sv:5:5
				wire reset;
				// Trace: ../../rtl/VX_dispatch.sv:8:5
				// removed modport instance ibuffer_if
				// Trace: ../../rtl/VX_dispatch.sv:9:5
				// removed modport instance gpr_rsp_if
				// Trace: ../../rtl/VX_dispatch.sv:12:5
				// removed modport instance alu_req_if
				// Trace: ../../rtl/VX_dispatch.sv:13:5
				// removed modport instance lsu_req_if
				// Trace: ../../rtl/VX_dispatch.sv:14:5
				// removed modport instance csr_req_if
				// Trace: ../../rtl/VX_dispatch.sv:18:5
				// removed modport instance gpu_req_if
				// Trace: ../../rtl/VX_dispatch.sv:20:5
				wire [0:0] tid;
				// Trace: ../../rtl/VX_dispatch.sv:21:5
				wire alu_req_ready;
				// Trace: ../../rtl/VX_dispatch.sv:22:5
				wire lsu_req_ready;
				// Trace: ../../rtl/VX_dispatch.sv:23:5
				wire csr_req_ready;
				// Trace: ../../rtl/VX_dispatch.sv:27:5
				wire gpu_req_ready;
				// Trace: ../../rtl/VX_dispatch.sv:29:5
				VX_lzc #(.N(2)) tid_select(
					.in_i(VX_pipeline.issue.dispatch_if.tmask),
					.cnt_o(tid)
				);
				// Trace: ../../rtl/VX_dispatch.sv:37:5
				wire [31:0] next_PC = VX_pipeline.issue.dispatch_if.PC + 4;
				// Trace: ../../rtl/VX_dispatch.sv:41:5
				wire alu_req_valid = VX_pipeline.issue.dispatch_if.valid && (VX_pipeline.issue.dispatch_if.ex_type == 3'h1);
				// Trace: ../../rtl/VX_dispatch.sv:42:5
				wire [3:0] alu_op_type = VX_pipeline.issue.dispatch_if.op_type;
				// Trace: ../../rtl/VX_dispatch.sv:44:5
				VX_skid_buffer #(
					.DATAW(287),
					.OUT_REG(1)
				) alu_buffer(
					.clk(clk),
					.reset(reset),
					.valid_in(alu_req_valid),
					.ready_in(alu_req_ready),
					.data_in({VX_pipeline.issue.dispatch_if.uuid, VX_pipeline.issue.dispatch_if.wid, VX_pipeline.issue.dispatch_if.tmask, VX_pipeline.issue.dispatch_if.PC, next_PC, alu_op_type, VX_pipeline.issue.dispatch_if.op_mod, VX_pipeline.issue.dispatch_if.imm, VX_pipeline.issue.dispatch_if.use_PC, VX_pipeline.issue.dispatch_if.use_imm, VX_pipeline.issue.dispatch_if.rd, VX_pipeline.issue.dispatch_if.wb, tid, VX_pipeline.issue.gpr_rsp_if.rs1_data, VX_pipeline.issue.gpr_rsp_if.rs2_data}),
					.data_out({VX_pipeline.alu_req_if.uuid, VX_pipeline.alu_req_if.wid, VX_pipeline.alu_req_if.tmask, VX_pipeline.alu_req_if.PC, VX_pipeline.alu_req_if.next_PC, VX_pipeline.alu_req_if.op_type, VX_pipeline.alu_req_if.op_mod, VX_pipeline.alu_req_if.imm, VX_pipeline.alu_req_if.use_PC, VX_pipeline.alu_req_if.use_imm, VX_pipeline.alu_req_if.rd, VX_pipeline.alu_req_if.wb, VX_pipeline.alu_req_if.tid, VX_pipeline.alu_req_if.rs1_data, VX_pipeline.alu_req_if.rs2_data}),
					.valid_out(VX_pipeline.alu_req_if.valid),
					.ready_out(VX_pipeline.alu_req_if.ready)
				);
				// Trace: ../../rtl/VX_dispatch.sv:60:5
				wire lsu_req_valid = VX_pipeline.issue.dispatch_if.valid && (VX_pipeline.issue.dispatch_if.ex_type == 3'h2);
				// Trace: ../../rtl/VX_dispatch.sv:61:5
				wire [3:0] lsu_op_type = VX_pipeline.issue.dispatch_if.op_type;
				// Trace: ../../rtl/VX_dispatch.sv:62:5
				wire lsu_is_fence = 3'h1 == VX_pipeline.issue.dispatch_if.op_mod;
				// Trace: ../../rtl/VX_dispatch.sv:63:5
				wire lsu_is_prefetch = 3'h2 == VX_pipeline.issue.dispatch_if.op_mod;
				// Trace: ../../rtl/VX_dispatch.sv:65:5
				VX_skid_buffer #(
					.DATAW(251),
					.OUT_REG(1)
				) lsu_buffer(
					.clk(clk),
					.reset(reset),
					.valid_in(lsu_req_valid),
					.ready_in(lsu_req_ready),
					.data_in({VX_pipeline.issue.dispatch_if.uuid, VX_pipeline.issue.dispatch_if.wid, VX_pipeline.issue.dispatch_if.tmask, VX_pipeline.issue.dispatch_if.PC, lsu_op_type, lsu_is_fence, VX_pipeline.issue.dispatch_if.imm, VX_pipeline.issue.dispatch_if.rd, VX_pipeline.issue.dispatch_if.wb, VX_pipeline.issue.gpr_rsp_if.rs1_data, VX_pipeline.issue.gpr_rsp_if.rs2_data, lsu_is_prefetch}),
					.data_out({VX_pipeline.lsu_req_if.uuid, VX_pipeline.lsu_req_if.wid, VX_pipeline.lsu_req_if.tmask, VX_pipeline.lsu_req_if.PC, VX_pipeline.lsu_req_if.op_type, VX_pipeline.lsu_req_if.is_fence, VX_pipeline.lsu_req_if.offset, VX_pipeline.lsu_req_if.rd, VX_pipeline.lsu_req_if.wb, VX_pipeline.lsu_req_if.base_addr, VX_pipeline.lsu_req_if.store_data, VX_pipeline.lsu_req_if.is_prefetch}),
					.valid_out(VX_pipeline.lsu_req_if.valid),
					.ready_out(VX_pipeline.lsu_req_if.ready)
				);
				// Trace: ../../rtl/VX_dispatch.sv:81:5
				wire csr_req_valid = VX_pipeline.issue.dispatch_if.valid && (VX_pipeline.issue.dispatch_if.ex_type == 3'h3);
				// Trace: ../../rtl/VX_dispatch.sv:82:5
				wire [1:0] csr_op_type = sv2v_cast_2(VX_pipeline.issue.dispatch_if.op_type);
				// Trace: ../../rtl/VX_dispatch.sv:83:5
				wire [11:0] csr_addr = VX_pipeline.issue.dispatch_if.imm[11:0];
				// Trace: ../../rtl/VX_dispatch.sv:84:5
				wire [4:0] csr_imm = VX_pipeline.issue.dispatch_if.imm[12+:5];
				// Trace: ../../rtl/VX_dispatch.sv:85:5
				wire [31:0] csr_rs1_data = VX_pipeline.issue.gpr_rsp_if.rs1_data[tid * 32+:32];
				// Trace: ../../rtl/VX_dispatch.sv:87:5
				VX_skid_buffer #(
					.DATAW(137),
					.OUT_REG(1)
				) csr_buffer(
					.clk(clk),
					.reset(reset),
					.valid_in(csr_req_valid),
					.ready_in(csr_req_ready),
					.data_in({VX_pipeline.issue.dispatch_if.uuid, VX_pipeline.issue.dispatch_if.wid, VX_pipeline.issue.dispatch_if.tmask, VX_pipeline.issue.dispatch_if.PC, csr_op_type, csr_addr, VX_pipeline.issue.dispatch_if.rd, VX_pipeline.issue.dispatch_if.wb, VX_pipeline.issue.dispatch_if.use_imm, csr_imm, csr_rs1_data}),
					.data_out({VX_pipeline.csr_req_if.uuid, VX_pipeline.csr_req_if.wid, VX_pipeline.csr_req_if.tmask, VX_pipeline.csr_req_if.PC, VX_pipeline.csr_req_if.op_type, VX_pipeline.csr_req_if.addr, VX_pipeline.csr_req_if.rd, VX_pipeline.csr_req_if.wb, VX_pipeline.csr_req_if.use_imm, VX_pipeline.csr_req_if.imm, VX_pipeline.csr_req_if.rs1_data}),
					.valid_out(VX_pipeline.csr_req_if.valid),
					.ready_out(VX_pipeline.csr_req_if.ready)
				);
				// Trace: ../../rtl/VX_dispatch.sv:126:5
				wire gpu_req_valid = VX_pipeline.issue.dispatch_if.valid && (VX_pipeline.issue.dispatch_if.ex_type == 3'h5);
				// Trace: ../../rtl/VX_dispatch.sv:127:5
				wire [3:0] gpu_op_type = VX_pipeline.issue.dispatch_if.op_type;
				// Trace: ../../rtl/VX_dispatch.sv:129:5
				VX_skid_buffer #(
					.DATAW(317),
					.OUT_REG(1)
				) gpu_buffer(
					.clk(clk),
					.reset(reset),
					.valid_in(gpu_req_valid),
					.ready_in(gpu_req_ready),
					.data_in({VX_pipeline.issue.dispatch_if.uuid, VX_pipeline.issue.dispatch_if.wid, VX_pipeline.issue.dispatch_if.tmask, VX_pipeline.issue.dispatch_if.PC, next_PC, gpu_op_type, VX_pipeline.issue.dispatch_if.op_mod, VX_pipeline.issue.dispatch_if.rd, VX_pipeline.issue.dispatch_if.wb, tid, VX_pipeline.issue.gpr_rsp_if.rs1_data, VX_pipeline.issue.gpr_rsp_if.rs2_data, VX_pipeline.issue.gpr_rsp_if.rs3_data}),
					.data_out({VX_pipeline.gpu_req_if.uuid, VX_pipeline.gpu_req_if.wid, VX_pipeline.gpu_req_if.tmask, VX_pipeline.gpu_req_if.PC, VX_pipeline.gpu_req_if.next_PC, VX_pipeline.gpu_req_if.op_type, VX_pipeline.gpu_req_if.op_mod, VX_pipeline.gpu_req_if.rd, VX_pipeline.gpu_req_if.wb, VX_pipeline.gpu_req_if.tid, VX_pipeline.gpu_req_if.rs1_data, VX_pipeline.gpu_req_if.rs2_data, VX_pipeline.gpu_req_if.rs3_data}),
					.valid_out(VX_pipeline.gpu_req_if.valid),
					.ready_out(VX_pipeline.gpu_req_if.ready)
				);
				// Trace: ../../rtl/VX_dispatch.sv:144:5
				reg ready_r;
				// Trace: ../../rtl/VX_dispatch.sv:145:5
				always @(*)
					// Trace: ../../rtl/VX_dispatch.sv:146:9
					case (VX_pipeline.issue.dispatch_if.ex_type)
						3'h1:
							// Trace: ../../rtl/VX_dispatch.sv:147:18
							ready_r = alu_req_ready;
						3'h2:
							// Trace: ../../rtl/VX_dispatch.sv:148:18
							ready_r = lsu_req_ready;
						3'h3:
							// Trace: ../../rtl/VX_dispatch.sv:149:18
							ready_r = csr_req_ready;
						3'h5:
							// Trace: ../../rtl/VX_dispatch.sv:153:18
							ready_r = gpu_req_ready;
						default:
							// Trace: ../../rtl/VX_dispatch.sv:154:18
							ready_r = 1'b1;
					endcase
				// Trace: ../../rtl/VX_dispatch.sv:157:5
				assign VX_pipeline.issue.dispatch_if.ready = ready_r;
			end
			assign dispatch.clk = clk;
			assign dispatch.reset = dispatch_reset;
		end
	endgenerate
	assign issue.clk = clk;
	assign issue.reset = issue_reset;
	// Trace: ../../rtl/VX_pipeline.sv:201:5
	// expanded module instance: execute
	localparam _param_B78CA_CORE_ID = CORE_ID;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [25:0] sv2v_cast_26;
		input reg [25:0] inp;
		sv2v_cast_26 = inp;
	endfunction
	function automatic signed [25:0] sv2v_cast_26_signed;
		input reg signed [25:0] inp;
		sv2v_cast_26_signed = inp;
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	generate
		if (1) begin : execute
			// Trace: ../../rtl/VX_execute.sv:4:15
			localparam CORE_ID = _param_B78CA_CORE_ID;
			// Trace: ../../rtl/VX_execute.sv:8:5
			wire clk;
			// Trace: ../../rtl/VX_execute.sv:9:5
			wire reset;
			// Trace: ../../rtl/VX_execute.sv:12:5
			// removed modport instance dcache_req_if
			// Trace: ../../rtl/VX_execute.sv:13:5
			// removed modport instance dcache_rsp_if
			// Trace: ../../rtl/VX_execute.sv:16:5
			// removed modport instance cmt_to_csr_if
			// Trace: ../../rtl/VX_execute.sv:19:5
			// removed modport instance fetch_to_csr_if
			// Trace: ../../rtl/VX_execute.sv:27:5
			// removed modport instance alu_req_if
			// Trace: ../../rtl/VX_execute.sv:28:5
			// removed modport instance lsu_req_if
			// Trace: ../../rtl/VX_execute.sv:29:5
			// removed modport instance csr_req_if
			// Trace: ../../rtl/VX_execute.sv:33:5
			// removed modport instance gpu_req_if
			// Trace: ../../rtl/VX_execute.sv:36:5
			// removed modport instance branch_ctl_if
			// Trace: ../../rtl/VX_execute.sv:37:5
			// removed modport instance warp_ctl_if
			// Trace: ../../rtl/VX_execute.sv:38:5
			// removed modport instance alu_commit_if
			// Trace: ../../rtl/VX_execute.sv:39:5
			// removed modport instance ld_commit_if
			// Trace: ../../rtl/VX_execute.sv:40:5
			// removed modport instance st_commit_if
			// Trace: ../../rtl/VX_execute.sv:41:5
			// removed modport instance csr_commit_if
			// Trace: ../../rtl/VX_execute.sv:45:5
			// removed modport instance gpu_commit_if
			// Trace: ../../rtl/VX_execute.sv:47:5
			wire busy;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_execute.sv:133:22
			wire alu_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_execute.sv:133:55
			VX_reset_relay __alu_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(alu_reset)
			);
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_execute.sv:134:22
			wire lsu_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_execute.sv:134:55
			VX_reset_relay __lsu_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(lsu_reset)
			);
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_execute.sv:135:22
			wire csr_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_execute.sv:135:55
			VX_reset_relay __csr_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(csr_reset)
			);
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_execute.sv:136:22
			wire gpu_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/VX_execute.sv:136:55
			VX_reset_relay __gpu_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(gpu_reset)
			);
			// Trace: ../../rtl/VX_execute.sv:138:5
			// expanded module instance: alu_unit
			localparam _param_4B10A_CORE_ID = CORE_ID;
			if (1) begin : alu_unit
				// Trace: ../../rtl/VX_alu_unit.sv:4:15
				localparam CORE_ID = _param_4B10A_CORE_ID;
				// Trace: ../../rtl/VX_alu_unit.sv:6:5
				wire clk;
				// Trace: ../../rtl/VX_alu_unit.sv:7:5
				wire reset;
				// Trace: ../../rtl/VX_alu_unit.sv:10:5
				// removed modport instance alu_req_if
				// Trace: ../../rtl/VX_alu_unit.sv:13:5
				// removed modport instance branch_ctl_if
				// Trace: ../../rtl/VX_alu_unit.sv:14:5
				// removed modport instance alu_commit_if
				// Trace: ../../rtl/VX_alu_unit.sv:19:5
				reg [63:0] alu_result;
				// Trace: ../../rtl/VX_alu_unit.sv:20:5
				wire [63:0] add_result;
				// Trace: ../../rtl/VX_alu_unit.sv:21:5
				wire [65:0] sub_result;
				// Trace: ../../rtl/VX_alu_unit.sv:22:5
				wire [63:0] shr_result;
				// Trace: ../../rtl/VX_alu_unit.sv:23:5
				reg [63:0] msc_result;
				// Trace: ../../rtl/VX_alu_unit.sv:25:5
				wire ready_in;
				// Trace: ../../rtl/VX_alu_unit.sv:28:5
				wire is_br_op = VX_pipeline.alu_req_if.op_mod[0];
				// Trace: ../../rtl/VX_alu_unit.sv:29:5
				wire [3:0] alu_op = VX_pipeline.alu_req_if.op_type;
				// Trace: ../../rtl/VX_alu_unit.sv:30:5
				wire [3:0] br_op = VX_pipeline.alu_req_if.op_type;
				// Trace: ../../rtl/VX_alu_unit.sv:31:5
				wire alu_signed = alu_op[0];
				// Trace: ../../rtl/VX_alu_unit.sv:32:5
				wire [1:0] alu_op_class = alu_op[3:2];
				// Trace: ../../rtl/VX_alu_unit.sv:33:5
				wire is_sub = alu_op == 4'b1011;
				// Trace: ../../rtl/VX_alu_unit.sv:35:5
				wire [63:0] alu_in1 = VX_pipeline.alu_req_if.rs1_data;
				// Trace: ../../rtl/VX_alu_unit.sv:36:5
				wire [63:0] alu_in2 = VX_pipeline.alu_req_if.rs2_data;
				// Trace: ../../rtl/VX_alu_unit.sv:38:5
				wire [63:0] alu_in1_PC = (VX_pipeline.alu_req_if.use_PC ? {2 {VX_pipeline.alu_req_if.PC}} : alu_in1);
				// Trace: ../../rtl/VX_alu_unit.sv:39:5
				wire [63:0] alu_in2_imm = (VX_pipeline.alu_req_if.use_imm ? {2 {VX_pipeline.alu_req_if.imm}} : alu_in2);
				// Trace: ../../rtl/VX_alu_unit.sv:40:5
				wire [63:0] alu_in2_less = (VX_pipeline.alu_req_if.use_imm && ~is_br_op ? {2 {VX_pipeline.alu_req_if.imm}} : alu_in2);
				// Trace: ../../rtl/VX_alu_unit.sv:42:5
				genvar i;
				for (i = 0; i < 2; i = i + 1) begin : genblk1
					// Trace: ../../rtl/VX_alu_unit.sv:43:9
					assign add_result[i * 32+:32] = alu_in1_PC[i * 32+:32] + alu_in2_imm[i * 32+:32];
				end
				// Trace: ../../rtl/VX_alu_unit.sv:46:5
				for (i = 0; i < 2; i = i + 1) begin : genblk2
					// Trace: ../../rtl/VX_alu_unit.sv:47:9
					wire [32:0] sub_in1 = {alu_signed & alu_in1[(i * 32) + 31], alu_in1[i * 32+:32]};
					// Trace: ../../rtl/VX_alu_unit.sv:48:9
					wire [32:0] sub_in2 = {alu_signed & alu_in2_less[(i * 32) + 31], alu_in2_less[i * 32+:32]};
					// Trace: ../../rtl/VX_alu_unit.sv:49:9
					assign sub_result[i * 33+:33] = sub_in1 - sub_in2;
				end
				// Trace: ../../rtl/VX_alu_unit.sv:52:5
				for (i = 0; i < 2; i = i + 1) begin : genblk3
					// Trace: ../../rtl/VX_alu_unit.sv:53:9
					wire [32:0] shr_in1 = {alu_signed & alu_in1[(i * 32) + 31], alu_in1[i * 32+:32]};
					// Trace: ../../rtl/VX_alu_unit.sv:54:9
					assign shr_result[i * 32+:32] = sv2v_cast_32_signed($signed(shr_in1) >>> alu_in2_imm[(i * 32) + 4-:5]);
				end
				// Trace: ../../rtl/VX_alu_unit.sv:57:5
				for (i = 0; i < 2; i = i + 1) begin : genblk4
					// Trace: ../../rtl/VX_alu_unit.sv:58:9
					always @(*)
						// Trace: ../../rtl/VX_alu_unit.sv:59:13
						case (alu_op)
							4'b1100:
								// Trace: ../../rtl/VX_alu_unit.sv:60:32
								msc_result[i * 32+:32] = alu_in1[i * 32+:32] & alu_in2_imm[i * 32+:32];
							4'b1101:
								// Trace: ../../rtl/VX_alu_unit.sv:61:32
								msc_result[i * 32+:32] = alu_in1[i * 32+:32] | alu_in2_imm[i * 32+:32];
							4'b1110:
								// Trace: ../../rtl/VX_alu_unit.sv:62:32
								msc_result[i * 32+:32] = alu_in1[i * 32+:32] ^ alu_in2_imm[i * 32+:32];
							default:
								// Trace: ../../rtl/VX_alu_unit.sv:64:27
								msc_result[i * 32+:32] = alu_in1[i * 32+:32] << alu_in2_imm[(i * 32) + 4-:5];
						endcase
				end
				// Trace: ../../rtl/VX_alu_unit.sv:69:5
				for (i = 0; i < 2; i = i + 1) begin : genblk5
					// Trace: ../../rtl/VX_alu_unit.sv:70:9
					always @(*)
						// Trace: ../../rtl/VX_alu_unit.sv:71:13
						case (alu_op_class)
							2'b00:
								// Trace: ../../rtl/VX_alu_unit.sv:72:24
								alu_result[i * 32+:32] = add_result[i * 32+:32];
							2'b01:
								// Trace: ../../rtl/VX_alu_unit.sv:73:24
								alu_result[i * 32+:32] = {31'b0000000000000000000000000000000, sub_result[(i * 33) + 32]};
							2'b10:
								// Trace: ../../rtl/VX_alu_unit.sv:74:24
								alu_result[i * 32+:32] = (is_sub ? sub_result[(i * 33) + 31-:32] : shr_result[i * 32+:32]);
							default:
								// Trace: ../../rtl/VX_alu_unit.sv:77:26
								alu_result[i * 32+:32] = msc_result[i * 32+:32];
						endcase
				end
				// Trace: ../../rtl/VX_alu_unit.sv:84:5
				wire is_jal = is_br_op && ((br_op == 4'b1000) || (br_op == 4'b1001));
				// Trace: ../../rtl/VX_alu_unit.sv:85:5
				wire [63:0] alu_jal_result = (is_jal ? {2 {VX_pipeline.alu_req_if.next_PC}} : alu_result);
				// Trace: ../../rtl/VX_alu_unit.sv:87:5
				wire [31:0] br_dest = add_result[VX_pipeline.alu_req_if.tid * 32+:32];
				// Trace: ../../rtl/VX_alu_unit.sv:88:5
				wire [32:0] cmp_result = sub_result[VX_pipeline.alu_req_if.tid * 33+:33];
				// Trace: ../../rtl/VX_alu_unit.sv:90:5
				wire is_less = cmp_result[32];
				// Trace: ../../rtl/VX_alu_unit.sv:91:5
				wire is_equal = ~(|cmp_result[31:0]);
				// Trace: ../../rtl/VX_alu_unit.sv:95:5
				wire alu_valid_in;
				// Trace: ../../rtl/VX_alu_unit.sv:96:5
				wire alu_ready_in;
				// Trace: ../../rtl/VX_alu_unit.sv:97:5
				wire alu_valid_out;
				// Trace: ../../rtl/VX_alu_unit.sv:98:5
				wire alu_ready_out;
				// Trace: ../../rtl/VX_alu_unit.sv:99:5
				wire [43:0] alu_uuid;
				// Trace: ../../rtl/VX_alu_unit.sv:100:5
				wire [0:0] alu_wid;
				// Trace: ../../rtl/VX_alu_unit.sv:101:5
				wire [1:0] alu_tmask;
				// Trace: ../../rtl/VX_alu_unit.sv:102:5
				wire [31:0] alu_PC;
				// Trace: ../../rtl/VX_alu_unit.sv:103:5
				wire [4:0] alu_rd;
				// Trace: ../../rtl/VX_alu_unit.sv:104:5
				wire alu_wb;
				// Trace: ../../rtl/VX_alu_unit.sv:105:5
				wire [63:0] alu_data;
				// Trace: ../../rtl/VX_alu_unit.sv:107:5
				wire [3:0] br_op_r;
				// Trace: ../../rtl/VX_alu_unit.sv:108:5
				wire [31:0] br_dest_r;
				// Trace: ../../rtl/VX_alu_unit.sv:109:5
				wire is_less_r;
				// Trace: ../../rtl/VX_alu_unit.sv:110:5
				wire is_equal_r;
				// Trace: ../../rtl/VX_alu_unit.sv:111:5
				wire is_br_op_r;
				// Trace: ../../rtl/VX_alu_unit.sv:113:5
				assign alu_ready_in = alu_ready_out || ~alu_valid_out;
				// Trace: ../../rtl/VX_alu_unit.sv:115:5
				VX_pipe_register #(
					.DATAW(189),
					.RESETW(1)
				) pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(alu_ready_in),
					.data_in({alu_valid_in, VX_pipeline.alu_req_if.uuid, VX_pipeline.alu_req_if.wid, VX_pipeline.alu_req_if.tmask, VX_pipeline.alu_req_if.PC, VX_pipeline.alu_req_if.rd, VX_pipeline.alu_req_if.wb, alu_jal_result, is_br_op, br_op, is_less, is_equal, br_dest}),
					.data_out({alu_valid_out, alu_uuid, alu_wid, alu_tmask, alu_PC, alu_rd, alu_wb, alu_data, is_br_op_r, br_op_r, is_less_r, is_equal_r, br_dest_r})
				);
				// Trace: ../../rtl/VX_alu_unit.sv:127:5
				wire br_neg = br_op_r[1];
				// Trace: ../../rtl/VX_alu_unit.sv:128:5
				wire br_less = br_op_r[2];
				// Trace: ../../rtl/VX_alu_unit.sv:129:5
				wire br_static = br_op_r[3];
				// Trace: ../../rtl/VX_alu_unit.sv:131:5
				assign VX_pipeline.branch_ctl_if.valid = (alu_valid_out && alu_ready_out) && is_br_op_r;
				// Trace: ../../rtl/VX_alu_unit.sv:132:5
				assign VX_pipeline.branch_ctl_if.taken = ((br_less ? is_less_r : is_equal_r) ^ br_neg) | br_static;
				// Trace: ../../rtl/VX_alu_unit.sv:133:5
				assign VX_pipeline.branch_ctl_if.wid = alu_wid;
				// Trace: ../../rtl/VX_alu_unit.sv:134:5
				assign VX_pipeline.branch_ctl_if.dest = br_dest_r;
				// Trace: ../../rtl/VX_alu_unit.sv:138:5
				wire mul_valid_in;
				// Trace: ../../rtl/VX_alu_unit.sv:139:5
				wire mul_ready_in;
				// Trace: ../../rtl/VX_alu_unit.sv:140:5
				wire mul_valid_out;
				// Trace: ../../rtl/VX_alu_unit.sv:141:5
				wire mul_ready_out;
				// Trace: ../../rtl/VX_alu_unit.sv:142:5
				wire [43:0] mul_uuid;
				// Trace: ../../rtl/VX_alu_unit.sv:143:5
				wire [0:0] mul_wid;
				// Trace: ../../rtl/VX_alu_unit.sv:144:5
				wire [1:0] mul_tmask;
				// Trace: ../../rtl/VX_alu_unit.sv:145:5
				wire [31:0] mul_PC;
				// Trace: ../../rtl/VX_alu_unit.sv:146:5
				wire [4:0] mul_rd;
				// Trace: ../../rtl/VX_alu_unit.sv:147:5
				wire mul_wb;
				// Trace: ../../rtl/VX_alu_unit.sv:148:5
				wire [63:0] mul_data;
				// Trace: ../../rtl/VX_alu_unit.sv:150:5
				wire [2:0] mul_op = sv2v_cast_3(VX_pipeline.alu_req_if.op_type);
				// Trace: ../../rtl/VX_alu_unit.sv:152:5
				VX_muldiv muldiv(
					.clk(clk),
					.reset(reset),
					.alu_op(mul_op),
					.uuid_in(VX_pipeline.alu_req_if.uuid),
					.wid_in(VX_pipeline.alu_req_if.wid),
					.tmask_in(VX_pipeline.alu_req_if.tmask),
					.PC_in(VX_pipeline.alu_req_if.PC),
					.rd_in(VX_pipeline.alu_req_if.rd),
					.wb_in(VX_pipeline.alu_req_if.wb),
					.alu_in1(VX_pipeline.alu_req_if.rs1_data),
					.alu_in2(VX_pipeline.alu_req_if.rs2_data),
					.wid_out(mul_wid),
					.uuid_out(mul_uuid),
					.tmask_out(mul_tmask),
					.PC_out(mul_PC),
					.rd_out(mul_rd),
					.wb_out(mul_wb),
					.data_out(mul_data),
					.valid_in(mul_valid_in),
					.ready_in(mul_ready_in),
					.valid_out(mul_valid_out),
					.ready_out(mul_ready_out)
				);
				// Trace: ../../rtl/VX_alu_unit.sv:183:5
				wire is_mul_op = VX_pipeline.alu_req_if.op_mod[1];
				// Trace: ../../rtl/VX_alu_unit.sv:185:5
				assign ready_in = (is_mul_op ? mul_ready_in : alu_ready_in);
				// Trace: ../../rtl/VX_alu_unit.sv:187:5
				assign alu_valid_in = VX_pipeline.alu_req_if.valid && ~is_mul_op;
				// Trace: ../../rtl/VX_alu_unit.sv:188:5
				assign mul_valid_in = VX_pipeline.alu_req_if.valid && is_mul_op;
				// Trace: ../../rtl/VX_alu_unit.sv:190:5
				assign VX_pipeline.alu_commit_if.valid = alu_valid_out || mul_valid_out;
				// Trace: ../../rtl/VX_alu_unit.sv:191:5
				assign VX_pipeline.alu_commit_if.uuid = (alu_valid_out ? alu_uuid : mul_uuid);
				// Trace: ../../rtl/VX_alu_unit.sv:192:5
				assign VX_pipeline.alu_commit_if.wid = (alu_valid_out ? alu_wid : mul_wid);
				// Trace: ../../rtl/VX_alu_unit.sv:193:5
				assign VX_pipeline.alu_commit_if.tmask = (alu_valid_out ? alu_tmask : mul_tmask);
				// Trace: ../../rtl/VX_alu_unit.sv:194:5
				assign VX_pipeline.alu_commit_if.PC = (alu_valid_out ? alu_PC : mul_PC);
				// Trace: ../../rtl/VX_alu_unit.sv:195:5
				assign VX_pipeline.alu_commit_if.rd = (alu_valid_out ? alu_rd : mul_rd);
				// Trace: ../../rtl/VX_alu_unit.sv:196:5
				assign VX_pipeline.alu_commit_if.wb = (alu_valid_out ? alu_wb : mul_wb);
				// Trace: ../../rtl/VX_alu_unit.sv:197:5
				assign VX_pipeline.alu_commit_if.data = (alu_valid_out ? alu_data : mul_data);
				// Trace: ../../rtl/VX_alu_unit.sv:199:5
				assign alu_ready_out = VX_pipeline.alu_commit_if.ready;
				// Trace: ../../rtl/VX_alu_unit.sv:200:5
				assign mul_ready_out = VX_pipeline.alu_commit_if.ready & ~alu_valid_out;
				// Trace: ../../rtl/VX_alu_unit.sv:221:5
				assign VX_pipeline.alu_commit_if.eop = 1'b1;
				// Trace: ../../rtl/VX_alu_unit.sv:224:5
				assign VX_pipeline.alu_req_if.ready = ready_in;
			end
			assign alu_unit.clk = clk;
			assign alu_unit.reset = alu_reset;
			// Trace: ../../rtl/VX_execute.sv:148:5
			// expanded module instance: lsu_unit
			localparam _param_54826_CORE_ID = CORE_ID;
			if (1) begin : lsu_unit
				// Trace: ../../rtl/VX_lsu_unit.sv:4:15
				localparam CORE_ID = _param_54826_CORE_ID;
				// Trace: ../../rtl/VX_lsu_unit.sv:8:5
				wire clk;
				// Trace: ../../rtl/VX_lsu_unit.sv:9:5
				wire reset;
				// Trace: ../../rtl/VX_lsu_unit.sv:12:5
				// removed modport instance dcache_req_if
				// Trace: ../../rtl/VX_lsu_unit.sv:13:5
				// removed modport instance dcache_rsp_if
				// Trace: ../../rtl/VX_lsu_unit.sv:16:5
				// removed modport instance lsu_req_if
				// Trace: ../../rtl/VX_lsu_unit.sv:19:5
				// removed modport instance ld_commit_if
				// Trace: ../../rtl/VX_lsu_unit.sv:20:5
				// removed modport instance st_commit_if
				// Trace: ../../rtl/VX_lsu_unit.sv:22:5
				localparam MEM_ASHIFT = 6;
				// Trace: ../../rtl/VX_lsu_unit.sv:23:5
				localparam MEM_ADDRW = 26;
				// Trace: ../../rtl/VX_lsu_unit.sv:24:5
				localparam REQ_ASHIFT = 2;
				// Trace: ../../rtl/VX_lsu_unit.sv:30:5
				wire req_valid;
				// Trace: ../../rtl/VX_lsu_unit.sv:31:5
				wire [43:0] req_uuid;
				// Trace: ../../rtl/VX_lsu_unit.sv:32:5
				wire [1:0] req_tmask;
				// Trace: ../../rtl/VX_lsu_unit.sv:33:5
				wire [63:0] req_addr;
				// Trace: ../../rtl/VX_lsu_unit.sv:34:5
				wire [3:0] req_type;
				// Trace: ../../rtl/VX_lsu_unit.sv:35:5
				wire [63:0] req_data;
				// Trace: ../../rtl/VX_lsu_unit.sv:36:5
				wire [4:0] req_rd;
				// Trace: ../../rtl/VX_lsu_unit.sv:37:5
				wire req_wb;
				// Trace: ../../rtl/VX_lsu_unit.sv:38:5
				wire [0:0] req_wid;
				// Trace: ../../rtl/VX_lsu_unit.sv:39:5
				wire [31:0] req_pc;
				// Trace: ../../rtl/VX_lsu_unit.sv:40:5
				wire req_is_dup;
				// Trace: ../../rtl/VX_lsu_unit.sv:41:5
				wire req_is_prefetch;
				// Trace: ../../rtl/VX_lsu_unit.sv:43:5
				wire mbuf_empty;
				// Trace: ../../rtl/VX_lsu_unit.sv:45:5
				wire [3:0] lsu_addr_type;
				wire [3:0] req_addr_type;
				// Trace: ../../rtl/VX_lsu_unit.sv:48:5
				wire [63:0] full_addr;
				// Trace: ../../rtl/VX_lsu_unit.sv:49:5
				genvar i;
				for (i = 0; i < 2; i = i + 1) begin : genblk1
					// Trace: ../../rtl/VX_lsu_unit.sv:50:9
					assign full_addr[i * 32+:32] = VX_pipeline.lsu_req_if.base_addr[i * 32+:32] + VX_pipeline.lsu_req_if.offset;
				end
				// Trace: ../../rtl/VX_lsu_unit.sv:54:5
				wire [0:0] addr_matches;
				// Trace: ../../rtl/VX_lsu_unit.sv:55:5
				for (i = 0; i < 1; i = i + 1) begin : genblk2
					// Trace: ../../rtl/VX_lsu_unit.sv:56:9
					assign addr_matches[i] = (VX_pipeline.lsu_req_if.base_addr[(i + 1) * 32+:32] == VX_pipeline.lsu_req_if.base_addr[0+:32]) || ~VX_pipeline.lsu_req_if.tmask[i + 1];
				end
				// Trace: ../../rtl/VX_lsu_unit.sv:59:5
				wire lsu_is_dup = VX_pipeline.lsu_req_if.tmask[0] && &addr_matches;
				// Trace: ../../rtl/VX_lsu_unit.sv:61:5
				for (i = 0; i < 2; i = i + 1) begin : genblk3
					// Trace: ../../rtl/VX_lsu_unit.sv:63:9
					wire is_addr_nc = full_addr[(i * 32) + MEM_ASHIFT+:MEM_ADDRW] >= sv2v_cast_26(32'hff000000 >> MEM_ASHIFT);
					if (1) begin : genblk1
						// Trace: ../../rtl/VX_lsu_unit.sv:66:13
						wire is_addr_sm = (full_addr[(i * 32) + MEM_ASHIFT+:MEM_ADDRW] >= sv2v_cast_26_signed(33'sd4278185984 >> MEM_ASHIFT)) & (full_addr[(i * 32) + MEM_ASHIFT+:MEM_ADDRW] < sv2v_cast_26(32'hff000000 >> MEM_ASHIFT));
						// Trace: ../../rtl/VX_lsu_unit.sv:68:13
						assign lsu_addr_type[i * 2+:2] = {is_addr_nc, is_addr_sm};
					end
				end
				// Trace: ../../rtl/VX_lsu_unit.sv:75:5
				wire fence_wait = VX_pipeline.lsu_req_if.is_fence && (req_valid || !mbuf_empty);
				// Trace: ../../rtl/VX_lsu_unit.sv:77:5
				wire ready_in;
				// Trace: ../../rtl/VX_lsu_unit.sv:78:5
				wire stall_in = ~ready_in && req_valid;
				// Trace: ../../rtl/VX_lsu_unit.sv:80:5
				wire lsu_valid = VX_pipeline.lsu_req_if.valid && ~fence_wait;
				// Trace: ../../rtl/VX_lsu_unit.sv:82:5
				wire lsu_wb = VX_pipeline.lsu_req_if.wb | VX_pipeline.lsu_req_if.is_prefetch;
				// Trace: ../../rtl/VX_lsu_unit.sv:84:5
				VX_pipe_register #(
					.DATAW(224),
					.RESETW(1)
				) req_pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(!stall_in),
					.data_in({lsu_valid, lsu_is_dup, VX_pipeline.lsu_req_if.is_prefetch, VX_pipeline.lsu_req_if.uuid, VX_pipeline.lsu_req_if.wid, VX_pipeline.lsu_req_if.tmask, VX_pipeline.lsu_req_if.PC, full_addr, lsu_addr_type, VX_pipeline.lsu_req_if.op_type, VX_pipeline.lsu_req_if.rd, lsu_wb, VX_pipeline.lsu_req_if.store_data}),
					.data_out({req_valid, req_is_dup, req_is_prefetch, req_uuid, req_wid, req_tmask, req_pc, req_addr, req_addr_type, req_type, req_rd, req_wb, req_data})
				);
				// Trace: ../../rtl/VX_lsu_unit.sv:96:5
				assign VX_pipeline.lsu_req_if.ready = ~stall_in && ~fence_wait;
				// Trace: ../../rtl/VX_lsu_unit.sv:98:5
				wire [43:0] rsp_uuid;
				// Trace: ../../rtl/VX_lsu_unit.sv:99:5
				wire [0:0] rsp_wid;
				// Trace: ../../rtl/VX_lsu_unit.sv:100:5
				wire [31:0] rsp_pc;
				// Trace: ../../rtl/VX_lsu_unit.sv:101:5
				wire [4:0] rsp_rd;
				// Trace: ../../rtl/VX_lsu_unit.sv:102:5
				wire rsp_wb;
				// Trace: ../../rtl/VX_lsu_unit.sv:103:5
				wire [3:0] rsp_type;
				// Trace: ../../rtl/VX_lsu_unit.sv:104:5
				wire rsp_is_dup;
				// Trace: ../../rtl/VX_lsu_unit.sv:105:5
				wire rsp_is_prefetch;
				// Trace: ../../rtl/VX_lsu_unit.sv:107:5
				reg [7:0] rsp_rem_mask;
				// Trace: ../../rtl/VX_lsu_unit.sv:108:5
				wire [1:0] rsp_rem_mask_n;
				// Trace: ../../rtl/VX_lsu_unit.sv:109:5
				wire [1:0] rsp_tmask;
				// Trace: ../../rtl/VX_lsu_unit.sv:111:5
				reg [1:0] req_sent_mask;
				// Trace: ../../rtl/VX_lsu_unit.sv:112:5
				reg is_req_start;
				// Trace: ../../rtl/VX_lsu_unit.sv:114:5
				wire [1:0] mbuf_waddr;
				wire [1:0] mbuf_raddr;
				// Trace: ../../rtl/VX_lsu_unit.sv:115:5
				wire mbuf_full;
				// Trace: ../../rtl/VX_lsu_unit.sv:120:5
				wire [3:0] req_offset;
				wire [3:0] rsp_offset;
				// Trace: ../../rtl/VX_lsu_unit.sv:121:5
				for (i = 0; i < 2; i = i + 1) begin : genblk4
					// Trace: ../../rtl/VX_lsu_unit.sv:122:9
					assign req_offset[i * 2+:2] = req_addr[(i * 32) + 1-:2];
				end
				// Trace: ../../rtl/VX_lsu_unit.sv:125:5
				wire [1:0] dcache_req_fire = VX_pipeline.dcache_req_if.valid & VX_pipeline.dcache_req_if.ready;
				// Trace: ../../rtl/VX_lsu_unit.sv:127:5
				wire dcache_rsp_fire = VX_pipeline.dcache_rsp_if.valid && VX_pipeline.dcache_rsp_if.ready;
				// Trace: ../../rtl/VX_lsu_unit.sv:129:5
				wire [1:0] req_tmask_dup = req_tmask & {~req_is_dup, 1'b1};
				// Trace: ../../rtl/VX_lsu_unit.sv:131:5
				wire mbuf_push = ((~mbuf_full && |(({2 {req_valid}} & req_tmask_dup) & VX_pipeline.dcache_req_if.ready)) && is_req_start) && req_wb;
				// Trace: ../../rtl/VX_lsu_unit.sv:136:5
				wire mbuf_pop = dcache_rsp_fire && (0 == rsp_rem_mask_n);
				// Trace: ../../rtl/VX_lsu_unit.sv:138:5
				assign mbuf_raddr = VX_pipeline.dcache_rsp_if.tag[2+:2];
				// Trace: ../../rtl/VX_lsu_unit.sv:142:5
				wire req_wb2 = req_wb && ~req_is_prefetch;
				// Trace: ../../rtl/VX_lsu_unit.sv:144:5
				VX_index_buffer #(
					.DATAW(95),
					.SIZE(4)
				) req_metadata(
					.clk(clk),
					.reset(reset),
					.write_addr(mbuf_waddr),
					.acquire_slot(mbuf_push),
					.read_addr(mbuf_raddr),
					.write_data({req_uuid, req_wid, req_pc, req_tmask, req_rd, req_wb2, req_type, req_offset, req_is_dup, req_is_prefetch}),
					.read_data({rsp_uuid, rsp_wid, rsp_pc, rsp_tmask, rsp_rd, rsp_wb, rsp_type, rsp_offset, rsp_is_dup, rsp_is_prefetch}),
					.release_addr(mbuf_raddr),
					.release_slot(mbuf_pop),
					.full(mbuf_full),
					.empty(mbuf_empty)
				);
				// Trace: ../../rtl/VX_lsu_unit.sv:161:5
				wire dcache_req_ready = &((VX_pipeline.dcache_req_if.ready | req_sent_mask) | ~req_tmask_dup);
				// Trace: ../../rtl/VX_lsu_unit.sv:163:5
				wire [1:0] req_sent_mask_n = req_sent_mask | dcache_req_fire;
				// Trace: ../../rtl/VX_lsu_unit.sv:165:5
				always @(posedge clk)
					// Trace: ../../rtl/VX_lsu_unit.sv:166:9
					if (reset) begin
						// Trace: ../../rtl/VX_lsu_unit.sv:167:13
						req_sent_mask <= 0;
						// Trace: ../../rtl/VX_lsu_unit.sv:168:13
						is_req_start <= 1;
					end
					else
						// Trace: ../../rtl/VX_lsu_unit.sv:170:13
						if (dcache_req_ready) begin
							// Trace: ../../rtl/VX_lsu_unit.sv:171:17
							req_sent_mask <= 0;
							// Trace: ../../rtl/VX_lsu_unit.sv:172:17
							is_req_start <= 1;
						end
						else begin
							// Trace: ../../rtl/VX_lsu_unit.sv:174:17
							req_sent_mask <= req_sent_mask_n;
							// Trace: ../../rtl/VX_lsu_unit.sv:175:17
							is_req_start <= 0 == req_sent_mask_n;
						end
				// Trace: ../../rtl/VX_lsu_unit.sv:181:5
				reg [1:0] req_tag_hold;
				// Trace: ../../rtl/VX_lsu_unit.sv:182:5
				wire [1:0] req_tag = (is_req_start ? mbuf_waddr : req_tag_hold);
				// Trace: ../../rtl/VX_lsu_unit.sv:183:5
				always @(posedge clk)
					// Trace: ../../rtl/VX_lsu_unit.sv:184:9
					if (mbuf_push)
						// Trace: ../../rtl/VX_lsu_unit.sv:185:13
						req_tag_hold <= mbuf_waddr;
				// Trace: ../../rtl/VX_lsu_unit.sv:189:5
				assign rsp_rem_mask_n = rsp_rem_mask[mbuf_raddr * 2+:2] & ~VX_pipeline.dcache_rsp_if.tmask;
				// Trace: ../../rtl/VX_lsu_unit.sv:191:5
				always @(posedge clk) begin
					// Trace: ../../rtl/VX_lsu_unit.sv:192:9
					if (mbuf_push)
						// Trace: ../../rtl/VX_lsu_unit.sv:193:13
						rsp_rem_mask[mbuf_waddr * 2+:2] <= req_tmask_dup;
					if (dcache_rsp_fire)
						// Trace: ../../rtl/VX_lsu_unit.sv:196:13
						rsp_rem_mask[mbuf_raddr * 2+:2] <= rsp_rem_mask_n;
				end
				// Trace: ../../rtl/VX_lsu_unit.sv:201:5
				wire req_dep_ready = (req_wb && ~(mbuf_full && is_req_start)) || (~req_wb && VX_pipeline.st_commit_if.ready);
				// Trace: ../../rtl/VX_lsu_unit.sv:206:5
				for (i = 0; i < 2; i = i + 1) begin : genblk5
					// Trace: ../../rtl/VX_lsu_unit.sv:208:9
					reg [3:0] mem_req_byteen;
					// Trace: ../../rtl/VX_lsu_unit.sv:209:9
					reg [31:0] mem_req_data;
					// Trace: ../../rtl/VX_lsu_unit.sv:211:9
					always @(*) begin
						// Trace: ../../rtl/VX_lsu_unit.sv:212:13
						mem_req_byteen = {4 {req_wb}};
						// Trace: ../../rtl/VX_lsu_unit.sv:213:13
						case (req_type[1:0])
							0:
								// Trace: ../../rtl/VX_lsu_unit.sv:214:20
								mem_req_byteen[req_offset[i * 2+:2]] = 1;
							1: begin
								// Trace: ../../rtl/VX_lsu_unit.sv:216:21
								mem_req_byteen[req_offset[i * 2+:2]] = 1;
								// Trace: ../../rtl/VX_lsu_unit.sv:217:21
								mem_req_byteen[{req_offset[(i * 2) + 1], 1'b1}] = 1;
							end
							default:
								// Trace: ../../rtl/VX_lsu_unit.sv:219:27
								mem_req_byteen = {4 {1'b1}};
						endcase
					end
					// Trace: ../../rtl/VX_lsu_unit.sv:223:9
					always @(*) begin
						// Trace: ../../rtl/VX_lsu_unit.sv:224:13
						mem_req_data = req_data[i * 32+:32];
						// Trace: ../../rtl/VX_lsu_unit.sv:225:13
						case (req_offset[i * 2+:2])
							1:
								// Trace: ../../rtl/VX_lsu_unit.sv:226:20
								mem_req_data[31:8] = req_data[(i * 32) + 23-:24];
							2:
								// Trace: ../../rtl/VX_lsu_unit.sv:227:20
								mem_req_data[31:16] = req_data[(i * 32) + 15-:16];
							3:
								// Trace: ../../rtl/VX_lsu_unit.sv:228:20
								mem_req_data[31:24] = req_data[(i * 32) + 7-:8];
							default:
								;
						endcase
					end
					// Trace: ../../rtl/VX_lsu_unit.sv:233:9
					assign VX_pipeline.dcache_req_if.valid[i] = ((req_valid && req_dep_ready) && req_tmask_dup[i]) && !req_sent_mask[i];
					// Trace: ../../rtl/VX_lsu_unit.sv:234:9
					assign VX_pipeline.dcache_req_if.rw[i] = ~req_wb;
					// Trace: ../../rtl/VX_lsu_unit.sv:235:9
					assign VX_pipeline.dcache_req_if.addr[i * 30+:30] = req_addr[(i * 32) + 31-:30];
					// Trace: ../../rtl/VX_lsu_unit.sv:236:9
					assign VX_pipeline.dcache_req_if.byteen[i * 4+:4] = mem_req_byteen;
					// Trace: ../../rtl/VX_lsu_unit.sv:237:9
					assign VX_pipeline.dcache_req_if.data[i * 32+:32] = mem_req_data;
					// Trace: ../../rtl/VX_lsu_unit.sv:238:9
					assign VX_pipeline.dcache_req_if.tag[i * 48+:48] = {req_uuid, req_tag, req_addr_type[i * 2+:2]};
				end
				// Trace: ../../rtl/VX_lsu_unit.sv:241:5
				assign ready_in = req_dep_ready && dcache_req_ready;
				// Trace: ../../rtl/VX_lsu_unit.sv:245:5
				wire is_store_rsp = (req_valid && ~req_wb) && dcache_req_ready;
				// Trace: ../../rtl/VX_lsu_unit.sv:247:5
				assign VX_pipeline.st_commit_if.valid = is_store_rsp;
				// Trace: ../../rtl/VX_lsu_unit.sv:248:5
				assign VX_pipeline.st_commit_if.uuid = req_uuid;
				// Trace: ../../rtl/VX_lsu_unit.sv:249:5
				assign VX_pipeline.st_commit_if.wid = req_wid;
				// Trace: ../../rtl/VX_lsu_unit.sv:250:5
				assign VX_pipeline.st_commit_if.tmask = req_tmask;
				// Trace: ../../rtl/VX_lsu_unit.sv:251:5
				assign VX_pipeline.st_commit_if.PC = req_pc;
				// Trace: ../../rtl/VX_lsu_unit.sv:252:5
				assign VX_pipeline.st_commit_if.rd = 0;
				// Trace: ../../rtl/VX_lsu_unit.sv:253:5
				assign VX_pipeline.st_commit_if.wb = 0;
				// Trace: ../../rtl/VX_lsu_unit.sv:254:5
				assign VX_pipeline.st_commit_if.eop = 1'b1;
				// Trace: ../../rtl/VX_lsu_unit.sv:255:5
				assign VX_pipeline.st_commit_if.data = 0;
				// Trace: ../../rtl/VX_lsu_unit.sv:259:5
				reg [63:0] rsp_data;
				// Trace: ../../rtl/VX_lsu_unit.sv:260:5
				wire [1:0] rsp_tmask_qual;
				// Trace: ../../rtl/VX_lsu_unit.sv:262:5
				for (i = 0; i < 2; i = i + 1) begin : genblk6
					// Trace: ../../rtl/VX_lsu_unit.sv:263:9
					wire [31:0] rsp_data32 = ((i == 0) || rsp_is_dup ? VX_pipeline.dcache_rsp_if.data[0+:32] : VX_pipeline.dcache_rsp_if.data[i * 32+:32]);
					// Trace: ../../rtl/VX_lsu_unit.sv:264:9
					wire [15:0] rsp_data16 = (rsp_offset[(i * 2) + 1] ? rsp_data32[31:16] : rsp_data32[15:0]);
					// Trace: ../../rtl/VX_lsu_unit.sv:265:9
					wire [7:0] rsp_data8 = (rsp_offset[i * 2] ? rsp_data16[15:8] : rsp_data16[7:0]);
					// Trace: ../../rtl/VX_lsu_unit.sv:267:9
					always @(*)
						// Trace: ../../rtl/VX_lsu_unit.sv:268:13
						case (rsp_type[2:0])
							3'b000:
								// Trace: ../../rtl/VX_lsu_unit.sv:269:27
								rsp_data[i * 32+:32] = sv2v_cast_32_signed($signed(rsp_data8));
							3'b001:
								// Trace: ../../rtl/VX_lsu_unit.sv:270:27
								rsp_data[i * 32+:32] = sv2v_cast_32_signed($signed(rsp_data16));
							3'b100:
								// Trace: ../../rtl/VX_lsu_unit.sv:271:27
								rsp_data[i * 32+:32] = sv2v_cast_32($unsigned(rsp_data8));
							3'b101:
								// Trace: ../../rtl/VX_lsu_unit.sv:272:27
								rsp_data[i * 32+:32] = sv2v_cast_32($unsigned(rsp_data16));
							default:
								// Trace: ../../rtl/VX_lsu_unit.sv:273:22
								rsp_data[i * 32+:32] = rsp_data32;
						endcase
				end
				// Trace: ../../rtl/VX_lsu_unit.sv:278:5
				assign rsp_tmask_qual = (rsp_is_dup ? rsp_tmask : VX_pipeline.dcache_rsp_if.tmask);
				// Trace: ../../rtl/VX_lsu_unit.sv:282:5
				wire load_rsp_stall = ~VX_pipeline.ld_commit_if.ready && VX_pipeline.ld_commit_if.valid;
				// Trace: ../../rtl/VX_lsu_unit.sv:284:5
				VX_pipe_register #(
					.DATAW(151),
					.RESETW(1)
				) rsp_pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(!load_rsp_stall),
					.data_in({VX_pipeline.dcache_rsp_if.valid, rsp_uuid, rsp_wid, rsp_tmask_qual, rsp_pc, rsp_rd, rsp_wb, rsp_data, mbuf_pop}),
					.data_out({VX_pipeline.ld_commit_if.valid, VX_pipeline.ld_commit_if.uuid, VX_pipeline.ld_commit_if.wid, VX_pipeline.ld_commit_if.tmask, VX_pipeline.ld_commit_if.PC, VX_pipeline.ld_commit_if.rd, VX_pipeline.ld_commit_if.wb, VX_pipeline.ld_commit_if.data, VX_pipeline.ld_commit_if.eop})
				);
				// Trace: ../../rtl/VX_lsu_unit.sv:296:5
				assign VX_pipeline.dcache_rsp_if.ready = ~load_rsp_stall;
			end
			assign lsu_unit.clk = clk;
			assign lsu_unit.reset = lsu_reset;
			// Trace: ../../rtl/VX_execute.sv:166:5
			// expanded module instance: csr_unit
			localparam _param_BED2E_CORE_ID = CORE_ID;
			if (1) begin : csr_unit
				// Trace: ../../rtl/VX_csr_unit.sv:4:15
				localparam CORE_ID = _param_BED2E_CORE_ID;
				// Trace: ../../rtl/VX_csr_unit.sv:6:5
				wire clk;
				// Trace: ../../rtl/VX_csr_unit.sv:7:5
				wire reset;
				// Trace: ../../rtl/VX_csr_unit.sv:17:5
				// removed modport instance cmt_to_csr_if
				// Trace: ../../rtl/VX_csr_unit.sv:18:5
				// removed modport instance fetch_to_csr_if
				// Trace: ../../rtl/VX_csr_unit.sv:19:5
				// removed modport instance csr_req_if
				// Trace: ../../rtl/VX_csr_unit.sv:20:5
				// removed modport instance csr_commit_if
				// Trace: ../../rtl/VX_csr_unit.sv:30:5
				wire [1:0] pending;
				// Trace: ../../rtl/VX_csr_unit.sv:31:5
				wire busy;
				// Trace: ../../rtl/VX_csr_unit.sv:33:5
				wire csr_we_s1;
				// Trace: ../../rtl/VX_csr_unit.sv:34:5
				wire [11:0] csr_addr_s1;
				// Trace: ../../rtl/VX_csr_unit.sv:35:5
				wire [31:0] csr_read_data;
				// Trace: ../../rtl/VX_csr_unit.sv:36:5
				wire [31:0] csr_read_data_s1;
				// Trace: ../../rtl/VX_csr_unit.sv:37:5
				wire [31:0] csr_updated_data_s1;
				// Trace: ../../rtl/VX_csr_unit.sv:39:5
				wire write_enable = VX_pipeline.csr_commit_if.valid && csr_we_s1;
				// Trace: ../../rtl/VX_csr_unit.sv:41:5
				wire [31:0] csr_req_data = (VX_pipeline.csr_req_if.use_imm ? sv2v_cast_32(VX_pipeline.csr_req_if.imm) : VX_pipeline.csr_req_if.rs1_data);
				// Trace: ../../rtl/VX_csr_unit.sv:43:5
				// expanded module instance: csr_data
				localparam _param_9D0B6_CORE_ID = CORE_ID;
				if (1) begin : csr_data
					// Trace: ../../rtl/VX_csr_data.sv:4:15
					localparam CORE_ID = _param_9D0B6_CORE_ID;
					// Trace: ../../rtl/VX_csr_data.sv:6:5
					wire clk;
					// Trace: ../../rtl/VX_csr_data.sv:7:5
					wire reset;
					// Trace: ../../rtl/VX_csr_data.sv:17:5
					// removed modport instance cmt_to_csr_if
					// Trace: ../../rtl/VX_csr_data.sv:18:5
					// removed modport instance fetch_to_csr_if
					// Trace: ../../rtl/VX_csr_data.sv:27:5
					wire read_enable;
					// Trace: ../../rtl/VX_csr_data.sv:28:5
					wire [43:0] read_uuid;
					// Trace: ../../rtl/VX_csr_data.sv:29:5
					wire [11:0] read_addr;
					// Trace: ../../rtl/VX_csr_data.sv:30:5
					wire [0:0] read_wid;
					// Trace: ../../rtl/VX_csr_data.sv:31:5
					wire [31:0] read_data;
					// Trace: ../../rtl/VX_csr_data.sv:33:5
					wire write_enable;
					// Trace: ../../rtl/VX_csr_data.sv:34:5
					wire [43:0] write_uuid;
					// Trace: ../../rtl/VX_csr_data.sv:35:5
					wire [11:0] write_addr;
					// Trace: ../../rtl/VX_csr_data.sv:36:5
					wire [0:0] write_wid;
					// Trace: ../../rtl/VX_csr_data.sv:37:5
					wire [31:0] write_data;
					// Trace: ../../rtl/VX_csr_data.sv:39:5
					wire busy;
					// Trace: ../../rtl/VX_csr_data.sv:41:5
					// removed import fpu_types::*;
					// Trace: ../../rtl/VX_csr_data.sv:43:5
					reg [11:0] csr_satp;
					// Trace: ../../rtl/VX_csr_data.sv:44:5
					reg [11:0] csr_mstatus;
					// Trace: ../../rtl/VX_csr_data.sv:45:5
					reg [11:0] csr_medeleg;
					// Trace: ../../rtl/VX_csr_data.sv:46:5
					reg [11:0] csr_mideleg;
					// Trace: ../../rtl/VX_csr_data.sv:47:5
					reg [11:0] csr_mie;
					// Trace: ../../rtl/VX_csr_data.sv:48:5
					reg [11:0] csr_mtvec;
					// Trace: ../../rtl/VX_csr_data.sv:49:5
					reg [11:0] csr_mepc;
					// Trace: ../../rtl/VX_csr_data.sv:50:5
					reg [11:0] csr_pmpcfg [0:0];
					// Trace: ../../rtl/VX_csr_data.sv:51:5
					reg [11:0] csr_pmpaddr [0:0];
					// Trace: ../../rtl/VX_csr_data.sv:52:5
					reg [63:0] csr_cycle;
					// Trace: ../../rtl/VX_csr_data.sv:53:5
					reg [63:0] csr_instret;
					// Trace: ../../rtl/VX_csr_data.sv:55:5
					// removed localparam type fpu_types_fflags_t
					reg [15:0] fcsr;
					// Trace: ../../rtl/VX_csr_data.sv:57:5
					always @(posedge clk)
						// Trace: ../../rtl/VX_csr_data.sv:58:9
						if (reset)
							// Trace: ../../rtl/VX_csr_data.sv:59:13
							fcsr <= 1'sb0;
						else
							// Trace: ../../rtl/VX_csr_data.sv:67:13
							if (write_enable)
								// Trace: ../../rtl/VX_csr_data.sv:68:17
								case (write_addr)
									12'h001:
										// Trace: ../../rtl/VX_csr_data.sv:69:36
										fcsr[(write_wid * 8) + 4-:5] <= write_data[4:0];
									12'h002:
										// Trace: ../../rtl/VX_csr_data.sv:70:36
										fcsr[(write_wid * 8) + 7-:3] <= write_data[2:0];
									12'h003:
										// Trace: ../../rtl/VX_csr_data.sv:71:36
										fcsr[write_wid * 8+:8] <= write_data[7:0];
									12'h180:
										// Trace: ../../rtl/VX_csr_data.sv:72:36
										csr_satp <= write_data[11:0];
									12'h300:
										// Trace: ../../rtl/VX_csr_data.sv:73:36
										csr_mstatus <= write_data[11:0];
									12'h302:
										// Trace: ../../rtl/VX_csr_data.sv:74:36
										csr_medeleg <= write_data[11:0];
									12'h303:
										// Trace: ../../rtl/VX_csr_data.sv:75:36
										csr_mideleg <= write_data[11:0];
									12'h304:
										// Trace: ../../rtl/VX_csr_data.sv:76:36
										csr_mie <= write_data[11:0];
									12'h305:
										// Trace: ../../rtl/VX_csr_data.sv:77:36
										csr_mtvec <= write_data[11:0];
									12'h341:
										// Trace: ../../rtl/VX_csr_data.sv:78:36
										csr_mepc <= write_data[11:0];
									12'h3a0:
										// Trace: ../../rtl/VX_csr_data.sv:79:36
										csr_pmpcfg[0] <= write_data[11:0];
									12'h3b0:
										// Trace: ../../rtl/VX_csr_data.sv:80:36
										csr_pmpaddr[0] <= write_data[11:0];
									default:
										// Trace: macro expansion of ASSERT at ../../rtl/VX_csr_data.sv:88:122
										if (~write_enable)
											;
								endcase
					// Trace: ../../rtl/VX_csr_data.sv:106:5
					always @(posedge clk)
						// Trace: ../../rtl/VX_csr_data.sv:107:8
						if (reset) begin
							// Trace: ../../rtl/VX_csr_data.sv:108:13
							csr_cycle <= 0;
							// Trace: ../../rtl/VX_csr_data.sv:109:13
							csr_instret <= 0;
						end
						else begin
							// Trace: ../../rtl/VX_csr_data.sv:111:13
							if (busy)
								// Trace: ../../rtl/VX_csr_data.sv:112:17
								csr_cycle <= csr_cycle + 1;
							if (VX_pipeline.cmt_to_csr_if.valid)
								// Trace: ../../rtl/VX_csr_data.sv:115:17
								csr_instret <= csr_instret + sv2v_cast_64(VX_pipeline.cmt_to_csr_if.commit_size);
						end
					// Trace: ../../rtl/VX_csr_data.sv:120:5
					reg [31:0] read_data_r;
					// Trace: ../../rtl/VX_csr_data.sv:121:5
					reg read_addr_valid_r;
					// Trace: ../../rtl/VX_csr_data.sv:123:5
					always @(*) begin
						// Trace: ../../rtl/VX_csr_data.sv:124:9
						read_data_r = 1'sbx;
						// Trace: ../../rtl/VX_csr_data.sv:125:9
						read_addr_valid_r = 1;
						// Trace: ../../rtl/VX_csr_data.sv:126:9
						case (read_addr)
							12'h001:
								// Trace: ../../rtl/VX_csr_data.sv:127:31
								read_data_r = sv2v_cast_32(fcsr[(read_wid * 8) + 4-:5]);
							12'h002:
								// Trace: ../../rtl/VX_csr_data.sv:128:31
								read_data_r = sv2v_cast_32(fcsr[(read_wid * 8) + 7-:3]);
							12'h003:
								// Trace: ../../rtl/VX_csr_data.sv:129:31
								read_data_r = sv2v_cast_32(fcsr[read_wid * 8+:8]);
							12'hcc0, 12'hcc1, 12'hcc3:
								// Trace: ../../rtl/VX_csr_data.sv:133:31
								read_data_r = sv2v_cast_32(read_wid);
							12'hcc2, 12'hf14:
								// Trace: ../../rtl/VX_csr_data.sv:136:31
								read_data_r = (CORE_ID * 2) + sv2v_cast_32(read_wid);
							12'hcc5:
								// Trace: ../../rtl/VX_csr_data.sv:137:31
								read_data_r = CORE_ID;
							12'hcc4:
								// Trace: ../../rtl/VX_csr_data.sv:139:31
								read_data_r = sv2v_cast_32(VX_pipeline.fetch_to_csr_if.thread_masks[read_wid * 2+:2]);
							12'hfc0:
								// Trace: ../../rtl/VX_csr_data.sv:141:31
								read_data_r = 2;
							12'hfc1:
								// Trace: ../../rtl/VX_csr_data.sv:142:31
								read_data_r = 2;
							12'hfc2:
								// Trace: ../../rtl/VX_csr_data.sv:143:31
								read_data_r = 1;
							12'hb00:
								// Trace: ../../rtl/VX_csr_data.sv:145:31
								read_data_r = csr_cycle[31:0];
							12'hb80:
								// Trace: ../../rtl/VX_csr_data.sv:146:31
								read_data_r = sv2v_cast_32(csr_cycle[43:32]);
							12'hb02:
								// Trace: ../../rtl/VX_csr_data.sv:147:31
								read_data_r = csr_instret[31:0];
							12'hb82:
								// Trace: ../../rtl/VX_csr_data.sv:148:31
								read_data_r = sv2v_cast_32(csr_instret[43:32]);
							12'h180:
								// Trace: ../../rtl/VX_csr_data.sv:222:30
								read_data_r = sv2v_cast_32(csr_satp);
							12'h300:
								// Trace: ../../rtl/VX_csr_data.sv:224:30
								read_data_r = sv2v_cast_32(csr_mstatus);
							12'h301:
								// Trace: ../../rtl/VX_csr_data.sv:225:30
								read_data_r = 9441536;
							12'h302:
								// Trace: ../../rtl/VX_csr_data.sv:226:30
								read_data_r = sv2v_cast_32(csr_medeleg);
							12'h303:
								// Trace: ../../rtl/VX_csr_data.sv:227:30
								read_data_r = sv2v_cast_32(csr_mideleg);
							12'h304:
								// Trace: ../../rtl/VX_csr_data.sv:228:30
								read_data_r = sv2v_cast_32(csr_mie);
							12'h305:
								// Trace: ../../rtl/VX_csr_data.sv:229:30
								read_data_r = sv2v_cast_32(csr_mtvec);
							12'h341:
								// Trace: ../../rtl/VX_csr_data.sv:231:30
								read_data_r = sv2v_cast_32(csr_mepc);
							12'h3a0:
								// Trace: ../../rtl/VX_csr_data.sv:233:30
								read_data_r = sv2v_cast_32(csr_pmpcfg[0]);
							12'h3b0:
								// Trace: ../../rtl/VX_csr_data.sv:234:30
								read_data_r = sv2v_cast_32(csr_pmpaddr[0]);
							12'hf11:
								// Trace: ../../rtl/VX_csr_data.sv:236:30
								read_data_r = 0;
							12'hf12:
								// Trace: ../../rtl/VX_csr_data.sv:237:30
								read_data_r = 0;
							12'hf13:
								// Trace: ../../rtl/VX_csr_data.sv:238:30
								read_data_r = 0;
							default:
								// Trace: ../../rtl/VX_csr_data.sv:241:17
								if (((read_addr >= 12'hb00) && (read_addr < 2848)) || ((read_addr >= 12'hb80) && (read_addr < 2976)))
									// Trace: ../../rtl/VX_csr_data.sv:243:22
									read_addr_valid_r = 1;
								else
									// Trace: ../../rtl/VX_csr_data.sv:252:21
									read_addr_valid_r = 0;
						endcase
					end
					// Trace: ../../rtl/VX_csr_data.sv:259:5
					assign read_data = read_data_r;
				end
				assign csr_data.clk = clk;
				assign csr_data.reset = reset;
				assign csr_data.read_enable = VX_pipeline.csr_req_if.valid;
				assign csr_data.read_uuid = VX_pipeline.csr_req_if.uuid;
				assign csr_data.read_addr = VX_pipeline.csr_req_if.addr;
				assign csr_data.read_wid = VX_pipeline.csr_req_if.wid;
				assign csr_read_data = csr_data.read_data;
				assign csr_data.write_enable = write_enable;
				assign csr_data.write_uuid = VX_pipeline.csr_commit_if.uuid;
				assign csr_data.write_addr = csr_addr_s1;
				assign csr_data.write_wid = VX_pipeline.csr_commit_if.wid;
				assign csr_data.write_data = csr_updated_data_s1;
				assign csr_data.busy = busy;
				// Trace: ../../rtl/VX_csr_unit.sv:76:5
				wire write_hazard = ((csr_addr_s1 == VX_pipeline.csr_req_if.addr) && (VX_pipeline.csr_commit_if.wid == VX_pipeline.csr_req_if.wid)) && VX_pipeline.csr_commit_if.valid;
				// Trace: ../../rtl/VX_csr_unit.sv:80:5
				wire [31:0] csr_read_data_qual = (write_hazard ? csr_updated_data_s1 : csr_read_data);
				// Trace: ../../rtl/VX_csr_unit.sv:82:5
				reg [31:0] csr_updated_data;
				// Trace: ../../rtl/VX_csr_unit.sv:83:5
				reg csr_we_s0_unqual;
				// Trace: ../../rtl/VX_csr_unit.sv:85:5
				always @(*) begin
					// Trace: ../../rtl/VX_csr_unit.sv:86:9
					csr_we_s0_unqual = csr_req_data != 0;
					// Trace: ../../rtl/VX_csr_unit.sv:87:9
					case (VX_pipeline.csr_req_if.op_type)
						2'h1: begin
							// Trace: ../../rtl/VX_csr_unit.sv:89:17
							csr_updated_data = csr_req_data;
							// Trace: ../../rtl/VX_csr_unit.sv:90:17
							csr_we_s0_unqual = 1;
						end
						2'h2:
							// Trace: ../../rtl/VX_csr_unit.sv:93:17
							csr_updated_data = csr_read_data_qual | csr_req_data;
						default:
							// Trace: ../../rtl/VX_csr_unit.sv:97:17
							csr_updated_data = csr_read_data_qual & ~csr_req_data;
					endcase
				end
				// Trace: ../../rtl/VX_csr_unit.sv:105:5
				wire stall_in = 0;
				// Trace: ../../rtl/VX_csr_unit.sv:108:5
				wire csr_req_valid = VX_pipeline.csr_req_if.valid && !stall_in;
				// Trace: ../../rtl/VX_csr_unit.sv:110:5
				wire stall_out = ~VX_pipeline.csr_commit_if.ready && VX_pipeline.csr_commit_if.valid;
				// Trace: ../../rtl/VX_csr_unit.sv:112:5
				VX_pipe_register #(
					.DATAW(163),
					.RESETW(1)
				) pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(!stall_out),
					.data_in({csr_req_valid, VX_pipeline.csr_req_if.uuid, VX_pipeline.csr_req_if.wid, VX_pipeline.csr_req_if.tmask, VX_pipeline.csr_req_if.PC, VX_pipeline.csr_req_if.rd, VX_pipeline.csr_req_if.wb, csr_we_s0_unqual, VX_pipeline.csr_req_if.addr, csr_read_data_qual, csr_updated_data}),
					.data_out({VX_pipeline.csr_commit_if.valid, VX_pipeline.csr_commit_if.uuid, VX_pipeline.csr_commit_if.wid, VX_pipeline.csr_commit_if.tmask, VX_pipeline.csr_commit_if.PC, VX_pipeline.csr_commit_if.rd, VX_pipeline.csr_commit_if.wb, csr_we_s1, csr_addr_s1, csr_read_data_s1, csr_updated_data_s1})
				);
				// Trace: ../../rtl/VX_csr_unit.sv:123:5
				genvar i;
				for (i = 0; i < 2; i = i + 1) begin : genblk1
					// Trace: ../../rtl/VX_csr_unit.sv:124:9
					assign VX_pipeline.csr_commit_if.data[i * 32+:32] = (csr_addr_s1 == 12'hcc0 ? i : ((csr_addr_s1 == 12'hcc1) || (csr_addr_s1 == 12'hcc2) ? (csr_read_data_s1 * 2) + i : csr_read_data_s1));
				end
				// Trace: ../../rtl/VX_csr_unit.sv:130:5
				assign VX_pipeline.csr_commit_if.eop = 1'b1;
				// Trace: ../../rtl/VX_csr_unit.sv:133:5
				assign VX_pipeline.csr_req_if.ready = ~(stall_out || stall_in);
				// Trace: ../../rtl/VX_csr_unit.sv:136:5
				reg [1:0] pending_r;
				// Trace: ../../rtl/VX_csr_unit.sv:137:5
				always @(posedge clk)
					// Trace: ../../rtl/VX_csr_unit.sv:138:9
					if (reset)
						// Trace: ../../rtl/VX_csr_unit.sv:139:13
						pending_r <= 0;
					else begin
						// Trace: ../../rtl/VX_csr_unit.sv:141:13
						if (VX_pipeline.csr_commit_if.valid && VX_pipeline.csr_commit_if.ready)
							// Trace: ../../rtl/VX_csr_unit.sv:142:18
							pending_r[VX_pipeline.csr_commit_if.wid] <= 0;
						if (VX_pipeline.csr_req_if.valid && VX_pipeline.csr_req_if.ready)
							// Trace: ../../rtl/VX_csr_unit.sv:145:18
							pending_r[VX_pipeline.csr_req_if.wid] <= 1;
					end
				// Trace: ../../rtl/VX_csr_unit.sv:149:5
				assign pending = pending_r;
			end
			assign csr_unit.clk = clk;
			assign csr_unit.reset = csr_reset;
			assign csr_unit.busy = busy;
			// Trace: ../../rtl/VX_execute.sv:211:5
			// expanded module instance: gpu_unit
			localparam _param_FC85A_CORE_ID = CORE_ID;
			if (1) begin : gpu_unit
				// Trace: ../../rtl/VX_gpu_unit.sv:4:15
				localparam CORE_ID = _param_FC85A_CORE_ID;
				// Trace: ../../rtl/VX_gpu_unit.sv:8:5
				wire clk;
				// Trace: ../../rtl/VX_gpu_unit.sv:9:5
				wire reset;
				// Trace: ../../rtl/VX_gpu_unit.sv:12:5
				// removed modport instance gpu_req_if
				// Trace: ../../rtl/VX_gpu_unit.sv:25:5
				// removed modport instance warp_ctl_if
				// Trace: ../../rtl/VX_gpu_unit.sv:26:5
				// removed modport instance gpu_commit_if
				// Trace: ../../rtl/VX_gpu_unit.sv:28:5
				// removed import gpu_types::*;
				// Trace: ../../rtl/VX_gpu_unit.sv:32:5
				// removed localparam type gpu_types_gpu_barrier_t
				// removed localparam type gpu_types_gpu_split_t
				// removed localparam type gpu_types_gpu_tmc_t
				// removed localparam type gpu_types_gpu_wspawn_t
				localparam WCTL_DATAW = 80;
				// Trace: ../../rtl/VX_gpu_unit.sv:33:5
				localparam RSP_DATAW = WCTL_DATAW;
				// Trace: ../../rtl/VX_gpu_unit.sv:35:5
				wire rsp_valid;
				// Trace: ../../rtl/VX_gpu_unit.sv:36:5
				wire [43:0] rsp_uuid;
				// Trace: ../../rtl/VX_gpu_unit.sv:37:5
				wire [0:0] rsp_wid;
				// Trace: ../../rtl/VX_gpu_unit.sv:38:5
				wire [1:0] rsp_tmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:39:5
				wire [31:0] rsp_PC;
				// Trace: ../../rtl/VX_gpu_unit.sv:40:5
				wire [4:0] rsp_rd;
				// Trace: ../../rtl/VX_gpu_unit.sv:41:5
				wire rsp_wb;
				// Trace: ../../rtl/VX_gpu_unit.sv:43:5
				wire [79:0] rsp_data;
				wire [79:0] rsp_data_r;
				// Trace: ../../rtl/VX_gpu_unit.sv:45:5
				wire [2:0] tmc;
				// Trace: ../../rtl/VX_gpu_unit.sv:46:5
				wire [34:0] wspawn;
				// Trace: ../../rtl/VX_gpu_unit.sv:47:5
				wire [3:0] barrier;
				// Trace: ../../rtl/VX_gpu_unit.sv:48:5
				wire [37:0] split;
				// Trace: ../../rtl/VX_gpu_unit.sv:50:5
				wire [79:0] warp_ctl_data;
				// Trace: ../../rtl/VX_gpu_unit.sv:51:5
				wire is_warp_ctl;
				// Trace: ../../rtl/VX_gpu_unit.sv:53:5
				wire stall_in;
				wire stall_out;
				// Trace: ../../rtl/VX_gpu_unit.sv:55:5
				wire is_wspawn = VX_pipeline.gpu_req_if.op_type == 4'h1;
				// Trace: ../../rtl/VX_gpu_unit.sv:56:5
				wire is_tmc = VX_pipeline.gpu_req_if.op_type == 4'h0;
				// Trace: ../../rtl/VX_gpu_unit.sv:57:5
				wire is_split = VX_pipeline.gpu_req_if.op_type == 4'h2;
				// Trace: ../../rtl/VX_gpu_unit.sv:58:5
				wire is_bar = VX_pipeline.gpu_req_if.op_type == 4'h4;
				// Trace: ../../rtl/VX_gpu_unit.sv:59:5
				wire is_pred = VX_pipeline.gpu_req_if.op_type == 4'h5;
				// Trace: ../../rtl/VX_gpu_unit.sv:61:5
				wire [31:0] rs1_data = VX_pipeline.gpu_req_if.rs1_data[VX_pipeline.gpu_req_if.tid * 32+:32];
				// Trace: ../../rtl/VX_gpu_unit.sv:62:5
				wire [31:0] rs2_data = VX_pipeline.gpu_req_if.rs2_data[VX_pipeline.gpu_req_if.tid * 32+:32];
				// Trace: ../../rtl/VX_gpu_unit.sv:64:5
				wire [1:0] taken_tmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:65:5
				wire [1:0] not_taken_tmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:67:5
				genvar i;
				for (i = 0; i < 2; i = i + 1) begin : genblk1
					// Trace: ../../rtl/VX_gpu_unit.sv:68:9
					wire taken = VX_pipeline.gpu_req_if.rs1_data[i * 32+:32] != 0;
					// Trace: ../../rtl/VX_gpu_unit.sv:69:9
					assign taken_tmask[i] = VX_pipeline.gpu_req_if.tmask[i] & taken;
					// Trace: ../../rtl/VX_gpu_unit.sv:70:9
					assign not_taken_tmask[i] = VX_pipeline.gpu_req_if.tmask[i] & ~taken;
				end
				// Trace: ../../rtl/VX_gpu_unit.sv:75:5
				wire [1:0] pred_mask = (taken_tmask != 0 ? taken_tmask : VX_pipeline.gpu_req_if.tmask);
				// Trace: ../../rtl/VX_gpu_unit.sv:77:5
				assign tmc[2] = is_tmc || is_pred;
				// Trace: ../../rtl/VX_gpu_unit.sv:78:5
				assign tmc[1-:2] = (is_pred ? pred_mask : rs1_data[1:0]);
				// Trace: ../../rtl/VX_gpu_unit.sv:82:5
				wire [31:0] wspawn_pc = rs2_data;
				// Trace: ../../rtl/VX_gpu_unit.sv:83:5
				wire [1:0] wspawn_wmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:84:5
				for (i = 0; i < 2; i = i + 1) begin : genblk2
					// Trace: ../../rtl/VX_gpu_unit.sv:85:9
					assign wspawn_wmask[i] = i < rs1_data;
				end
				// Trace: ../../rtl/VX_gpu_unit.sv:87:5
				assign wspawn[34] = is_wspawn;
				// Trace: ../../rtl/VX_gpu_unit.sv:88:5
				assign wspawn[33-:2] = wspawn_wmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:89:5
				assign wspawn[31-:32] = wspawn_pc;
				// Trace: ../../rtl/VX_gpu_unit.sv:93:5
				assign split[37] = is_split;
				// Trace: ../../rtl/VX_gpu_unit.sv:94:5
				assign split[36] = |taken_tmask && |not_taken_tmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:95:5
				assign split[35-:2] = taken_tmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:96:5
				assign split[33-:2] = not_taken_tmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:97:5
				assign split[31-:32] = VX_pipeline.gpu_req_if.next_PC;
				// Trace: ../../rtl/VX_gpu_unit.sv:101:5
				assign barrier[3] = is_bar;
				// Trace: ../../rtl/VX_gpu_unit.sv:102:5
				assign barrier[2-:2] = rs1_data[1:0];
				// Trace: ../../rtl/VX_gpu_unit.sv:103:5
				assign barrier[0-:1] = sv2v_cast_1(rs2_data - 1);
				// Trace: ../../rtl/VX_gpu_unit.sv:106:5
				assign warp_ctl_data = {tmc, wspawn, split, barrier};
				// Trace: ../../rtl/VX_gpu_unit.sv:170:5
				assign stall_in = stall_out;
				// Trace: ../../rtl/VX_gpu_unit.sv:171:5
				assign is_warp_ctl = 1;
				// Trace: ../../rtl/VX_gpu_unit.sv:173:5
				assign rsp_valid = VX_pipeline.gpu_req_if.valid;
				// Trace: ../../rtl/VX_gpu_unit.sv:174:5
				assign rsp_uuid = VX_pipeline.gpu_req_if.uuid;
				// Trace: ../../rtl/VX_gpu_unit.sv:175:5
				assign rsp_wid = VX_pipeline.gpu_req_if.wid;
				// Trace: ../../rtl/VX_gpu_unit.sv:176:5
				assign rsp_tmask = VX_pipeline.gpu_req_if.tmask;
				// Trace: ../../rtl/VX_gpu_unit.sv:177:5
				assign rsp_PC = VX_pipeline.gpu_req_if.PC;
				// Trace: ../../rtl/VX_gpu_unit.sv:178:5
				assign rsp_rd = 0;
				// Trace: ../../rtl/VX_gpu_unit.sv:179:5
				assign rsp_wb = 0;
				// Trace: ../../rtl/VX_gpu_unit.sv:180:5
				function automatic [79:0] sv2v_cast_790CE;
					input reg [79:0] inp;
					sv2v_cast_790CE = inp;
				endfunction
				assign rsp_data = sv2v_cast_790CE(warp_ctl_data);
				// Trace: ../../rtl/VX_gpu_unit.sv:184:5
				wire is_warp_ctl_r;
				// Trace: ../../rtl/VX_gpu_unit.sv:187:5
				assign stall_out = ~VX_pipeline.gpu_commit_if.ready && VX_pipeline.gpu_commit_if.valid;
				// Trace: ../../rtl/VX_gpu_unit.sv:189:5
				VX_pipe_register #(
					.DATAW(167),
					.RESETW(1)
				) pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(!stall_out),
					.data_in({rsp_valid, rsp_uuid, rsp_wid, rsp_tmask, rsp_PC, rsp_rd, rsp_wb, rsp_data, is_warp_ctl}),
					.data_out({VX_pipeline.gpu_commit_if.valid, VX_pipeline.gpu_commit_if.uuid, VX_pipeline.gpu_commit_if.wid, VX_pipeline.gpu_commit_if.tmask, VX_pipeline.gpu_commit_if.PC, VX_pipeline.gpu_commit_if.rd, VX_pipeline.gpu_commit_if.wb, rsp_data_r, is_warp_ctl_r})
				);
				// Trace: ../../rtl/VX_gpu_unit.sv:200:5
				assign VX_pipeline.gpu_commit_if.data = rsp_data_r[63:0];
				// Trace: ../../rtl/VX_gpu_unit.sv:201:5
				assign VX_pipeline.gpu_commit_if.eop = 1'b1;
				// Trace: ../../rtl/VX_gpu_unit.sv:205:5
				assign {VX_pipeline.warp_ctl_if.tmc, VX_pipeline.warp_ctl_if.wspawn, VX_pipeline.warp_ctl_if.split, VX_pipeline.warp_ctl_if.barrier} = rsp_data_r[79:0];
				// Trace: ../../rtl/VX_gpu_unit.sv:207:5
				assign VX_pipeline.warp_ctl_if.valid = (VX_pipeline.gpu_commit_if.valid && VX_pipeline.gpu_commit_if.ready) && is_warp_ctl_r;
				// Trace: ../../rtl/VX_gpu_unit.sv:208:5
				assign VX_pipeline.warp_ctl_if.wid = VX_pipeline.gpu_commit_if.wid;
				// Trace: ../../rtl/VX_gpu_unit.sv:211:5
				assign VX_pipeline.gpu_req_if.ready = ~stall_in;
			end
			assign gpu_unit.clk = clk;
			assign gpu_unit.reset = gpu_reset;
			// Trace: ../../rtl/VX_execute.sv:231:5
			wire ebreak;
			// Trace: ../../rtl/VX_execute.sv:232:5
			assign ebreak = ((VX_pipeline.alu_req_if.valid && VX_pipeline.alu_req_if.ready) && VX_pipeline.alu_req_if.op_mod[0]) && ((VX_pipeline.alu_req_if.op_type == 4'b1011) || (VX_pipeline.alu_req_if.op_type == 4'b1010));
		end
	endgenerate
	assign execute.clk = clk;
	assign execute.reset = execute_reset;
	assign execute.busy = busy;
	// Trace: ../../rtl/VX_pipeline.sv:242:5
	// expanded module instance: commit
	localparam _param_D837E_CORE_ID = CORE_ID;
	generate
		if (1) begin : commit
			// Trace: ../../rtl/VX_commit.sv:4:15
			localparam CORE_ID = _param_D837E_CORE_ID;
			// Trace: ../../rtl/VX_commit.sv:6:5
			wire clk;
			// Trace: ../../rtl/VX_commit.sv:7:5
			wire reset;
			// Trace: ../../rtl/VX_commit.sv:10:5
			// removed modport instance alu_commit_if
			// Trace: ../../rtl/VX_commit.sv:11:5
			// removed modport instance ld_commit_if
			// Trace: ../../rtl/VX_commit.sv:12:5
			// removed modport instance st_commit_if
			// Trace: ../../rtl/VX_commit.sv:13:5
			// removed modport instance csr_commit_if
			// Trace: ../../rtl/VX_commit.sv:17:5
			// removed modport instance gpu_commit_if
			// Trace: ../../rtl/VX_commit.sv:20:5
			// removed modport instance writeback_if
			// Trace: ../../rtl/VX_commit.sv:21:5
			// removed modport instance cmt_to_csr_if
			// Trace: ../../rtl/VX_commit.sv:25:5
			wire alu_commit_fire = VX_pipeline.alu_commit_if.valid && VX_pipeline.alu_commit_if.ready;
			// Trace: ../../rtl/VX_commit.sv:26:5
			wire ld_commit_fire = VX_pipeline.ld_commit_if.valid && VX_pipeline.ld_commit_if.ready;
			// Trace: ../../rtl/VX_commit.sv:27:5
			wire st_commit_fire = VX_pipeline.st_commit_if.valid && VX_pipeline.st_commit_if.ready;
			// Trace: ../../rtl/VX_commit.sv:28:5
			wire csr_commit_fire = VX_pipeline.csr_commit_if.valid && VX_pipeline.csr_commit_if.ready;
			// Trace: ../../rtl/VX_commit.sv:32:5
			wire gpu_commit_fire = VX_pipeline.gpu_commit_if.valid && VX_pipeline.gpu_commit_if.ready;
			// Trace: ../../rtl/VX_commit.sv:34:5
			wire commit_fire = (((alu_commit_fire || ld_commit_fire) || st_commit_fire) || csr_commit_fire) || gpu_commit_fire;
			// Trace: ../../rtl/VX_commit.sv:46:5
			wire [9:0] commit_tmask;
			// Trace: ../../rtl/VX_commit.sv:49:5
			wire [3:0] commit_size;
			// Trace: ../../rtl/VX_commit.sv:51:5
			assign commit_tmask = {{2 {alu_commit_fire}} & VX_pipeline.alu_commit_if.tmask, {2 {ld_commit_fire}} & VX_pipeline.ld_commit_if.tmask, {2 {st_commit_fire}} & VX_pipeline.st_commit_if.tmask, {2 {csr_commit_fire}} & VX_pipeline.csr_commit_if.tmask, {2 {gpu_commit_fire}} & VX_pipeline.gpu_commit_if.tmask};
			// Trace: macro expansion of POP_COUNT at ../../rtl/VX_commit.sv:62:37
			VX_popcount #(.N(10)) __commit_size(
				.in_i(commit_tmask),
				.cnt_o(commit_size)
			);
			// Trace: ../../rtl/VX_commit.sv:64:5
			VX_pipe_register #(
				.DATAW(5),
				.RESETW(1)
			) pipe_reg(
				.clk(clk),
				.reset(reset),
				.enable(1'b1),
				.data_in({commit_fire, commit_size}),
				.data_out({VX_pipeline.cmt_to_csr_if.valid, VX_pipeline.cmt_to_csr_if.commit_size})
			);
			// Trace: ../../rtl/VX_commit.sv:77:5
			// expanded module instance: writeback
			localparam _param_35426_CORE_ID = CORE_ID;
			if (1) begin : writeback
				// Trace: ../../rtl/VX_writeback.sv:4:15
				localparam CORE_ID = _param_35426_CORE_ID;
				// Trace: ../../rtl/VX_writeback.sv:6:5
				wire clk;
				// Trace: ../../rtl/VX_writeback.sv:7:5
				wire reset;
				// Trace: ../../rtl/VX_writeback.sv:10:5
				// removed modport instance alu_commit_if
				// Trace: ../../rtl/VX_writeback.sv:11:5
				// removed modport instance ld_commit_if
				// Trace: ../../rtl/VX_writeback.sv:12:5
				// removed modport instance csr_commit_if
				// Trace: ../../rtl/VX_writeback.sv:16:5
				// removed modport instance gpu_commit_if
				// Trace: ../../rtl/VX_writeback.sv:19:5
				// removed modport instance writeback_if
				// Trace: ../../rtl/VX_writeback.sv:24:5
				localparam DATAW = 105;
				// Trace: ../../rtl/VX_writeback.sv:28:5
				localparam NUM_RSPS = 4;
				// Trace: ../../rtl/VX_writeback.sv:31:5
				wire wb_valid;
				// Trace: ../../rtl/VX_writeback.sv:32:5
				wire [0:0] wb_wid;
				// Trace: ../../rtl/VX_writeback.sv:33:5
				wire [31:0] wb_PC;
				// Trace: ../../rtl/VX_writeback.sv:34:5
				wire [1:0] wb_tmask;
				// Trace: ../../rtl/VX_writeback.sv:35:5
				wire [4:0] wb_rd;
				// Trace: ../../rtl/VX_writeback.sv:36:5
				wire [63:0] wb_data;
				// Trace: ../../rtl/VX_writeback.sv:37:5
				wire wb_eop;
				// Trace: ../../rtl/VX_writeback.sv:39:5
				wire [3:0] rsp_valid;
				// Trace: ../../rtl/VX_writeback.sv:40:5
				wire [419:0] rsp_data;
				// Trace: ../../rtl/VX_writeback.sv:41:5
				wire [3:0] rsp_ready;
				// Trace: ../../rtl/VX_writeback.sv:42:5
				wire stall;
				// Trace: ../../rtl/VX_writeback.sv:44:5
				assign rsp_valid = {VX_pipeline.gpu_commit_if.valid && VX_pipeline.gpu_commit_if.wb, VX_pipeline.csr_commit_if.valid && VX_pipeline.csr_commit_if.wb, VX_pipeline.alu_commit_if.valid && VX_pipeline.alu_commit_if.wb, VX_pipeline.ld_commit_if.valid && VX_pipeline.ld_commit_if.wb};
				// Trace: ../../rtl/VX_writeback.sv:54:5
				assign rsp_data = {VX_pipeline.gpu_commit_if.wid, VX_pipeline.gpu_commit_if.PC, VX_pipeline.gpu_commit_if.tmask, VX_pipeline.gpu_commit_if.rd, VX_pipeline.gpu_commit_if.data, VX_pipeline.gpu_commit_if.eop, VX_pipeline.csr_commit_if.wid, VX_pipeline.csr_commit_if.PC, VX_pipeline.csr_commit_if.tmask, VX_pipeline.csr_commit_if.rd, VX_pipeline.csr_commit_if.data, VX_pipeline.csr_commit_if.eop, VX_pipeline.alu_commit_if.wid, VX_pipeline.alu_commit_if.PC, VX_pipeline.alu_commit_if.tmask, VX_pipeline.alu_commit_if.rd, VX_pipeline.alu_commit_if.data, VX_pipeline.alu_commit_if.eop, VX_pipeline.ld_commit_if.wid, VX_pipeline.ld_commit_if.PC, VX_pipeline.ld_commit_if.tmask, VX_pipeline.ld_commit_if.rd, VX_pipeline.ld_commit_if.data, VX_pipeline.ld_commit_if.eop};
				// Trace: ../../rtl/VX_writeback.sv:64:5
				VX_stream_arbiter #(
					.NUM_REQS(NUM_RSPS),
					.DATAW(DATAW),
					.BUFFERED(1),
					.TYPE("R")
				) rsp_arb(
					.clk(clk),
					.reset(reset),
					.valid_in(rsp_valid),
					.data_in(rsp_data),
					.ready_in(rsp_ready),
					.valid_out(wb_valid),
					.data_out({wb_wid, wb_PC, wb_tmask, wb_rd, wb_data, wb_eop}),
					.ready_out(~stall)
				);
				// Trace: ../../rtl/VX_writeback.sv:80:5
				assign VX_pipeline.ld_commit_if.ready = rsp_ready[0] || ~VX_pipeline.ld_commit_if.wb;
				// Trace: ../../rtl/VX_writeback.sv:87:5
				assign VX_pipeline.alu_commit_if.ready = rsp_ready[1] || ~VX_pipeline.alu_commit_if.wb;
				// Trace: ../../rtl/VX_writeback.sv:88:5
				assign VX_pipeline.csr_commit_if.ready = rsp_ready[2] || ~VX_pipeline.csr_commit_if.wb;
				// Trace: ../../rtl/VX_writeback.sv:89:5
				assign VX_pipeline.gpu_commit_if.ready = rsp_ready[3] || ~VX_pipeline.gpu_commit_if.wb;
				// Trace: ../../rtl/VX_writeback.sv:92:5
				assign stall = ~VX_pipeline.writeback_if.ready && VX_pipeline.writeback_if.valid;
				// Trace: ../../rtl/VX_writeback.sv:94:5
				VX_pipe_register #(
					.DATAW(106),
					.RESETW(1)
				) pipe_reg(
					.clk(clk),
					.reset(reset),
					.enable(~stall),
					.data_in({wb_valid, wb_wid, wb_PC, wb_tmask, wb_rd, wb_data, wb_eop}),
					.data_out({VX_pipeline.writeback_if.valid, VX_pipeline.writeback_if.wid, VX_pipeline.writeback_if.PC, VX_pipeline.writeback_if.tmask, VX_pipeline.writeback_if.rd, VX_pipeline.writeback_if.data, VX_pipeline.writeback_if.eop})
				);
				// Trace: ../../rtl/VX_writeback.sv:106:5
				reg [31:0] last_wb_value [31:0];
				// Trace: ../../rtl/VX_writeback.sv:107:5
				always @(posedge clk)
					// Trace: ../../rtl/VX_writeback.sv:108:9
					if (VX_pipeline.writeback_if.valid && VX_pipeline.writeback_if.ready)
						// Trace: ../../rtl/VX_writeback.sv:109:13
						last_wb_value[VX_pipeline.writeback_if.rd] <= VX_pipeline.writeback_if.data[0+:32];
			end
			assign writeback.clk = clk;
			assign writeback.reset = reset;
			// Trace: ../../rtl/VX_commit.sv:94:5
			assign VX_pipeline.st_commit_if.ready = 1'b1;
		end
	endgenerate
	assign commit.clk = clk;
	assign commit.reset = commit_reset;
endmodule
// removed module with interface ports: VX_scoreboard
module VX_smem_arb (
	clk,
	reset,
	req_valid_in,
	req_rw_in,
	req_byteen_in,
	req_addr_in,
	req_data_in,
	req_tag_in,
	req_ready_in,
	req_valid_out,
	req_rw_out,
	req_byteen_out,
	req_addr_out,
	req_data_out,
	req_tag_out,
	req_ready_out,
	rsp_valid_in,
	rsp_tmask_in,
	rsp_data_in,
	rsp_tag_in,
	rsp_ready_in,
	rsp_valid_out,
	rsp_tmask_out,
	rsp_data_out,
	rsp_tag_out,
	rsp_ready_out
);
	// Trace: ../../rtl/VX_smem_arb.sv:4:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/VX_smem_arb.sv:5:15
	parameter LANES = 1;
	// Trace: ../../rtl/VX_smem_arb.sv:6:15
	parameter DATA_SIZE = 1;
	// Trace: ../../rtl/VX_smem_arb.sv:7:15
	parameter TAG_IN_WIDTH = 1;
	// Trace: ../../rtl/VX_smem_arb.sv:8:15
	parameter TAG_SEL_IDX = 0;
	// Trace: ../../rtl/VX_smem_arb.sv:9:15
	parameter BUFFERED_REQ = 0;
	// Trace: ../../rtl/VX_smem_arb.sv:10:15
	parameter BUFFERED_RSP = 0;
	// Trace: ../../rtl/VX_smem_arb.sv:11:15
	parameter TYPE = "P";
	// Trace: ../../rtl/VX_smem_arb.sv:13:15
	parameter ADDR_WIDTH = 32 - $clog2(DATA_SIZE);
	// Trace: ../../rtl/VX_smem_arb.sv:14:15
	parameter DATA_WIDTH = 8 * DATA_SIZE;
	// Trace: ../../rtl/VX_smem_arb.sv:15:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: ../../rtl/VX_smem_arb.sv:16:15
	parameter TAG_OUT_WIDTH = TAG_IN_WIDTH - LOG_NUM_REQS;
	// Trace: ../../rtl/VX_smem_arb.sv:18:5
	input wire clk;
	// Trace: ../../rtl/VX_smem_arb.sv:19:5
	input wire reset;
	// Trace: ../../rtl/VX_smem_arb.sv:22:5
	input wire [LANES - 1:0] req_valid_in;
	// Trace: ../../rtl/VX_smem_arb.sv:23:5
	input wire [LANES - 1:0] req_rw_in;
	// Trace: ../../rtl/VX_smem_arb.sv:24:5
	input wire [(LANES * DATA_SIZE) - 1:0] req_byteen_in;
	// Trace: ../../rtl/VX_smem_arb.sv:25:5
	input wire [(LANES * ADDR_WIDTH) - 1:0] req_addr_in;
	// Trace: ../../rtl/VX_smem_arb.sv:26:5
	input wire [(LANES * DATA_WIDTH) - 1:0] req_data_in;
	// Trace: ../../rtl/VX_smem_arb.sv:27:5
	input wire [(LANES * TAG_IN_WIDTH) - 1:0] req_tag_in;
	// Trace: ../../rtl/VX_smem_arb.sv:28:5
	output wire [LANES - 1:0] req_ready_in;
	// Trace: ../../rtl/VX_smem_arb.sv:31:5
	output wire [(NUM_REQS * LANES) - 1:0] req_valid_out;
	// Trace: ../../rtl/VX_smem_arb.sv:32:5
	output wire [(NUM_REQS * LANES) - 1:0] req_rw_out;
	// Trace: ../../rtl/VX_smem_arb.sv:33:5
	output wire [((NUM_REQS * LANES) * DATA_SIZE) - 1:0] req_byteen_out;
	// Trace: ../../rtl/VX_smem_arb.sv:34:5
	output wire [((NUM_REQS * LANES) * ADDR_WIDTH) - 1:0] req_addr_out;
	// Trace: ../../rtl/VX_smem_arb.sv:35:5
	output wire [((NUM_REQS * LANES) * DATA_WIDTH) - 1:0] req_data_out;
	// Trace: ../../rtl/VX_smem_arb.sv:36:5
	output wire [((NUM_REQS * LANES) * TAG_OUT_WIDTH) - 1:0] req_tag_out;
	// Trace: ../../rtl/VX_smem_arb.sv:37:5
	input wire [(NUM_REQS * LANES) - 1:0] req_ready_out;
	// Trace: ../../rtl/VX_smem_arb.sv:40:5
	input wire [NUM_REQS - 1:0] rsp_valid_in;
	// Trace: ../../rtl/VX_smem_arb.sv:41:5
	input wire [(NUM_REQS * LANES) - 1:0] rsp_tmask_in;
	// Trace: ../../rtl/VX_smem_arb.sv:42:5
	input wire [((NUM_REQS * LANES) * DATA_WIDTH) - 1:0] rsp_data_in;
	// Trace: ../../rtl/VX_smem_arb.sv:43:5
	input wire [(NUM_REQS * TAG_OUT_WIDTH) - 1:0] rsp_tag_in;
	// Trace: ../../rtl/VX_smem_arb.sv:44:5
	output wire [NUM_REQS - 1:0] rsp_ready_in;
	// Trace: ../../rtl/VX_smem_arb.sv:47:5
	output wire rsp_valid_out;
	// Trace: ../../rtl/VX_smem_arb.sv:48:5
	output wire [LANES - 1:0] rsp_tmask_out;
	// Trace: ../../rtl/VX_smem_arb.sv:49:5
	output wire [(LANES * DATA_WIDTH) - 1:0] rsp_data_out;
	// Trace: ../../rtl/VX_smem_arb.sv:50:5
	output wire [TAG_IN_WIDTH - 1:0] rsp_tag_out;
	// Trace: ../../rtl/VX_smem_arb.sv:51:5
	input wire rsp_ready_out;
	// Trace: ../../rtl/VX_smem_arb.sv:53:5
	localparam REQ_DATAW = (((TAG_OUT_WIDTH + ADDR_WIDTH) + 1) + DATA_SIZE) + DATA_WIDTH;
	// Trace: ../../rtl/VX_smem_arb.sv:54:5
	localparam RSP_DATAW = (LANES * (1 + DATA_WIDTH)) + TAG_IN_WIDTH;
	// Trace: ../../rtl/VX_smem_arb.sv:56:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_REQS > 1) begin : genblk1
			// Trace: ../../rtl/VX_smem_arb.sv:58:9
			wire [(LANES * REQ_DATAW) - 1:0] req_data_in_merged;
			// Trace: ../../rtl/VX_smem_arb.sv:59:9
			wire [((NUM_REQS * LANES) * REQ_DATAW) - 1:0] req_data_out_merged;
			// Trace: ../../rtl/VX_smem_arb.sv:61:9
			wire [(LANES * LOG_NUM_REQS) - 1:0] req_sel;
			// Trace: ../../rtl/VX_smem_arb.sv:62:9
			wire [(LANES * TAG_OUT_WIDTH) - 1:0] req_tag_in_w;
			genvar i;
			for (i = 0; i < LANES; i = i + 1) begin : genblk1
				// Trace: ../../rtl/VX_smem_arb.sv:65:13
				assign req_sel[i * LOG_NUM_REQS+:LOG_NUM_REQS] = req_tag_in[(i * TAG_IN_WIDTH) + TAG_SEL_IDX+:LOG_NUM_REQS];
				// Trace: ../../rtl/VX_smem_arb.sv:67:13
				VX_bits_remove #(
					.N(TAG_IN_WIDTH),
					.S(LOG_NUM_REQS),
					.POS(TAG_SEL_IDX)
				) bits_remove(
					.data_in(req_tag_in[i * TAG_IN_WIDTH+:TAG_IN_WIDTH]),
					.data_out(req_tag_in_w[i * TAG_OUT_WIDTH+:TAG_OUT_WIDTH])
				);
				// Trace: ../../rtl/VX_smem_arb.sv:76:13
				assign req_data_in_merged[i * REQ_DATAW+:REQ_DATAW] = {req_tag_in_w[i * TAG_OUT_WIDTH+:TAG_OUT_WIDTH], req_addr_in[i * ADDR_WIDTH+:ADDR_WIDTH], req_rw_in[i], req_byteen_in[i * DATA_SIZE+:DATA_SIZE], req_data_in[i * DATA_WIDTH+:DATA_WIDTH]};
			end
			// Trace: ../../rtl/VX_smem_arb.sv:79:9
			VX_stream_demux #(
				.NUM_REQS(NUM_REQS),
				.LANES(LANES),
				.DATAW(REQ_DATAW),
				.BUFFERED(BUFFERED_REQ)
			) req_demux(
				.clk(clk),
				.reset(reset),
				.sel_in(req_sel),
				.valid_in(req_valid_in),
				.data_in(req_data_in_merged),
				.ready_in(req_ready_in),
				.valid_out(req_valid_out),
				.data_out(req_data_out_merged),
				.ready_out(req_ready_out)
			);
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk2
				genvar j;
				for (j = 0; j < LANES; j = j + 1) begin : genblk1
					// Trace: ../../rtl/VX_smem_arb.sv:98:17
					assign {req_tag_out[((i * LANES) + j) * TAG_OUT_WIDTH+:TAG_OUT_WIDTH], req_addr_out[((i * LANES) + j) * ADDR_WIDTH+:ADDR_WIDTH], req_rw_out[(i * LANES) + j], req_byteen_out[((i * LANES) + j) * DATA_SIZE+:DATA_SIZE], req_data_out[((i * LANES) + j) * DATA_WIDTH+:DATA_WIDTH]} = req_data_out_merged[((i * LANES) + j) * REQ_DATAW+:REQ_DATAW];
				end
			end
			// Trace: ../../rtl/VX_smem_arb.sv:104:9
			wire [(NUM_REQS * RSP_DATAW) - 1:0] rsp_data_in_merged;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk3
				// Trace: ../../rtl/VX_smem_arb.sv:107:13
				wire [TAG_IN_WIDTH - 1:0] rsp_tag_in_w;
				// Trace: ../../rtl/VX_smem_arb.sv:109:13
				VX_bits_insert #(
					.N(TAG_OUT_WIDTH),
					.S(LOG_NUM_REQS),
					.POS(TAG_SEL_IDX)
				) bits_insert(
					.data_in(rsp_tag_in[i * TAG_OUT_WIDTH+:TAG_OUT_WIDTH]),
					.sel_in(sv2v_cast_76B5F_signed(i)),
					.data_out(rsp_tag_in_w)
				);
				// Trace: ../../rtl/VX_smem_arb.sv:119:13
				assign rsp_data_in_merged[i * RSP_DATAW+:RSP_DATAW] = {rsp_tag_in_w, rsp_tmask_in[i * LANES+:LANES], rsp_data_in[DATA_WIDTH * (i * LANES)+:DATA_WIDTH * LANES]};
			end
			// Trace: ../../rtl/VX_smem_arb.sv:122:9
			VX_stream_arbiter #(
				.NUM_REQS(NUM_REQS),
				.LANES(1),
				.DATAW(RSP_DATAW),
				.BUFFERED(BUFFERED_RSP),
				.TYPE(TYPE)
			) rsp_arb(
				.clk(clk),
				.reset(reset),
				.valid_in(rsp_valid_in),
				.data_in(rsp_data_in_merged),
				.ready_in(rsp_ready_in),
				.valid_out(rsp_valid_out),
				.data_out({rsp_tag_out, rsp_tmask_out, rsp_data_out}),
				.ready_out(rsp_ready_out)
			);
		end
		else begin : genblk1
			// Trace: ../../rtl/VX_smem_arb.sv:144:9
			assign req_valid_out = req_valid_in;
			// Trace: ../../rtl/VX_smem_arb.sv:145:9
			assign req_tag_out = req_tag_in;
			// Trace: ../../rtl/VX_smem_arb.sv:146:9
			assign req_addr_out = req_addr_in;
			// Trace: ../../rtl/VX_smem_arb.sv:147:9
			assign req_rw_out = req_rw_in;
			// Trace: ../../rtl/VX_smem_arb.sv:148:9
			assign req_byteen_out = req_byteen_in;
			// Trace: ../../rtl/VX_smem_arb.sv:149:9
			assign req_data_out = req_data_in;
			// Trace: ../../rtl/VX_smem_arb.sv:150:9
			assign req_ready_in = req_ready_out;
			// Trace: ../../rtl/VX_smem_arb.sv:152:9
			assign rsp_valid_out = rsp_valid_in;
			// Trace: ../../rtl/VX_smem_arb.sv:153:9
			assign rsp_tmask_out = rsp_tmask_in;
			// Trace: ../../rtl/VX_smem_arb.sv:154:9
			assign rsp_tag_out = rsp_tag_in;
			// Trace: ../../rtl/VX_smem_arb.sv:155:9
			assign rsp_data_out = rsp_data_in;
			// Trace: ../../rtl/VX_smem_arb.sv:156:9
			assign rsp_ready_in = rsp_ready_out;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_warp_sched
// removed module with interface ports: VX_writeback
module Vortex (
	clk,
	reset,
	mem_req_valid,
	mem_req_rw,
	mem_req_byteen,
	mem_req_addr,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready,
	busy
);
	// Trace: ../../rtl/Vortex.sv:7:5
	input wire clk;
	// Trace: ../../rtl/Vortex.sv:8:5
	input wire reset;
	// Trace: ../../rtl/Vortex.sv:11:5
	output wire mem_req_valid;
	// Trace: ../../rtl/Vortex.sv:12:5
	output wire mem_req_rw;
	// Trace: ../../rtl/Vortex.sv:13:5
	output wire [(0 || 0 ? 16 : 64) - 1:0] mem_req_byteen;
	// Trace: ../../rtl/Vortex.sv:14:5
	output wire [(32 - $clog2((0 || 0 ? 16 : 64))) - 1:0] mem_req_addr;
	// Trace: ../../rtl/Vortex.sv:15:5
	output wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_req_data;
	// Trace: ../../rtl/Vortex.sv:16:5
	output wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_req_tag;
	// Trace: ../../rtl/Vortex.sv:17:5
	input wire mem_req_ready;
	// Trace: ../../rtl/Vortex.sv:20:5
	input wire mem_rsp_valid;
	// Trace: ../../rtl/Vortex.sv:21:5
	input wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_rsp_data;
	// Trace: ../../rtl/Vortex.sv:22:5
	input wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_rsp_tag;
	// Trace: ../../rtl/Vortex.sv:23:5
	output wire mem_rsp_ready;
	// Trace: ../../rtl/Vortex.sv:26:5
	output wire busy;
	// Trace: ../../rtl/Vortex.sv:30:5
	wire [0:0] per_cluster_mem_req_valid;
	// Trace: ../../rtl/Vortex.sv:31:5
	wire [0:0] per_cluster_mem_req_rw;
	// Trace: ../../rtl/Vortex.sv:32:5
	wire [(0 || 0 ? 16 : 64) - 1:0] per_cluster_mem_req_byteen;
	// Trace: ../../rtl/Vortex.sv:33:5
	wire [(32 - $clog2((0 || 0 ? 16 : 64))) - 1:0] per_cluster_mem_req_addr;
	// Trace: ../../rtl/Vortex.sv:34:5
	wire [((0 || 0 ? 16 : 64) * 8) - 1:0] per_cluster_mem_req_data;
	// Trace: ../../rtl/Vortex.sv:35:5
	wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] per_cluster_mem_req_tag;
	// Trace: ../../rtl/Vortex.sv:36:5
	wire [0:0] per_cluster_mem_req_ready;
	// Trace: ../../rtl/Vortex.sv:38:5
	wire [0:0] per_cluster_mem_rsp_valid;
	// Trace: ../../rtl/Vortex.sv:39:5
	wire [((0 || 0 ? 16 : 64) * 8) - 1:0] per_cluster_mem_rsp_data;
	// Trace: ../../rtl/Vortex.sv:40:5
	wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] per_cluster_mem_rsp_tag;
	// Trace: ../../rtl/Vortex.sv:41:5
	wire [0:0] per_cluster_mem_rsp_ready;
	// Trace: ../../rtl/Vortex.sv:43:5
	wire [0:0] per_cluster_busy;
	// Trace: ../../rtl/Vortex.sv:45:5
	genvar i;
	generate
		for (i = 0; i < 1; i = i + 1) begin : genblk1
			// Trace: macro expansion of RESET_RELAY at ../../rtl/Vortex.sv:47:30
			wire cluster_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/Vortex.sv:47:63
			VX_reset_relay __cluster_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(cluster_reset)
			);
			// Trace: ../../rtl/Vortex.sv:49:9
			VX_cluster #(.CLUSTER_ID(i)) cluster(
				.clk(clk),
				.reset(cluster_reset),
				.mem_req_valid(per_cluster_mem_req_valid[i]),
				.mem_req_rw(per_cluster_mem_req_rw[i]),
				.mem_req_byteen(per_cluster_mem_req_byteen[i * (0 || 0 ? 16 : 64)+:(0 || 0 ? 16 : 64)]),
				.mem_req_addr(per_cluster_mem_req_addr[i * (32 - $clog2((0 || 0 ? 16 : 64)))+:32 - $clog2((0 || 0 ? 16 : 64))]),
				.mem_req_data(per_cluster_mem_req_data[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8]),
				.mem_req_tag(per_cluster_mem_req_tag[i * ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1)+:(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1]),
				.mem_req_ready(per_cluster_mem_req_ready[i]),
				.mem_rsp_valid(per_cluster_mem_rsp_valid[i]),
				.mem_rsp_data(per_cluster_mem_rsp_data[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8]),
				.mem_rsp_tag(per_cluster_mem_rsp_tag[i * ((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1)+:(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1]),
				.mem_rsp_ready(per_cluster_mem_rsp_ready[i]),
				.busy(per_cluster_busy[i])
			);
		end
	endgenerate
	// Trace: ../../rtl/Vortex.sv:74:5
	assign busy = |per_cluster_busy;
	// Trace: ../../rtl/Vortex.sv:76:5
	generate
		if (1) begin : genblk2
			// Trace: macro expansion of RESET_RELAY at ../../rtl/Vortex.sv:145:30
			wire mem_arb_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/Vortex.sv:145:63
			VX_reset_relay __mem_arb_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(mem_arb_reset)
			);
			// Trace: ../../rtl/Vortex.sv:147:9
			VX_mem_arb #(
				.NUM_REQS(1),
				.DATA_WIDTH((0 || 0 ? 16 : 64) * 8),
				.ADDR_WIDTH(32 - $clog2((0 || 0 ? 16 : 64))),
				.TAG_IN_WIDTH((1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 1),
				.TYPE("R"),
				.BUFFERED_REQ(1),
				.BUFFERED_RSP(1)
			) mem_arb(
				.clk(clk),
				.reset(mem_arb_reset),
				.req_valid_in(per_cluster_mem_req_valid),
				.req_rw_in(per_cluster_mem_req_rw),
				.req_byteen_in(per_cluster_mem_req_byteen),
				.req_addr_in(per_cluster_mem_req_addr),
				.req_data_in(per_cluster_mem_req_data),
				.req_tag_in(per_cluster_mem_req_tag),
				.req_ready_in(per_cluster_mem_req_ready),
				.req_valid_out(mem_req_valid),
				.req_rw_out(mem_req_rw),
				.req_byteen_out(mem_req_byteen),
				.req_addr_out(mem_req_addr),
				.req_data_out(mem_req_data),
				.req_tag_out(mem_req_tag),
				.req_ready_out(mem_req_ready),
				.rsp_valid_out(per_cluster_mem_rsp_valid),
				.rsp_data_out(per_cluster_mem_rsp_data),
				.rsp_tag_out(per_cluster_mem_rsp_tag),
				.rsp_ready_out(per_cluster_mem_rsp_ready),
				.rsp_valid_in(mem_rsp_valid),
				.rsp_tag_in(mem_rsp_tag),
				.rsp_data_in(mem_rsp_data),
				.rsp_ready_in(mem_rsp_ready)
			);
		end
	endgenerate
endmodule


module local_mem (
	clk,
	reset,
	mem_req_valid,
	mem_req_rw,
	mem_req_byteen,
	mem_req_addr,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready,
	busy,
	tb_addr_out_of_bounds
);
	// Trace: ../../rtl/local_mem.sv:16:5
	input clk;
	input reset;
	// Trace: ../../rtl/local_mem.sv:20:5
	input wire mem_req_valid;
	// Trace: ../../rtl/local_mem.sv:21:5
	input wire mem_req_rw;
	// Trace: ../../rtl/local_mem.sv:22:5
	input wire [(0 || 0 ? 16 : 64) - 1:0] mem_req_byteen;
	// Trace: ../../rtl/local_mem.sv:23:5
	input wire [(32 - $clog2((0 || 0 ? 16 : 64))) - 1:0] mem_req_addr;
	// Trace: ../../rtl/local_mem.sv:24:5
	input wire [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_req_data;
	// Trace: ../../rtl/local_mem.sv:25:5
	input wire [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_req_tag;
	// Trace: ../../rtl/local_mem.sv:27:5
	output reg mem_req_ready;
	// Trace: ../../rtl/local_mem.sv:31:5
	output reg mem_rsp_valid;
	// Trace: ../../rtl/local_mem.sv:32:5
	output reg [((0 || 0 ? 16 : 64) * 8) - 1:0] mem_rsp_data;
	// Trace: ../../rtl/local_mem.sv:33:5
	output reg [(1 > (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 1 : (4 > ((1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48) ? 4 : (1 + $clog2((0 || 0 ? 16 : 64) / 4)) + 48)) + 0:0] mem_rsp_tag;
	// Trace: ../../rtl/local_mem.sv:35:5
	input wire mem_rsp_ready;
	// Trace: ../../rtl/local_mem.sv:39:5
	input wire busy;
	// Trace: ../../rtl/local_mem.sv:42:5
	output reg tb_addr_out_of_bounds;
	// Trace: ../../rtl/local_mem.sv:47:5
	reg wen_0_80000000;
	// Trace: ../../rtl/local_mem.sv:48:5
	reg [5:0] wsel_0_80000000;
	// Trace: ../../rtl/local_mem.sv:49:5
	reg [((0 || 0 ? 16 : 64) * 8) - 1:0] wdata_0_80000000;
	// Trace: ../../rtl/local_mem.sv:50:5
	reg [5:0] rsel_0_80000000;
	// Trace: ../../rtl/local_mem.sv:51:5
	reg [((0 || 0 ? 16 : 64) * 8) - 1:0] rdata_0_80000000;
	// Trace: ../../rtl/local_mem.sv:53:5
	reg [(64 * ((0 || 0 ? 16 : 64) * 8)) - 1:0] reg_val_0_80000000;
	// Trace: ../../rtl/local_mem.sv:54:5
	reg [(64 * ((0 || 0 ? 16 : 64) * 8)) - 1:0] next_reg_val_0_80000000;
	// Trace: ../../rtl/local_mem.sv:56:5
	always @(posedge clk) begin : REGISTER_LOGIC_0_80000000
		// Trace: ../../rtl/local_mem.sv:57:9
		if (reset) begin
			// Trace: ../../rtl/local_mem.sv:60:13
			reg_val_0_80000000[31-:32] <= 32'hfc102573;
			// Trace: ../../rtl/local_mem.sv:61:13
			reg_val_0_80000000[63-:32] <= 32'h00000597;
			// Trace: ../../rtl/local_mem.sv:62:13
			reg_val_0_80000000[95-:32] <= 32'h09c58593;
			// Trace: ../../rtl/local_mem.sv:63:13
			reg_val_0_80000000[127-:32] <= 32'h00b5106b;
			// Trace: ../../rtl/local_mem.sv:64:13
			reg_val_0_80000000[159-:32] <= 32'h090000ef;
			// Trace: ../../rtl/local_mem.sv:65:13
			reg_val_0_80000000[191-:32] <= 32'h00100513;
			// Trace: ../../rtl/local_mem.sv:66:13
			reg_val_0_80000000[223-:32] <= 32'h0005006b;
			// Trace: ../../rtl/local_mem.sv:67:13
			reg_val_0_80000000[255-:32] <= 32'hfc102573;
			// Trace: ../../rtl/local_mem.sv:68:13
			reg_val_0_80000000[287-:32] <= 32'h00000597;
			// Trace: ../../rtl/local_mem.sv:69:13
			reg_val_0_80000000[319-:32] <= 32'h12058593;
			// Trace: ../../rtl/local_mem.sv:70:13
			reg_val_0_80000000[351-:32] <= 32'h00b5106b;
			// Trace: ../../rtl/local_mem.sv:71:13
			reg_val_0_80000000[383-:32] <= 32'h114000ef;
			// Trace: ../../rtl/local_mem.sv:72:13
			reg_val_0_80000000[415-:32] <= 32'h00100513;
			// Trace: ../../rtl/local_mem.sv:73:13
			reg_val_0_80000000[447-:32] <= 32'h0005006b;
			// Trace: ../../rtl/local_mem.sv:74:13
			reg_val_0_80000000[479-:32] <= 32'h00001517;
			// Trace: ../../rtl/local_mem.sv:75:13
			reg_val_0_80000000[511-:32] <= 32'h40850513;
			// Trace: ../../rtl/local_mem.sv:76:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 31-:32] <= 32'h00001617;
			// Trace: ../../rtl/local_mem.sv:77:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 63-:32] <= 32'h48060613;
			// Trace: ../../rtl/local_mem.sv:78:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 95-:32] <= 32'h40a60633;
			// Trace: ../../rtl/local_mem.sv:79:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 127-:32] <= 32'h00000593;
			// Trace: ../../rtl/local_mem.sv:80:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 159-:32] <= 32'h29d000ef;
			// Trace: ../../rtl/local_mem.sv:81:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 191-:32] <= 32'h00000517;
			// Trace: ../../rtl/local_mem.sv:82:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 223-:32] <= 32'h1dc50513;
			// Trace: ../../rtl/local_mem.sv:83:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 255-:32] <= 32'h12d000ef;
			// Trace: ../../rtl/local_mem.sv:84:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 287-:32] <= 32'h13c000ef;
			// Trace: ../../rtl/local_mem.sv:85:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 319-:32] <= 32'h008000ef;
			// Trace: ../../rtl/local_mem.sv:86:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 351-:32] <= 32'h1350006f;
			// Trace: ../../rtl/local_mem.sv:87:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 383-:32] <= 32'hfff00793;
			// Trace: ../../rtl/local_mem.sv:88:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 415-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:89:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 447-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:90:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 479-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:91:13
			reg_val_0_80000000[((0 || 0 ? 16 : 64) * 8) + 511-:32] <= 32'h00000793;
			// Trace: ../../rtl/local_mem.sv:92:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00078863;
			// Trace: ../../rtl/local_mem.sv:93:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h80000537;
			// Trace: ../../rtl/local_mem.sv:94:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h23050513;
			// Trace: ../../rtl/local_mem.sv:95:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h0fd0006f;
			// Trace: ../../rtl/local_mem.sv:96:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:97:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00040193;
			// Trace: ../../rtl/local_mem.sv:98:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:99:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h0005006b;
			// Trace: ../../rtl/local_mem.sv:100:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:101:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h0005006b;
			// Trace: ../../rtl/local_mem.sv:102:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00001197;
			// Trace: ../../rtl/local_mem.sv:103:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h76018193;
			// Trace: ../../rtl/local_mem.sv:104:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hff000137;
			// Trace: ../../rtl/local_mem.sv:105:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hcc102573;
			// Trace: ../../rtl/local_mem.sv:106:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00a51593;
			// Trace: ../../rtl/local_mem.sv:107:13
			reg_val_0_80000000[(2 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h40b10133;
			// Trace: ../../rtl/local_mem.sv:108:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000593;
			// Trace: ../../rtl/local_mem.sv:109:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h02b50533;
			// Trace: ../../rtl/local_mem.sv:110:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00001217;
			// Trace: ../../rtl/local_mem.sv:111:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h43720213;
			// Trace: ../../rtl/local_mem.sv:112:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00a20233;
			// Trace: ../../rtl/local_mem.sv:113:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hfc027213;
			// Trace: ../../rtl/local_mem.sv:114:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hcc3026f3;
			// Trace: ../../rtl/local_mem.sv:115:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00068663;
			// Trace: ../../rtl/local_mem.sv:116:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:117:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h0005006b;
			// Trace: ../../rtl/local_mem.sv:118:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:119:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:120:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:121:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:122:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:123:13
			reg_val_0_80000000[(3 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:124:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:125:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:126:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:127:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:128:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:129:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:130:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:131:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00100073;
			// Trace: ../../rtl/local_mem.sv:132:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:133:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:134:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00060513;
			// Trace: ../../rtl/local_mem.sv:135:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:136:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:137:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:138:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hf1402573;
			// Trace: ../../rtl/local_mem.sv:139:13
			reg_val_0_80000000[(4 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:140:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hff010113;
			// Trace: ../../rtl/local_mem.sv:141:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00112623;
			// Trace: ../../rtl/local_mem.sv:142:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00812423;
			// Trace: ../../rtl/local_mem.sv:143:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hfff00793;
			// Trace: ../../rtl/local_mem.sv:144:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:145:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000613;
			// Trace: ../../rtl/local_mem.sv:146:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00020513;
			// Trace: ../../rtl/local_mem.sv:147:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00001597;
			// Trace: ../../rtl/local_mem.sv:148:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hea458593;
			// Trace: ../../rtl/local_mem.sv:149:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00020413;
			// Trace: ../../rtl/local_mem.sv:150:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h069000ef;
			// Trace: ../../rtl/local_mem.sv:151:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:152:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000613;
			// Trace: ../../rtl/local_mem.sv:153:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000593;
			// Trace: ../../rtl/local_mem.sv:154:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00a40533;
			// Trace: ../../rtl/local_mem.sv:155:13
			reg_val_0_80000000[(5 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h171000ef;
			// Trace: ../../rtl/local_mem.sv:156:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hcc3027f3;
			// Trace: ../../rtl/local_mem.sv:157:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h0017b793;
			// Trace: ../../rtl/local_mem.sv:158:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:159:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00c12083;
			// Trace: ../../rtl/local_mem.sv:160:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00812403;
			// Trace: ../../rtl/local_mem.sv:161:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h01010113;
			// Trace: ../../rtl/local_mem.sv:162:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:163:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hff010113;
			// Trace: ../../rtl/local_mem.sv:164:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00812423;
			// Trace: ../../rtl/local_mem.sv:165:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h01212023;
			// Trace: ../../rtl/local_mem.sv:166:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00001417;
			// Trace: ../../rtl/local_mem.sv:167:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'he5840413;
			// Trace: ../../rtl/local_mem.sv:168:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00001917;
			// Trace: ../../rtl/local_mem.sv:169:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'he5090913;
			// Trace: ../../rtl/local_mem.sv:170:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h40890933;
			// Trace: ../../rtl/local_mem.sv:171:13
			reg_val_0_80000000[(6 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00112623;
			// Trace: ../../rtl/local_mem.sv:172:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00912223;
			// Trace: ../../rtl/local_mem.sv:173:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h40295913;
			// Trace: ../../rtl/local_mem.sv:174:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00090e63;
			// Trace: ../../rtl/local_mem.sv:175:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000493;
			// Trace: ../../rtl/local_mem.sv:176:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00042783;
			// Trace: ../../rtl/local_mem.sv:177:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00148493;
			// Trace: ../../rtl/local_mem.sv:178:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00440413;
			// Trace: ../../rtl/local_mem.sv:179:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h000780e7;
			// Trace: ../../rtl/local_mem.sv:180:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hfe9918e3;
			// Trace: ../../rtl/local_mem.sv:181:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00001417;
			// Trace: ../../rtl/local_mem.sv:182:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'he1c40413;
			// Trace: ../../rtl/local_mem.sv:183:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00001917;
			// Trace: ../../rtl/local_mem.sv:184:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'he1890913;
			// Trace: ../../rtl/local_mem.sv:185:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h40890933;
			// Trace: ../../rtl/local_mem.sv:186:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h40295913;
			// Trace: ../../rtl/local_mem.sv:187:13
			reg_val_0_80000000[(7 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00090e63;
			// Trace: ../../rtl/local_mem.sv:188:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000493;
			// Trace: ../../rtl/local_mem.sv:189:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00042783;
			// Trace: ../../rtl/local_mem.sv:190:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00148493;
			// Trace: ../../rtl/local_mem.sv:191:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00440413;
			// Trace: ../../rtl/local_mem.sv:192:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h000780e7;
			// Trace: ../../rtl/local_mem.sv:193:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hfe9918e3;
			// Trace: ../../rtl/local_mem.sv:194:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00c12083;
			// Trace: ../../rtl/local_mem.sv:195:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00812403;
			// Trace: ../../rtl/local_mem.sv:196:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00412483;
			// Trace: ../../rtl/local_mem.sv:197:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00012903;
			// Trace: ../../rtl/local_mem.sv:198:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h01010113;
			// Trace: ../../rtl/local_mem.sv:199:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:200:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hff010113;
			// Trace: ../../rtl/local_mem.sv:201:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00812423;
			// Trace: ../../rtl/local_mem.sv:202:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00001797;
			// Trace: ../../rtl/local_mem.sv:203:13
			reg_val_0_80000000[(8 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'hdcc78793;
			// Trace: ../../rtl/local_mem.sv:204:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00001417;
			// Trace: ../../rtl/local_mem.sv:205:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hdc440413;
			// Trace: ../../rtl/local_mem.sv:206:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h408787b3;
			// Trace: ../../rtl/local_mem.sv:207:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00912223;
			// Trace: ../../rtl/local_mem.sv:208:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00112623;
			// Trace: ../../rtl/local_mem.sv:209:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h4027d493;
			// Trace: ../../rtl/local_mem.sv:210:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h02048063;
			// Trace: ../../rtl/local_mem.sv:211:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hffc78793;
			// Trace: ../../rtl/local_mem.sv:212:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00878433;
			// Trace: ../../rtl/local_mem.sv:213:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00042783;
			// Trace: ../../rtl/local_mem.sv:214:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hfff48493;
			// Trace: ../../rtl/local_mem.sv:215:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hffc40413;
			// Trace: ../../rtl/local_mem.sv:216:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h000780e7;
			// Trace: ../../rtl/local_mem.sv:217:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hfe0498e3;
			// Trace: ../../rtl/local_mem.sv:218:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00c12083;
			// Trace: ../../rtl/local_mem.sv:219:13
			reg_val_0_80000000[(9 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00812403;
			// Trace: ../../rtl/local_mem.sv:220:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00412483;
			// Trace: ../../rtl/local_mem.sv:221:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h01010113;
			// Trace: ../../rtl/local_mem.sv:222:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:223:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hff010113;
			// Trace: ../../rtl/local_mem.sv:224:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00112623;
			// Trace: ../../rtl/local_mem.sv:225:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00812423;
			// Trace: ../../rtl/local_mem.sv:226:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00912223;
			// Trace: ../../rtl/local_mem.sv:227:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h01212023;
			// Trace: ../../rtl/local_mem.sv:228:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hcc5027f3;
			// Trace: ../../rtl/local_mem.sv:229:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'hcc302773;
			// Trace: ../../rtl/local_mem.sv:230:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hcc0026f3;
			// Trace: ../../rtl/local_mem.sv:231:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hfc0025f3;
			// Trace: ../../rtl/local_mem.sv:232:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00279613;
			// Trace: ../../rtl/local_mem.sv:233:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00001797;
			// Trace: ../../rtl/local_mem.sv:234:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h18c78793;
			// Trace: ../../rtl/local_mem.sv:235:13
			reg_val_0_80000000[(10 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00c787b3;
			// Trace: ../../rtl/local_mem.sv:236:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h0007a483;
			// Trace: ../../rtl/local_mem.sv:237:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h0104a403;
			// Trace: ../../rtl/local_mem.sv:238:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00c4a603;
			// Trace: ../../rtl/local_mem.sv:239:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00872933;
			// Trace: ../../rtl/local_mem.sv:240:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00040793;
			// Trace: ../../rtl/local_mem.sv:241:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00c90933;
			// Trace: ../../rtl/local_mem.sv:242:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h02e60433;
			// Trace: ../../rtl/local_mem.sv:243:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00f75463;
			// Trace: ../../rtl/local_mem.sv:244:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00070793;
			// Trace: ../../rtl/local_mem.sv:245:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00f40433;
			// Trace: ../../rtl/local_mem.sv:246:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h0084a703;
			// Trace: ../../rtl/local_mem.sv:247:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h02b40433;
			// Trace: ../../rtl/local_mem.sv:248:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h02d907b3;
			// Trace: ../../rtl/local_mem.sv:249:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00e40433;
			// Trace: ../../rtl/local_mem.sv:250:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00f40433;
			// Trace: ../../rtl/local_mem.sv:251:13
			reg_val_0_80000000[(11 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00890933;
			// Trace: ../../rtl/local_mem.sv:252:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h01245e63;
			// Trace: ../../rtl/local_mem.sv:253:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h0004a783;
			// Trace: ../../rtl/local_mem.sv:254:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h0044a583;
			// Trace: ../../rtl/local_mem.sv:255:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00040513;
			// Trace: ../../rtl/local_mem.sv:256:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00140413;
			// Trace: ../../rtl/local_mem.sv:257:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h000780e7;
			// Trace: ../../rtl/local_mem.sv:258:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hfe8916e3;
			// Trace: ../../rtl/local_mem.sv:259:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h0144a703;
			// Trace: ../../rtl/local_mem.sv:260:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000793;
			// Trace: ../../rtl/local_mem.sv:261:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00e7c06b;
			// Trace: ../../rtl/local_mem.sv:262:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00c12083;
			// Trace: ../../rtl/local_mem.sv:263:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00812403;
			// Trace: ../../rtl/local_mem.sv:264:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00412483;
			// Trace: ../../rtl/local_mem.sv:265:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00012903;
			// Trace: ../../rtl/local_mem.sv:266:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h01010113;
			// Trace: ../../rtl/local_mem.sv:267:13
			reg_val_0_80000000[(12 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:268:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hcc5027f3;
			// Trace: ../../rtl/local_mem.sv:269:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hcc202573;
			// Trace: ../../rtl/local_mem.sv:270:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00279713;
			// Trace: ../../rtl/local_mem.sv:271:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00001797;
			// Trace: ../../rtl/local_mem.sv:272:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h0f478793;
			// Trace: ../../rtl/local_mem.sv:273:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00e787b3;
			// Trace: ../../rtl/local_mem.sv:274:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h0007a783;
			// Trace: ../../rtl/local_mem.sv:275:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h0087a703;
			// Trace: ../../rtl/local_mem.sv:276:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h0007a303;
			// Trace: ../../rtl/local_mem.sv:277:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h0047a583;
			// Trace: ../../rtl/local_mem.sv:278:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00e50533;
			// Trace: ../../rtl/local_mem.sv:279:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00030067;
			// Trace: ../../rtl/local_mem.sv:280:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hff010113;
			// Trace: ../../rtl/local_mem.sv:281:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00112623;
			// Trace: ../../rtl/local_mem.sv:282:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hfff00793;
			// Trace: ../../rtl/local_mem.sv:283:13
			reg_val_0_80000000[(13 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:284:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hf0dff0ef;
			// Trace: ../../rtl/local_mem.sv:285:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hcc3027f3;
			// Trace: ../../rtl/local_mem.sv:286:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h0017b793;
			// Trace: ../../rtl/local_mem.sv:287:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:288:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00c12083;
			// Trace: ../../rtl/local_mem.sv:289:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h01010113;
			// Trace: ../../rtl/local_mem.sv:290:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:291:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hfe010113;
			// Trace: ../../rtl/local_mem.sv:292:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00112e23;
			// Trace: ../../rtl/local_mem.sv:293:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00812c23;
			// Trace: ../../rtl/local_mem.sv:294:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00912a23;
			// Trace: ../../rtl/local_mem.sv:295:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01212823;
			// Trace: ../../rtl/local_mem.sv:296:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h01312623;
			// Trace: ../../rtl/local_mem.sv:297:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h01412423;
			// Trace: ../../rtl/local_mem.sv:298:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hcc5027f3;
			// Trace: ../../rtl/local_mem.sv:299:13
			reg_val_0_80000000[(14 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'hcc302773;
			// Trace: ../../rtl/local_mem.sv:300:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hcc0026f3;
			// Trace: ../../rtl/local_mem.sv:301:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hfc002573;
			// Trace: ../../rtl/local_mem.sv:302:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00279613;
			// Trace: ../../rtl/local_mem.sv:303:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00001797;
			// Trace: ../../rtl/local_mem.sv:304:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h07478793;
			// Trace: ../../rtl/local_mem.sv:305:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00c787b3;
			// Trace: ../../rtl/local_mem.sv:306:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h0007a403;
			// Trace: ../../rtl/local_mem.sv:307:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h01442483;
			// Trace: ../../rtl/local_mem.sv:308:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h01042603;
			// Trace: ../../rtl/local_mem.sv:309:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00972a33;
			// Trace: ../../rtl/local_mem.sv:310:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00048793;
			// Trace: ../../rtl/local_mem.sv:311:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00ca0a33;
			// Trace: ../../rtl/local_mem.sv:312:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h02e604b3;
			// Trace: ../../rtl/local_mem.sv:313:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00f75463;
			// Trace: ../../rtl/local_mem.sv:314:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00070793;
			// Trace: ../../rtl/local_mem.sv:315:13
			reg_val_0_80000000[(15 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00f484b3;
			// Trace: ../../rtl/local_mem.sv:316:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00042583;
			// Trace: ../../rtl/local_mem.sv:317:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00c42703;
			// Trace: ../../rtl/local_mem.sv:318:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h0005a903;
			// Trace: ../../rtl/local_mem.sv:319:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h0045a983;
			// Trace: ../../rtl/local_mem.sv:320:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h02a484b3;
			// Trace: ../../rtl/local_mem.sv:321:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h02da07b3;
			// Trace: ../../rtl/local_mem.sv:322:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00e484b3;
			// Trace: ../../rtl/local_mem.sv:323:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00f484b3;
			// Trace: ../../rtl/local_mem.sv:324:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h009a0a33;
			// Trace: ../../rtl/local_mem.sv:325:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h033909b3;
			// Trace: ../../rtl/local_mem.sv:326:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h0744c063;
			// Trace: ../../rtl/local_mem.sv:327:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h0800006f;
			// Trace: ../../rtl/local_mem.sv:328:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h01e44703;
			// Trace: ../../rtl/local_mem.sv:329:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h01d44683;
			// Trace: ../../rtl/local_mem.sv:330:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h40e4d733;
			// Trace: ../../rtl/local_mem.sv:331:13
			reg_val_0_80000000[(16 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h033707b3;
			// Trace: ../../rtl/local_mem.sv:332:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h40f487b3;
			// Trace: ../../rtl/local_mem.sv:333:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h06068063;
			// Trace: ../../rtl/local_mem.sv:334:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h01f44683;
			// Trace: ../../rtl/local_mem.sv:335:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h40d7d6b3;
			// Trace: ../../rtl/local_mem.sv:336:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h032688b3;
			// Trace: ../../rtl/local_mem.sv:337:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h0145ae03;
			// Trace: ../../rtl/local_mem.sv:338:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h0105a303;
			// Trace: ../../rtl/local_mem.sv:339:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00c5a603;
			// Trace: ../../rtl/local_mem.sv:340:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00442803;
			// Trace: ../../rtl/local_mem.sv:341:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00842503;
			// Trace: ../../rtl/local_mem.sv:342:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00148493;
			// Trace: ../../rtl/local_mem.sv:343:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01c70733;
			// Trace: ../../rtl/local_mem.sv:344:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h006686b3;
			// Trace: ../../rtl/local_mem.sv:345:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h411787b3;
			// Trace: ../../rtl/local_mem.sv:346:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00c78633;
			// Trace: ../../rtl/local_mem.sv:347:13
			reg_val_0_80000000[(17 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h000800e7;
			// Trace: ../../rtl/local_mem.sv:348:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h029a0663;
			// Trace: ../../rtl/local_mem.sv:349:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00042583;
			// Trace: ../../rtl/local_mem.sv:350:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h01c44783;
			// Trace: ../../rtl/local_mem.sv:351:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hfa0792e3;
			// Trace: ../../rtl/local_mem.sv:352:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h0334c733;
			// Trace: ../../rtl/local_mem.sv:353:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h01d44683;
			// Trace: ../../rtl/local_mem.sv:354:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h033707b3;
			// Trace: ../../rtl/local_mem.sv:355:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h40f487b3;
			// Trace: ../../rtl/local_mem.sv:356:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hfa0694e3;
			// Trace: ../../rtl/local_mem.sv:357:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h0327c6b3;
			// Trace: ../../rtl/local_mem.sv:358:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hfa9ff06f;
			// Trace: ../../rtl/local_mem.sv:359:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01842703;
			// Trace: ../../rtl/local_mem.sv:360:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000793;
			// Trace: ../../rtl/local_mem.sv:361:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00e7c06b;
			// Trace: ../../rtl/local_mem.sv:362:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h01c12083;
			// Trace: ../../rtl/local_mem.sv:363:13
			reg_val_0_80000000[(18 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h01812403;
			// Trace: ../../rtl/local_mem.sv:364:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h01412483;
			// Trace: ../../rtl/local_mem.sv:365:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h01012903;
			// Trace: ../../rtl/local_mem.sv:366:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00c12983;
			// Trace: ../../rtl/local_mem.sv:367:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00812a03;
			// Trace: ../../rtl/local_mem.sv:368:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h02010113;
			// Trace: ../../rtl/local_mem.sv:369:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:370:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hcc502773;
			// Trace: ../../rtl/local_mem.sv:371:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hcc2027f3;
			// Trace: ../../rtl/local_mem.sv:372:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00271693;
			// Trace: ../../rtl/local_mem.sv:373:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00001717;
			// Trace: ../../rtl/local_mem.sv:374:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hf5c70713;
			// Trace: ../../rtl/local_mem.sv:375:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00d70733;
			// Trace: ../../rtl/local_mem.sv:376:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00072503;
			// Trace: ../../rtl/local_mem.sv:377:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00052583;
			// Trace: ../../rtl/local_mem.sv:378:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00c52683;
			// Trace: ../../rtl/local_mem.sv:379:13
			reg_val_0_80000000[(19 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h01c54703;
			// Trace: ../../rtl/local_mem.sv:380:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h0005a883;
			// Trace: ../../rtl/local_mem.sv:381:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h0045a603;
			// Trace: ../../rtl/local_mem.sv:382:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00d787b3;
			// Trace: ../../rtl/local_mem.sv:383:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h02c88633;
			// Trace: ../../rtl/local_mem.sv:384:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h04070863;
			// Trace: ../../rtl/local_mem.sv:385:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h01e54703;
			// Trace: ../../rtl/local_mem.sv:386:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h01d54683;
			// Trace: ../../rtl/local_mem.sv:387:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h40e7d733;
			// Trace: ../../rtl/local_mem.sv:388:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h02c70633;
			// Trace: ../../rtl/local_mem.sv:389:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h40c787b3;
			// Trace: ../../rtl/local_mem.sv:390:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h04068663;
			// Trace: ../../rtl/local_mem.sv:391:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01f54683;
			// Trace: ../../rtl/local_mem.sv:392:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h40d7d833;
			// Trace: ../../rtl/local_mem.sv:393:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h0105a683;
			// Trace: ../../rtl/local_mem.sv:394:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h0145ae03;
			// Trace: ../../rtl/local_mem.sv:395:13
			reg_val_0_80000000[(20 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00c5a603;
			// Trace: ../../rtl/local_mem.sv:396:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00d806b3;
			// Trace: ../../rtl/local_mem.sv:397:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h03180833;
			// Trace: ../../rtl/local_mem.sv:398:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00452303;
			// Trace: ../../rtl/local_mem.sv:399:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00852503;
			// Trace: ../../rtl/local_mem.sv:400:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h01c70733;
			// Trace: ../../rtl/local_mem.sv:401:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h410787b3;
			// Trace: ../../rtl/local_mem.sv:402:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00c78633;
			// Trace: ../../rtl/local_mem.sv:403:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00030067;
			// Trace: ../../rtl/local_mem.sv:404:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h02c7c733;
			// Trace: ../../rtl/local_mem.sv:405:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h01d54683;
			// Trace: ../../rtl/local_mem.sv:406:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h02c70633;
			// Trace: ../../rtl/local_mem.sv:407:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h40c787b3;
			// Trace: ../../rtl/local_mem.sv:408:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hfa069ee3;
			// Trace: ../../rtl/local_mem.sv:409:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h0317c833;
			// Trace: ../../rtl/local_mem.sv:410:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hfbdff06f;
			// Trace: ../../rtl/local_mem.sv:411:13
			reg_val_0_80000000[(21 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'hff010113;
			// Trace: ../../rtl/local_mem.sv:412:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00112623;
			// Trace: ../../rtl/local_mem.sv:413:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hfff00793;
			// Trace: ../../rtl/local_mem.sv:414:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:415:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'he11ff0ef;
			// Trace: ../../rtl/local_mem.sv:416:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'hcc3027f3;
			// Trace: ../../rtl/local_mem.sv:417:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h0017b793;
			// Trace: ../../rtl/local_mem.sv:418:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:419:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00c12083;
			// Trace: ../../rtl/local_mem.sv:420:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h01010113;
			// Trace: ../../rtl/local_mem.sv:421:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:422:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hfd010113;
			// Trace: ../../rtl/local_mem.sv:423:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h02112623;
			// Trace: ../../rtl/local_mem.sv:424:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h02812423;
			// Trace: ../../rtl/local_mem.sv:425:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h02912223;
			// Trace: ../../rtl/local_mem.sv:426:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h03212023;
			// Trace: ../../rtl/local_mem.sv:427:13
			reg_val_0_80000000[(22 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'hfc2026f3;
			// Trace: ../../rtl/local_mem.sv:428:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hfc1028f3;
			// Trace: ../../rtl/local_mem.sv:429:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hfc0024f3;
			// Trace: ../../rtl/local_mem.sv:430:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'hcc5027f3;
			// Trace: ../../rtl/local_mem.sv:431:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h01f00713;
			// Trace: ../../rtl/local_mem.sv:432:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h08f74863;
			// Trace: ../../rtl/local_mem.sv:433:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h03148833;
			// Trace: ../../rtl/local_mem.sv:434:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00100713;
			// Trace: ../../rtl/local_mem.sv:435:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00a85463;
			// Trace: ../../rtl/local_mem.sv:436:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h03054733;
			// Trace: ../../rtl/local_mem.sv:437:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h08e6ca63;
			// Trace: ../../rtl/local_mem.sv:438:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h06e7dc63;
			// Trace: ../../rtl/local_mem.sv:439:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hfff68693;
			// Trace: ../../rtl/local_mem.sv:440:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h02e54333;
			// Trace: ../../rtl/local_mem.sv:441:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00030813;
			// Trace: ../../rtl/local_mem.sv:442:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00f69663;
			// Trace: ../../rtl/local_mem.sv:443:13
			reg_val_0_80000000[(23 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h02e56533;
			// Trace: ../../rtl/local_mem.sv:444:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00650833;
			// Trace: ../../rtl/local_mem.sv:445:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h02984933;
			// Trace: ../../rtl/local_mem.sv:446:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h02986433;
			// Trace: ../../rtl/local_mem.sv:447:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h07194c63;
			// Trace: ../../rtl/local_mem.sv:448:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00100513;
			// Trace: ../../rtl/local_mem.sv:449:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h031946b3;
			// Trace: ../../rtl/local_mem.sv:450:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00068663;
			// Trace: ../../rtl/local_mem.sv:451:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00068513;
			// Trace: ../../rtl/local_mem.sv:452:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h031966b3;
			// Trace: ../../rtl/local_mem.sv:453:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00001717;
			// Trace: ../../rtl/local_mem.sv:454:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'he1c70713;
			// Trace: ../../rtl/local_mem.sv:455:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00b12423;
			// Trace: ../../rtl/local_mem.sv:456:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00c12623;
			// Trace: ../../rtl/local_mem.sv:457:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00a12a23;
			// Trace: ../../rtl/local_mem.sv:458:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00d12c23;
			// Trace: ../../rtl/local_mem.sv:459:13
			reg_val_0_80000000[(24 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00012e23;
			// Trace: ../../rtl/local_mem.sv:460:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h02f30333;
			// Trace: ../../rtl/local_mem.sv:461:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00279793;
			// Trace: ../../rtl/local_mem.sv:462:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00f707b3;
			// Trace: ../../rtl/local_mem.sv:463:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00810713;
			// Trace: ../../rtl/local_mem.sv:464:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00e7a023;
			// Trace: ../../rtl/local_mem.sv:465:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00612823;
			// Trace: ../../rtl/local_mem.sv:466:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h03204c63;
			// Trace: ../../rtl/local_mem.sv:467:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h06041663;
			// Trace: ../../rtl/local_mem.sv:468:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h02c12083;
			// Trace: ../../rtl/local_mem.sv:469:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h02812403;
			// Trace: ../../rtl/local_mem.sv:470:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h02412483;
			// Trace: ../../rtl/local_mem.sv:471:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h02012903;
			// Trace: ../../rtl/local_mem.sv:472:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h03010113;
			// Trace: ../../rtl/local_mem.sv:473:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:474:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00068713;
			// Trace: ../../rtl/local_mem.sv:475:13
			reg_val_0_80000000[(25 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'hf6e7c8e3;
			// Trace: ../../rtl/local_mem.sv:476:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hfe1ff06f;
			// Trace: ../../rtl/local_mem.sv:477:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000693;
			// Trace: ../../rtl/local_mem.sv:478:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00100513;
			// Trace: ../../rtl/local_mem.sv:479:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hf99ff06f;
			// Trace: ../../rtl/local_mem.sv:480:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00090793;
			// Trace: ../../rtl/local_mem.sv:481:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h0128d463;
			// Trace: ../../rtl/local_mem.sv:482:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00088793;
			// Trace: ../../rtl/local_mem.sv:483:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00f12e23;
			// Trace: ../../rtl/local_mem.sv:484:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000717;
			// Trace: ../../rtl/local_mem.sv:485:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'hcd070713;
			// Trace: ../../rtl/local_mem.sv:486:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00e7906b;
			// Trace: ../../rtl/local_mem.sv:487:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hfff00793;
			// Trace: ../../rtl/local_mem.sv:488:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:489:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hbd9ff0ef;
			// Trace: ../../rtl/local_mem.sv:490:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hcc3027f3;
			// Trace: ../../rtl/local_mem.sv:491:13
			reg_val_0_80000000[(26 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h0017b793;
			// Trace: ../../rtl/local_mem.sv:492:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:493:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hf8040ee3;
			// Trace: ../../rtl/local_mem.sv:494:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h029904b3;
			// Trace: ../../rtl/local_mem.sv:495:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00100913;
			// Trace: ../../rtl/local_mem.sv:496:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00891833;
			// Trace: ../../rtl/local_mem.sv:497:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hfff80813;
			// Trace: ../../rtl/local_mem.sv:498:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00912823;
			// Trace: ../../rtl/local_mem.sv:499:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h0008006b;
			// Trace: ../../rtl/local_mem.sv:500:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hc61ff0ef;
			// Trace: ../../rtl/local_mem.sv:501:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h0009006b;
			// Trace: ../../rtl/local_mem.sv:502:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h02c12083;
			// Trace: ../../rtl/local_mem.sv:503:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h02812403;
			// Trace: ../../rtl/local_mem.sv:504:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h02412483;
			// Trace: ../../rtl/local_mem.sv:505:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h02012903;
			// Trace: ../../rtl/local_mem.sv:506:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h03010113;
			// Trace: ../../rtl/local_mem.sv:507:13
			reg_val_0_80000000[(27 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:508:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hfd010113;
			// Trace: ../../rtl/local_mem.sv:509:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h02112623;
			// Trace: ../../rtl/local_mem.sv:510:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h02812423;
			// Trace: ../../rtl/local_mem.sv:511:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h02912223;
			// Trace: ../../rtl/local_mem.sv:512:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h03212023;
			// Trace: ../../rtl/local_mem.sv:513:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hfc2028f3;
			// Trace: ../../rtl/local_mem.sv:514:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hfc102373;
			// Trace: ../../rtl/local_mem.sv:515:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hfc0024f3;
			// Trace: ../../rtl/local_mem.sv:516:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hcc5027f3;
			// Trace: ../../rtl/local_mem.sv:517:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h01f00713;
			// Trace: ../../rtl/local_mem.sv:518:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h0ef74663;
			// Trace: ../../rtl/local_mem.sv:519:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00052e03;
			// Trace: ../../rtl/local_mem.sv:520:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00452683;
			// Trace: ../../rtl/local_mem.sv:521:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00852803;
			// Trace: ../../rtl/local_mem.sv:522:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h02930eb3;
			// Trace: ../../rtl/local_mem.sv:523:13
			reg_val_0_80000000[(28 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00100713;
			// Trace: ../../rtl/local_mem.sv:524:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h02de06b3;
			// Trace: ../../rtl/local_mem.sv:525:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h03068833;
			// Trace: ../../rtl/local_mem.sv:526:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h010ed463;
			// Trace: ../../rtl/local_mem.sv:527:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h03d84733;
			// Trace: ../../rtl/local_mem.sv:528:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h0ce8ce63;
			// Trace: ../../rtl/local_mem.sv:529:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h0ce7d063;
			// Trace: ../../rtl/local_mem.sv:530:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hfff88893;
			// Trace: ../../rtl/local_mem.sv:531:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h02e84f33;
			// Trace: ../../rtl/local_mem.sv:532:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h000f0413;
			// Trace: ../../rtl/local_mem.sv:533:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00f89663;
			// Trace: ../../rtl/local_mem.sv:534:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h02e86733;
			// Trace: ../../rtl/local_mem.sv:535:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01e70433;
			// Trace: ../../rtl/local_mem.sv:536:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h02944933;
			// Trace: ../../rtl/local_mem.sv:537:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h02946433;
			// Trace: ../../rtl/local_mem.sv:538:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h0c694063;
			// Trace: ../../rtl/local_mem.sv:539:13
			reg_val_0_80000000[(29 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00100293;
			// Trace: ../../rtl/local_mem.sv:540:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h02694fb3;
			// Trace: ../../rtl/local_mem.sv:541:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h000f8663;
			// Trace: ../../rtl/local_mem.sv:542:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h000f8293;
			// Trace: ../../rtl/local_mem.sv:543:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h02696fb3;
			// Trace: ../../rtl/local_mem.sv:544:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'hd006f7d3;
			// Trace: ../../rtl/local_mem.sv:545:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hfffe0893;
			// Trace: ../../rtl/local_mem.sv:546:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hfff68e93;
			// Trace: ../../rtl/local_mem.sv:547:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'he0078853;
			// Trace: ../../rtl/local_mem.sv:548:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hd00e77d3;
			// Trace: ../../rtl/local_mem.sv:549:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00def6b3;
			// Trace: ../../rtl/local_mem.sv:550:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h01c8fe33;
			// Trace: ../../rtl/local_mem.sv:551:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'he0078753;
			// Trace: ../../rtl/local_mem.sv:552:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h41785813;
			// Trace: ../../rtl/local_mem.sv:553:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00001897;
			// Trace: ../../rtl/local_mem.sv:554:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hc8c88893;
			// Trace: ../../rtl/local_mem.sv:555:13
			reg_val_0_80000000[(30 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h41775713;
			// Trace: ../../rtl/local_mem.sv:556:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h0016b693;
			// Trace: ../../rtl/local_mem.sv:557:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h001e3e13;
			// Trace: ../../rtl/local_mem.sv:558:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'hf8180813;
			// Trace: ../../rtl/local_mem.sv:559:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hf8170713;
			// Trace: ../../rtl/local_mem.sv:560:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00a12023;
			// Trace: ../../rtl/local_mem.sv:561:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00b12223;
			// Trace: ../../rtl/local_mem.sv:562:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00c12423;
			// Trace: ../../rtl/local_mem.sv:563:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00512823;
			// Trace: ../../rtl/local_mem.sv:564:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h01f12a23;
			// Trace: ../../rtl/local_mem.sv:565:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00012c23;
			// Trace: ../../rtl/local_mem.sv:566:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00d10e23;
			// Trace: ../../rtl/local_mem.sv:567:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01c10ea3;
			// Trace: ../../rtl/local_mem.sv:568:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h01010f23;
			// Trace: ../../rtl/local_mem.sv:569:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00e10fa3;
			// Trace: ../../rtl/local_mem.sv:570:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h02ff0f33;
			// Trace: ../../rtl/local_mem.sv:571:13
			reg_val_0_80000000[(31 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00279793;
			// Trace: ../../rtl/local_mem.sv:572:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00f887b3;
			// Trace: ../../rtl/local_mem.sv:573:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h0027a023;
			// Trace: ../../rtl/local_mem.sv:574:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h01e12623;
			// Trace: ../../rtl/local_mem.sv:575:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h03204c63;
			// Trace: ../../rtl/local_mem.sv:576:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h06041663;
			// Trace: ../../rtl/local_mem.sv:577:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h02c12083;
			// Trace: ../../rtl/local_mem.sv:578:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h02812403;
			// Trace: ../../rtl/local_mem.sv:579:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h02412483;
			// Trace: ../../rtl/local_mem.sv:580:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h02012903;
			// Trace: ../../rtl/local_mem.sv:581:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h03010113;
			// Trace: ../../rtl/local_mem.sv:582:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:583:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00088713;
			// Trace: ../../rtl/local_mem.sv:584:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hf2e7c4e3;
			// Trace: ../../rtl/local_mem.sv:585:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hfe1ff06f;
			// Trace: ../../rtl/local_mem.sv:586:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000f93;
			// Trace: ../../rtl/local_mem.sv:587:13
			reg_val_0_80000000[(32 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00100293;
			// Trace: ../../rtl/local_mem.sv:588:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hf51ff06f;
			// Trace: ../../rtl/local_mem.sv:589:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00090793;
			// Trace: ../../rtl/local_mem.sv:590:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h01235463;
			// Trace: ../../rtl/local_mem.sv:591:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00030793;
			// Trace: ../../rtl/local_mem.sv:592:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00f12c23;
			// Trace: ../../rtl/local_mem.sv:593:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000717;
			// Trace: ../../rtl/local_mem.sv:594:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hd2870713;
			// Trace: ../../rtl/local_mem.sv:595:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00e7906b;
			// Trace: ../../rtl/local_mem.sv:596:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hfff00793;
			// Trace: ../../rtl/local_mem.sv:597:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:598:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hb35ff0ef;
			// Trace: ../../rtl/local_mem.sv:599:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hcc3027f3;
			// Trace: ../../rtl/local_mem.sv:600:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h0017b793;
			// Trace: ../../rtl/local_mem.sv:601:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h0007806b;
			// Trace: ../../rtl/local_mem.sv:602:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hf8040ee3;
			// Trace: ../../rtl/local_mem.sv:603:13
			reg_val_0_80000000[(33 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h029904b3;
			// Trace: ../../rtl/local_mem.sv:604:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00100913;
			// Trace: ../../rtl/local_mem.sv:605:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00891433;
			// Trace: ../../rtl/local_mem.sv:606:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'hfff40413;
			// Trace: ../../rtl/local_mem.sv:607:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00912623;
			// Trace: ../../rtl/local_mem.sv:608:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h0004006b;
			// Trace: ../../rtl/local_mem.sv:609:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hc45ff0ef;
			// Trace: ../../rtl/local_mem.sv:610:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h0009006b;
			// Trace: ../../rtl/local_mem.sv:611:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h02c12083;
			// Trace: ../../rtl/local_mem.sv:612:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h02812403;
			// Trace: ../../rtl/local_mem.sv:613:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h02412483;
			// Trace: ../../rtl/local_mem.sv:614:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h02012903;
			// Trace: ../../rtl/local_mem.sv:615:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h03010113;
			// Trace: ../../rtl/local_mem.sv:616:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:617:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hfe810113;
			// Trace: ../../rtl/local_mem.sv:618:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00112a23;
			// Trace: ../../rtl/local_mem.sv:619:13
			reg_val_0_80000000[(34 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h01412823;
			// Trace: ../../rtl/local_mem.sv:620:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h01312623;
			// Trace: ../../rtl/local_mem.sv:621:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h01212423;
			// Trace: ../../rtl/local_mem.sv:622:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00912223;
			// Trace: ../../rtl/local_mem.sv:623:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00812023;
			// Trace: ../../rtl/local_mem.sv:624:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00050a13;
			// Trace: ../../rtl/local_mem.sv:625:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00058993;
			// Trace: ../../rtl/local_mem.sv:626:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hfc002973;
			// Trace: ../../rtl/local_mem.sv:627:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hcc0024f3;
			// Trace: ../../rtl/local_mem.sv:628:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000413;
			// Trace: ../../rtl/local_mem.sv:629:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h409402b3;
			// Trace: ../../rtl/local_mem.sv:630:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h0012b313;
			// Trace: ../../rtl/local_mem.sv:631:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h0003206b;
			// Trace: ../../rtl/local_mem.sv:632:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00029663;
			// Trace: ../../rtl/local_mem.sv:633:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00098513;
			// Trace: ../../rtl/local_mem.sv:634:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h000a00e7;
			// Trace: ../../rtl/local_mem.sv:635:13
			reg_val_0_80000000[(35 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h0000306b;
			// Trace: ../../rtl/local_mem.sv:636:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00140413;
			// Trace: ../../rtl/local_mem.sv:637:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hff2440e3;
			// Trace: ../../rtl/local_mem.sv:638:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h01412083;
			// Trace: ../../rtl/local_mem.sv:639:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h01012a03;
			// Trace: ../../rtl/local_mem.sv:640:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00c12983;
			// Trace: ../../rtl/local_mem.sv:641:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00812903;
			// Trace: ../../rtl/local_mem.sv:642:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00412483;
			// Trace: ../../rtl/local_mem.sv:643:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00012403;
			// Trace: ../../rtl/local_mem.sv:644:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h01810113;
			// Trace: ../../rtl/local_mem.sv:645:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:646:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:647:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:648:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:649:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:650:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:651:13
			reg_val_0_80000000[(36 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:652:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:653:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:654:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:655:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:656:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:657:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:658:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:659:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:660:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:661:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:662:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:663:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:664:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:665:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:666:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:667:13
			reg_val_0_80000000[(37 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:668:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:669:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:670:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00050593;
			// Trace: ../../rtl/local_mem.sv:671:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000693;
			// Trace: ../../rtl/local_mem.sv:672:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000613;
			// Trace: ../../rtl/local_mem.sv:673:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:674:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h2300006f;
			// Trace: ../../rtl/local_mem.sv:675:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hff010113;
			// Trace: ../../rtl/local_mem.sv:676:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000593;
			// Trace: ../../rtl/local_mem.sv:677:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00812423;
			// Trace: ../../rtl/local_mem.sv:678:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00112623;
			// Trace: ../../rtl/local_mem.sv:679:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00050413;
			// Trace: ../../rtl/local_mem.sv:680:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h2b4000ef;
			// Trace: ../../rtl/local_mem.sv:681:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h800017b7;
			// Trace: ../../rtl/local_mem.sv:682:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h4387a503;
			// Trace: ../../rtl/local_mem.sv:683:13
			reg_val_0_80000000[(38 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h03c52783;
			// Trace: ../../rtl/local_mem.sv:684:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00078463;
			// Trace: ../../rtl/local_mem.sv:685:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h000780e7;
			// Trace: ../../rtl/local_mem.sv:686:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00040513;
			// Trace: ../../rtl/local_mem.sv:687:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hec8ff0ef;
			// Trace: ../../rtl/local_mem.sv:688:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00a5c7b3;
			// Trace: ../../rtl/local_mem.sv:689:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h0037f793;
			// Trace: ../../rtl/local_mem.sv:690:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00c508b3;
			// Trace: ../../rtl/local_mem.sv:691:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h06079263;
			// Trace: ../../rtl/local_mem.sv:692:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00300793;
			// Trace: ../../rtl/local_mem.sv:693:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h04c7fe63;
			// Trace: ../../rtl/local_mem.sv:694:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00357793;
			// Trace: ../../rtl/local_mem.sv:695:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00050713;
			// Trace: ../../rtl/local_mem.sv:696:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h06079863;
			// Trace: ../../rtl/local_mem.sv:697:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hffc8f613;
			// Trace: ../../rtl/local_mem.sv:698:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hfe060793;
			// Trace: ../../rtl/local_mem.sv:699:13
			reg_val_0_80000000[(39 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h08f76c63;
			// Trace: ../../rtl/local_mem.sv:700:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h02c77c63;
			// Trace: ../../rtl/local_mem.sv:701:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00058693;
			// Trace: ../../rtl/local_mem.sv:702:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00070793;
			// Trace: ../../rtl/local_mem.sv:703:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h0006a803;
			// Trace: ../../rtl/local_mem.sv:704:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00478793;
			// Trace: ../../rtl/local_mem.sv:705:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00468693;
			// Trace: ../../rtl/local_mem.sv:706:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hff07ae23;
			// Trace: ../../rtl/local_mem.sv:707:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hfec7e8e3;
			// Trace: ../../rtl/local_mem.sv:708:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hfff60793;
			// Trace: ../../rtl/local_mem.sv:709:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h40e787b3;
			// Trace: ../../rtl/local_mem.sv:710:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hffc7f793;
			// Trace: ../../rtl/local_mem.sv:711:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00478793;
			// Trace: ../../rtl/local_mem.sv:712:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00f70733;
			// Trace: ../../rtl/local_mem.sv:713:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00f585b3;
			// Trace: ../../rtl/local_mem.sv:714:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h01176863;
			// Trace: ../../rtl/local_mem.sv:715:13
			reg_val_0_80000000[(40 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:716:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00050713;
			// Trace: ../../rtl/local_mem.sv:717:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hff157ce3;
			// Trace: ../../rtl/local_mem.sv:718:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h0005c783;
			// Trace: ../../rtl/local_mem.sv:719:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00170713;
			// Trace: ../../rtl/local_mem.sv:720:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00158593;
			// Trace: ../../rtl/local_mem.sv:721:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hfef70fa3;
			// Trace: ../../rtl/local_mem.sv:722:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hff1768e3;
			// Trace: ../../rtl/local_mem.sv:723:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:724:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h0005c683;
			// Trace: ../../rtl/local_mem.sv:725:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00170713;
			// Trace: ../../rtl/local_mem.sv:726:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00377793;
			// Trace: ../../rtl/local_mem.sv:727:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hfed70fa3;
			// Trace: ../../rtl/local_mem.sv:728:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00158593;
			// Trace: ../../rtl/local_mem.sv:729:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hf80780e3;
			// Trace: ../../rtl/local_mem.sv:730:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h0005c683;
			// Trace: ../../rtl/local_mem.sv:731:13
			reg_val_0_80000000[(41 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00170713;
			// Trace: ../../rtl/local_mem.sv:732:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00377793;
			// Trace: ../../rtl/local_mem.sv:733:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hfed70fa3;
			// Trace: ../../rtl/local_mem.sv:734:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00158593;
			// Trace: ../../rtl/local_mem.sv:735:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hfc079ae3;
			// Trace: ../../rtl/local_mem.sv:736:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'hf65ff06f;
			// Trace: ../../rtl/local_mem.sv:737:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h0045a683;
			// Trace: ../../rtl/local_mem.sv:738:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h0005a283;
			// Trace: ../../rtl/local_mem.sv:739:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h0085af83;
			// Trace: ../../rtl/local_mem.sv:740:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00c5af03;
			// Trace: ../../rtl/local_mem.sv:741:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h0105ae83;
			// Trace: ../../rtl/local_mem.sv:742:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h0145ae03;
			// Trace: ../../rtl/local_mem.sv:743:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h0185a303;
			// Trace: ../../rtl/local_mem.sv:744:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h01c5a803;
			// Trace: ../../rtl/local_mem.sv:745:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00d72223;
			// Trace: ../../rtl/local_mem.sv:746:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h0205a683;
			// Trace: ../../rtl/local_mem.sv:747:13
			reg_val_0_80000000[(42 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00572023;
			// Trace: ../../rtl/local_mem.sv:748:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h01f72423;
			// Trace: ../../rtl/local_mem.sv:749:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h01e72623;
			// Trace: ../../rtl/local_mem.sv:750:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h01d72823;
			// Trace: ../../rtl/local_mem.sv:751:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h01c72a23;
			// Trace: ../../rtl/local_mem.sv:752:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00672c23;
			// Trace: ../../rtl/local_mem.sv:753:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h01072e23;
			// Trace: ../../rtl/local_mem.sv:754:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h02d72023;
			// Trace: ../../rtl/local_mem.sv:755:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h02470713;
			// Trace: ../../rtl/local_mem.sv:756:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h02458593;
			// Trace: ../../rtl/local_mem.sv:757:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'hfaf768e3;
			// Trace: ../../rtl/local_mem.sv:758:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'hf19ff06f;
			// Trace: ../../rtl/local_mem.sv:759:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00f00313;
			// Trace: ../../rtl/local_mem.sv:760:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00050713;
			// Trace: ../../rtl/local_mem.sv:761:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h02c37e63;
			// Trace: ../../rtl/local_mem.sv:762:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00f77793;
			// Trace: ../../rtl/local_mem.sv:763:13
			reg_val_0_80000000[(43 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h0a079063;
			// Trace: ../../rtl/local_mem.sv:764:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h08059263;
			// Trace: ../../rtl/local_mem.sv:765:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hff067693;
			// Trace: ../../rtl/local_mem.sv:766:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00f67613;
			// Trace: ../../rtl/local_mem.sv:767:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00e686b3;
			// Trace: ../../rtl/local_mem.sv:768:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00b72023;
			// Trace: ../../rtl/local_mem.sv:769:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00b72223;
			// Trace: ../../rtl/local_mem.sv:770:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00b72423;
			// Trace: ../../rtl/local_mem.sv:771:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00b72623;
			// Trace: ../../rtl/local_mem.sv:772:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h01070713;
			// Trace: ../../rtl/local_mem.sv:773:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'hfed766e3;
			// Trace: ../../rtl/local_mem.sv:774:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00061463;
			// Trace: ../../rtl/local_mem.sv:775:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:776:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h40c306b3;
			// Trace: ../../rtl/local_mem.sv:777:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00269693;
			// Trace: ../../rtl/local_mem.sv:778:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000297;
			// Trace: ../../rtl/local_mem.sv:779:13
			reg_val_0_80000000[(44 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h005686b3;
			// Trace: ../../rtl/local_mem.sv:780:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00c68067;
			// Trace: ../../rtl/local_mem.sv:781:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00b70723;
			// Trace: ../../rtl/local_mem.sv:782:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00b706a3;
			// Trace: ../../rtl/local_mem.sv:783:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00b70623;
			// Trace: ../../rtl/local_mem.sv:784:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00b705a3;
			// Trace: ../../rtl/local_mem.sv:785:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00b70523;
			// Trace: ../../rtl/local_mem.sv:786:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00b704a3;
			// Trace: ../../rtl/local_mem.sv:787:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00b70423;
			// Trace: ../../rtl/local_mem.sv:788:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00b703a3;
			// Trace: ../../rtl/local_mem.sv:789:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00b70323;
			// Trace: ../../rtl/local_mem.sv:790:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00b702a3;
			// Trace: ../../rtl/local_mem.sv:791:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00b70223;
			// Trace: ../../rtl/local_mem.sv:792:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00b701a3;
			// Trace: ../../rtl/local_mem.sv:793:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00b70123;
			// Trace: ../../rtl/local_mem.sv:794:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00b700a3;
			// Trace: ../../rtl/local_mem.sv:795:13
			reg_val_0_80000000[(45 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00b70023;
			// Trace: ../../rtl/local_mem.sv:796:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:797:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h0ff5f593;
			// Trace: ../../rtl/local_mem.sv:798:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00859693;
			// Trace: ../../rtl/local_mem.sv:799:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00d5e5b3;
			// Trace: ../../rtl/local_mem.sv:800:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h01059693;
			// Trace: ../../rtl/local_mem.sv:801:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00d5e5b3;
			// Trace: ../../rtl/local_mem.sv:802:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hf6dff06f;
			// Trace: ../../rtl/local_mem.sv:803:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00279693;
			// Trace: ../../rtl/local_mem.sv:804:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000297;
			// Trace: ../../rtl/local_mem.sv:805:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h005686b3;
			// Trace: ../../rtl/local_mem.sv:806:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00008293;
			// Trace: ../../rtl/local_mem.sv:807:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hfa0680e7;
			// Trace: ../../rtl/local_mem.sv:808:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00028093;
			// Trace: ../../rtl/local_mem.sv:809:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hff078793;
			// Trace: ../../rtl/local_mem.sv:810:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h40f70733;
			// Trace: ../../rtl/local_mem.sv:811:13
			reg_val_0_80000000[(46 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00f60633;
			// Trace: ../../rtl/local_mem.sv:812:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hf6c378e3;
			// Trace: ../../rtl/local_mem.sv:813:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hf3dff06f;
			// Trace: ../../rtl/local_mem.sv:814:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h800017b7;
			// Trace: ../../rtl/local_mem.sv:815:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h4387a703;
			// Trace: ../../rtl/local_mem.sv:816:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h14872783;
			// Trace: ../../rtl/local_mem.sv:817:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h04078c63;
			// Trace: ../../rtl/local_mem.sv:818:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h0047a703;
			// Trace: ../../rtl/local_mem.sv:819:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h01f00813;
			// Trace: ../../rtl/local_mem.sv:820:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h06e84e63;
			// Trace: ../../rtl/local_mem.sv:821:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00271813;
			// Trace: ../../rtl/local_mem.sv:822:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h02050663;
			// Trace: ../../rtl/local_mem.sv:823:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01078333;
			// Trace: ../../rtl/local_mem.sv:824:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h08c32423;
			// Trace: ../../rtl/local_mem.sv:825:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h1887a883;
			// Trace: ../../rtl/local_mem.sv:826:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00100613;
			// Trace: ../../rtl/local_mem.sv:827:13
			reg_val_0_80000000[(47 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00e61633;
			// Trace: ../../rtl/local_mem.sv:828:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00c8e8b3;
			// Trace: ../../rtl/local_mem.sv:829:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h1917a423;
			// Trace: ../../rtl/local_mem.sv:830:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h10d32423;
			// Trace: ../../rtl/local_mem.sv:831:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00200693;
			// Trace: ../../rtl/local_mem.sv:832:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h02d50463;
			// Trace: ../../rtl/local_mem.sv:833:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00170713;
			// Trace: ../../rtl/local_mem.sv:834:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00e7a223;
			// Trace: ../../rtl/local_mem.sv:835:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h010787b3;
			// Trace: ../../rtl/local_mem.sv:836:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00b7a423;
			// Trace: ../../rtl/local_mem.sv:837:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:838:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:839:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h14c70793;
			// Trace: ../../rtl/local_mem.sv:840:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h14f72423;
			// Trace: ../../rtl/local_mem.sv:841:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hfa5ff06f;
			// Trace: ../../rtl/local_mem.sv:842:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h18c7a683;
			// Trace: ../../rtl/local_mem.sv:843:13
			reg_val_0_80000000[(48 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00170713;
			// Trace: ../../rtl/local_mem.sv:844:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00e7a223;
			// Trace: ../../rtl/local_mem.sv:845:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00c6e633;
			// Trace: ../../rtl/local_mem.sv:846:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h18c7a623;
			// Trace: ../../rtl/local_mem.sv:847:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h010787b3;
			// Trace: ../../rtl/local_mem.sv:848:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00b7a423;
			// Trace: ../../rtl/local_mem.sv:849:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000513;
			// Trace: ../../rtl/local_mem.sv:850:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:851:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hfff00513;
			// Trace: ../../rtl/local_mem.sv:852:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:853:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'hfd010113;
			// Trace: ../../rtl/local_mem.sv:854:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h800017b7;
			// Trace: ../../rtl/local_mem.sv:855:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01412c23;
			// Trace: ../../rtl/local_mem.sv:856:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h4387aa03;
			// Trace: ../../rtl/local_mem.sv:857:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h03212023;
			// Trace: ../../rtl/local_mem.sv:858:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h02112623;
			// Trace: ../../rtl/local_mem.sv:859:13
			reg_val_0_80000000[(49 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h148a2903;
			// Trace: ../../rtl/local_mem.sv:860:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h02812423;
			// Trace: ../../rtl/local_mem.sv:861:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h02912223;
			// Trace: ../../rtl/local_mem.sv:862:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h01312e23;
			// Trace: ../../rtl/local_mem.sv:863:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h01512a23;
			// Trace: ../../rtl/local_mem.sv:864:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h01612823;
			// Trace: ../../rtl/local_mem.sv:865:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h01712623;
			// Trace: ../../rtl/local_mem.sv:866:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h01812423;
			// Trace: ../../rtl/local_mem.sv:867:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h04090063;
			// Trace: ../../rtl/local_mem.sv:868:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00050b13;
			// Trace: ../../rtl/local_mem.sv:869:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00058b93;
			// Trace: ../../rtl/local_mem.sv:870:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00100a93;
			// Trace: ../../rtl/local_mem.sv:871:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hfff00993;
			// Trace: ../../rtl/local_mem.sv:872:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00492483;
			// Trace: ../../rtl/local_mem.sv:873:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hfff48413;
			// Trace: ../../rtl/local_mem.sv:874:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h02044263;
			// Trace: ../../rtl/local_mem.sv:875:13
			reg_val_0_80000000[(50 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00249493;
			// Trace: ../../rtl/local_mem.sv:876:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h009904b3;
			// Trace: ../../rtl/local_mem.sv:877:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h040b8463;
			// Trace: ../../rtl/local_mem.sv:878:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h1044a783;
			// Trace: ../../rtl/local_mem.sv:879:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h05778063;
			// Trace: ../../rtl/local_mem.sv:880:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'hfff40413;
			// Trace: ../../rtl/local_mem.sv:881:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hffc48493;
			// Trace: ../../rtl/local_mem.sv:882:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hff3416e3;
			// Trace: ../../rtl/local_mem.sv:883:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h02c12083;
			// Trace: ../../rtl/local_mem.sv:884:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h02812403;
			// Trace: ../../rtl/local_mem.sv:885:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h02412483;
			// Trace: ../../rtl/local_mem.sv:886:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h02012903;
			// Trace: ../../rtl/local_mem.sv:887:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h01c12983;
			// Trace: ../../rtl/local_mem.sv:888:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h01812a03;
			// Trace: ../../rtl/local_mem.sv:889:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h01412a83;
			// Trace: ../../rtl/local_mem.sv:890:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h01012b03;
			// Trace: ../../rtl/local_mem.sv:891:13
			reg_val_0_80000000[(51 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00c12b83;
			// Trace: ../../rtl/local_mem.sv:892:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00812c03;
			// Trace: ../../rtl/local_mem.sv:893:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h03010113;
			// Trace: ../../rtl/local_mem.sv:894:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00008067;
			// Trace: ../../rtl/local_mem.sv:895:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00492783;
			// Trace: ../../rtl/local_mem.sv:896:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h0044a683;
			// Trace: ../../rtl/local_mem.sv:897:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hfff78793;
			// Trace: ../../rtl/local_mem.sv:898:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h04878e63;
			// Trace: ../../rtl/local_mem.sv:899:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h0004a223;
			// Trace: ../../rtl/local_mem.sv:900:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hfa0688e3;
			// Trace: ../../rtl/local_mem.sv:901:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h18892783;
			// Trace: ../../rtl/local_mem.sv:902:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h008a9733;
			// Trace: ../../rtl/local_mem.sv:903:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00492c03;
			// Trace: ../../rtl/local_mem.sv:904:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00f777b3;
			// Trace: ../../rtl/local_mem.sv:905:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h02079263;
			// Trace: ../../rtl/local_mem.sv:906:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h000680e7;
			// Trace: ../../rtl/local_mem.sv:907:13
			reg_val_0_80000000[(52 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00492703;
			// Trace: ../../rtl/local_mem.sv:908:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h148a2783;
			// Trace: ../../rtl/local_mem.sv:909:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h01871463;
			// Trace: ../../rtl/local_mem.sv:910:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'hf8f904e3;
			// Trace: ../../rtl/local_mem.sv:911:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hf80788e3;
			// Trace: ../../rtl/local_mem.sv:912:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00078913;
			// Trace: ../../rtl/local_mem.sv:913:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'hf5dff06f;
			// Trace: ../../rtl/local_mem.sv:914:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h18c92783;
			// Trace: ../../rtl/local_mem.sv:915:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h0844a583;
			// Trace: ../../rtl/local_mem.sv:916:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00f77733;
			// Trace: ../../rtl/local_mem.sv:917:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00071c63;
			// Trace: ../../rtl/local_mem.sv:918:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h000b0513;
			// Trace: ../../rtl/local_mem.sv:919:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h000680e7;
			// Trace: ../../rtl/local_mem.sv:920:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hfcdff06f;
			// Trace: ../../rtl/local_mem.sv:921:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00892223;
			// Trace: ../../rtl/local_mem.sv:922:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hfa9ff06f;
			// Trace: ../../rtl/local_mem.sv:923:13
			reg_val_0_80000000[(53 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00058513;
			// Trace: ../../rtl/local_mem.sv:924:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h000680e7;
			// Trace: ../../rtl/local_mem.sv:925:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hfb9ff06f;
			// Trace: ../../rtl/local_mem.sv:926:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:927:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:928:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00527a03;
			// Trace: ../../rtl/local_mem.sv:929:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h01017c01;
			// Trace: ../../rtl/local_mem.sv:930:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00020d1b;
			// Trace: ../../rtl/local_mem.sv:931:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:932:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000018;
			// Trace: ../../rtl/local_mem.sv:933:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'hfffffb84;
			// Trace: ../../rtl/local_mem.sv:934:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:935:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:936:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:937:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h0000002c;
			// Trace: ../../rtl/local_mem.sv:938:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'hfffffb78;
			// Trace: ../../rtl/local_mem.sv:939:13
			reg_val_0_80000000[(54 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:940:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:941:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:942:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000040;
			// Trace: ../../rtl/local_mem.sv:943:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'hfffffb6c;
			// Trace: ../../rtl/local_mem.sv:944:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:945:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:946:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:947:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000054;
			// Trace: ../../rtl/local_mem.sv:948:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'hfffffb60;
			// Trace: ../../rtl/local_mem.sv:949:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:950:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:951:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:952:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000068;
			// Trace: ../../rtl/local_mem.sv:953:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'hfffffb54;
			// Trace: ../../rtl/local_mem.sv:954:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:955:13
			reg_val_0_80000000[(55 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:956:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:957:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h0000007c;
			// Trace: ../../rtl/local_mem.sv:958:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'hfffffb48;
			// Trace: ../../rtl/local_mem.sv:959:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:960:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:961:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:962:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000090;
			// Trace: ../../rtl/local_mem.sv:963:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'hfffffb3c;
			// Trace: ../../rtl/local_mem.sv:964:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:965:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:966:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:967:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h000000a4;
			// Trace: ../../rtl/local_mem.sv:968:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'hfffffb30;
			// Trace: ../../rtl/local_mem.sv:969:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:970:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:971:13
			reg_val_0_80000000[(56 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:972:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h000000b8;
			// Trace: ../../rtl/local_mem.sv:973:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'hfffffb24;
			// Trace: ../../rtl/local_mem.sv:974:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:975:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:976:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:977:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h000000cc;
			// Trace: ../../rtl/local_mem.sv:978:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'hfffffb18;
			// Trace: ../../rtl/local_mem.sv:979:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:980:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:981:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:982:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h000000e0;
			// Trace: ../../rtl/local_mem.sv:983:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'hfffffb0c;
			// Trace: ../../rtl/local_mem.sv:984:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:985:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:986:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000010;
			// Trace: ../../rtl/local_mem.sv:987:13
			reg_val_0_80000000[(57 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h000000f4;
			// Trace: ../../rtl/local_mem.sv:988:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'hfffffb00;
			// Trace: ../../rtl/local_mem.sv:989:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000008;
			// Trace: ../../rtl/local_mem.sv:990:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:992:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:993:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:994:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:995:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:996:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:997:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:998:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:999:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1000:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1001:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1002:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1003:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1004:13
			reg_val_0_80000000[(58 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1005:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1006:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1007:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1008:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1009:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1010:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1011:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1012:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1013:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1014:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1015:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1016:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1017:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1018:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1019:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1020:13
			reg_val_0_80000000[(59 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1021:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1022:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1023:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1024:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1025:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1026:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1027:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1028:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1029:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1030:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1031:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1032:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1033:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1034:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1035:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1036:13
			reg_val_0_80000000[(60 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1037:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1038:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1039:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1040:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1041:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1042:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1043:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1044:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1045:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1046:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1047:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1048:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1049:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1050:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1051:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1052:13
			reg_val_0_80000000[(61 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1053:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1054:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1055:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1056:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1057:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1058:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1059:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1060:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1061:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1062:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1063:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1064:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1065:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1066:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1067:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1068:13
			reg_val_0_80000000[(62 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1069:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1070:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1071:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1072:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1073:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1074:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1075:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1076:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1077:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1078:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1079:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1080:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1081:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1082:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1083:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1084:13
			reg_val_0_80000000[(63 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
		end
		else
			// Trace: ../../rtl/local_mem.sv:1088:13
			reg_val_0_80000000 = next_reg_val_0_80000000;
	end
	// Trace: ../../rtl/local_mem.sv:1092:5
	always @(*) begin : WRITE_LOGIC_0_80000000
		// Trace: ../../rtl/local_mem.sv:1094:9
		begin : sv2v_autoblock_1
			// Trace: ../../rtl/local_mem.sv:1094:14
			reg signed [31:0] i;
			// Trace: ../../rtl/local_mem.sv:1094:14
			for (i = 0; i < 64; i = i + 1)
				begin
					// Trace: ../../rtl/local_mem.sv:1096:13
					next_reg_val_0_80000000[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8] = reg_val_0_80000000[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8];
				end
		end
		if (wen_0_80000000)
			// Trace: ../../rtl/local_mem.sv:1101:13
			next_reg_val_0_80000000[wsel_0_80000000 * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8] = wdata_0_80000000;
	end
	// Trace: ../../rtl/local_mem.sv:1105:5
	always @(*) begin : READ_LOGIC_0_80000000
		// Trace: ../../rtl/local_mem.sv:1107:9
		rdata_0_80000000 = reg_val_0_80000000[rsel_0_80000000 * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8];
	end
	// Trace: ../../rtl/local_mem.sv:1111:5
	reg wen_1_80001000;
	// Trace: ../../rtl/local_mem.sv:1112:5
	reg [0:0] wsel_1_80001000;
	// Trace: ../../rtl/local_mem.sv:1114:5
	reg [((0 || 0 ? 16 : 64) * 8) - 1:0] wdata_1_80001000;
	// Trace: ../../rtl/local_mem.sv:1115:5
	reg [0:0] rsel_1_80001000;
	// Trace: ../../rtl/local_mem.sv:1117:5
	reg [((0 || 0 ? 16 : 64) * 8) - 1:0] rdata_1_80001000;
	// Trace: ../../rtl/local_mem.sv:1119:5
	reg [(2 * ((0 || 0 ? 16 : 64) * 8)) - 1:0] reg_val_1_80001000;
	// Trace: ../../rtl/local_mem.sv:1120:5
	reg [(2 * ((0 || 0 ? 16 : 64) * 8)) - 1:0] next_reg_val_1_80001000;
	// Trace: ../../rtl/local_mem.sv:1122:5
	always @(posedge clk) begin : REGISTER_LOGIC_1_80001000
		// Trace: ../../rtl/local_mem.sv:1123:9
		if (reset) begin
			// Trace: ../../rtl/local_mem.sv:1126:13
			reg_val_1_80001000[31-:32] <= 32'h8000007c;
			// Trace: ../../rtl/local_mem.sv:1128:13
			reg_val_1_80001000[63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1129:13
			reg_val_1_80001000[95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1130:13
			reg_val_1_80001000[127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1131:13
			reg_val_1_80001000[159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1132:13
			reg_val_1_80001000[191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1133:13
			reg_val_1_80001000[223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1134:13
			reg_val_1_80001000[255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1135:13
			reg_val_1_80001000[287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1136:13
			reg_val_1_80001000[319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1137:13
			reg_val_1_80001000[351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1138:13
			reg_val_1_80001000[383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1139:13
			reg_val_1_80001000[415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1140:13
			reg_val_1_80001000[447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1141:13
			reg_val_1_80001000[479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1142:13
			reg_val_1_80001000[511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1143:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1144:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1145:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1146:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1147:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1148:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1149:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1150:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1151:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1152:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1153:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1154:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1155:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1156:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1157:13
			reg_val_1_80001000[((0 || 0 ? 16 : 64) * 8) + 511-:32] <= 32'h00000000;
		end
		else
			// Trace: ../../rtl/local_mem.sv:1161:13
			reg_val_1_80001000 = next_reg_val_1_80001000;
	end
	// Trace: ../../rtl/local_mem.sv:1165:5
	always @(*) begin : WRITE_LOGIC_1_80001000
		// Trace: ../../rtl/local_mem.sv:1167:9
		begin : sv2v_autoblock_2
			// Trace: ../../rtl/local_mem.sv:1167:14
			reg signed [31:0] i;
			// Trace: ../../rtl/local_mem.sv:1167:14
			for (i = 0; i < 1; i = i + 1)
				begin
					// Trace: ../../rtl/local_mem.sv:1169:13
					next_reg_val_1_80001000[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8] = reg_val_1_80001000[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8];
				end
		end
		if (wen_1_80001000)
			// Trace: ../../rtl/local_mem.sv:1174:13
			next_reg_val_1_80001000[wsel_1_80001000 * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8] = wdata_1_80001000;
	end
	// Trace: ../../rtl/local_mem.sv:1178:5
	always @(*) begin : READ_LOGIC_1_80001000
		// Trace: ../../rtl/local_mem.sv:1180:9
		rdata_1_80001000 = reg_val_1_80001000[rsel_1_80001000 * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8];
	end
	// Trace: ../../rtl/local_mem.sv:1184:5
	reg wen_2_80001008;
	// Trace: ../../rtl/local_mem.sv:1185:5
	reg [4:0] wsel_2_80001008;
	// Trace: ../../rtl/local_mem.sv:1186:5
	reg [((0 || 0 ? 16 : 64) * 8) - 1:0] wdata_2_80001008;
	// Trace: ../../rtl/local_mem.sv:1187:5
	reg [4:0] rsel_2_80001008;
	// Trace: ../../rtl/local_mem.sv:1188:5
	reg [((0 || 0 ? 16 : 64) * 8) - 1:0] rdata_2_80001008;
	// Trace: ../../rtl/local_mem.sv:1190:5
	reg [(32 * ((0 || 0 ? 16 : 64) * 8)) - 1:0] reg_val_2_80001008;
	// Trace: ../../rtl/local_mem.sv:1191:5
	reg [(32 * ((0 || 0 ? 16 : 64) * 8)) - 1:0] next_reg_val_2_80001008;
	// Trace: ../../rtl/local_mem.sv:1193:5
	always @(posedge clk) begin : REGISTER_LOGIC_2_80001008
		// Trace: ../../rtl/local_mem.sv:1194:9
		if (reset) begin
			// Trace: ../../rtl/local_mem.sv:1197:13
			reg_val_2_80001008[31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1198:13
			reg_val_2_80001008[63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1199:13
			reg_val_2_80001008[95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1200:13
			reg_val_2_80001008[127-:32] <= 32'h800012fc;
			// Trace: ../../rtl/local_mem.sv:1201:13
			reg_val_2_80001008[159-:32] <= 32'h80001364;
			// Trace: ../../rtl/local_mem.sv:1202:13
			reg_val_2_80001008[191-:32] <= 32'h800013cc;
			// Trace: ../../rtl/local_mem.sv:1203:13
			reg_val_2_80001008[223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1204:13
			reg_val_2_80001008[255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1205:13
			reg_val_2_80001008[287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1206:13
			reg_val_2_80001008[319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1207:13
			reg_val_2_80001008[351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1208:13
			reg_val_2_80001008[383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1209:13
			reg_val_2_80001008[415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1210:13
			reg_val_2_80001008[447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1211:13
			reg_val_2_80001008[479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1212:13
			reg_val_2_80001008[511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1213:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1214:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1215:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1216:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1217:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1218:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1219:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1220:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1221:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1222:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1223:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1224:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1225:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1226:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1227:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1228:13
			reg_val_2_80001008[((0 || 0 ? 16 : 64) * 8) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1229:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1230:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1231:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1232:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1233:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1234:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1235:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1236:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1237:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1238:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1239:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1240:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1241:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000001;
			// Trace: ../../rtl/local_mem.sv:1242:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1243:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'habcd330e;
			// Trace: ../../rtl/local_mem.sv:1244:13
			reg_val_2_80001008[(2 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'he66d1234;
			// Trace: ../../rtl/local_mem.sv:1245:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h0005deec;
			// Trace: ../../rtl/local_mem.sv:1246:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h0000000b;
			// Trace: ../../rtl/local_mem.sv:1247:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1248:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1249:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1250:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1251:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1252:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1253:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1254:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1255:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1256:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1257:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1258:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1259:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1260:13
			reg_val_2_80001008[(3 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1261:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1262:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1263:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1264:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1265:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1266:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1267:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1268:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1269:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1270:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1271:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1272:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1273:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1274:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1275:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1276:13
			reg_val_2_80001008[(4 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1277:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1278:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1279:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1280:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1281:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1282:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1283:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1284:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1285:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1286:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1287:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1288:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1289:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1290:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1291:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1292:13
			reg_val_2_80001008[(5 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1293:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1294:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1295:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1296:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1297:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1298:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1299:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1300:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1301:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1302:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1303:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1304:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1305:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1306:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1307:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1308:13
			reg_val_2_80001008[(6 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1309:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1310:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1311:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1312:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1313:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1314:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1315:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1316:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1317:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1318:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1319:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1320:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1321:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1322:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1323:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1324:13
			reg_val_2_80001008[(7 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1325:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1326:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1327:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1328:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1329:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1330:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1331:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1332:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1333:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1334:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1335:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1336:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1337:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1338:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1339:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1340:13
			reg_val_2_80001008[(8 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1341:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1342:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1343:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1344:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1345:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1346:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1347:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1348:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1349:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1350:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1351:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1352:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1353:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1354:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1355:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1356:13
			reg_val_2_80001008[(9 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1357:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1358:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1359:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1360:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1361:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1362:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1363:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1364:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1365:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1366:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1367:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1368:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1369:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1370:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1371:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1372:13
			reg_val_2_80001008[(10 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1373:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1374:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1375:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1376:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1377:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1378:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1379:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1380:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1381:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1382:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1383:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1384:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1385:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1386:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1387:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1388:13
			reg_val_2_80001008[(11 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1389:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1390:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1391:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1392:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1393:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1394:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1395:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1396:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1397:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1398:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1399:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1400:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1401:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1402:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1403:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1404:13
			reg_val_2_80001008[(12 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1405:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1406:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1407:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1408:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1409:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1410:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1411:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1412:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1413:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1414:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1415:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1416:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1417:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1418:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1419:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1420:13
			reg_val_2_80001008[(13 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1421:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1422:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1423:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1424:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1425:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1426:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1427:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1428:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1429:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1430:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1431:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1432:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1433:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1434:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1435:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1436:13
			reg_val_2_80001008[(14 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1437:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1438:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1439:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1440:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1441:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1442:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1443:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1444:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1445:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1446:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1447:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1448:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1449:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1450:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1451:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1452:13
			reg_val_2_80001008[(15 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1453:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1454:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1455:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1456:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1457:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1458:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1459:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1460:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1461:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1462:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1463:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1464:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1465:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h80001010;
			// Trace: ../../rtl/local_mem.sv:1466:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h80001010;
			// Trace: ../../rtl/local_mem.sv:1468:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1469:13
			reg_val_2_80001008[(16 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1470:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1471:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1472:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1473:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1474:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1475:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1476:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1477:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1478:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1479:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1480:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1481:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1482:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1483:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1484:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1485:13
			reg_val_2_80001008[(17 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1486:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1487:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1488:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1489:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1490:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1491:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1492:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1493:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1494:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1495:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1496:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1497:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1498:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1499:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1500:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1501:13
			reg_val_2_80001008[(18 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1502:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1503:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1504:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1505:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1506:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1507:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1508:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1509:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1510:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1511:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1512:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1513:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1514:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1515:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1516:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1517:13
			reg_val_2_80001008[(19 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1518:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1519:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1520:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1521:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1522:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1523:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1524:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1525:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1526:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1527:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1528:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1529:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1530:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1531:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1532:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1533:13
			reg_val_2_80001008[(20 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1534:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1535:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1536:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1537:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1538:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1539:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1540:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1541:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1542:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1543:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1544:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1545:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1546:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1547:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1548:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1549:13
			reg_val_2_80001008[(21 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1550:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1551:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1552:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1553:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1554:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1555:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1556:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1557:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1558:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1559:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1560:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1561:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1562:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1563:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1564:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1565:13
			reg_val_2_80001008[(22 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1566:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1567:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1568:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1569:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1570:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1571:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1572:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1573:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1574:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1575:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1576:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1577:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1578:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1579:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1580:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1581:13
			reg_val_2_80001008[(23 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1582:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1583:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1584:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1585:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1586:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1587:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1588:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1589:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1590:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1591:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1592:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1593:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1594:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1595:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1596:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1597:13
			reg_val_2_80001008[(24 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1598:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1599:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1600:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1601:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1602:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1603:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1604:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1605:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1606:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1607:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1608:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1609:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1610:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1611:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1612:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1613:13
			reg_val_2_80001008[(25 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1614:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1615:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1616:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1617:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1618:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1619:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1620:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1621:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1622:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1623:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1624:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1625:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1626:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1627:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1628:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1629:13
			reg_val_2_80001008[(26 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1630:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1631:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1632:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1633:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1634:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1635:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1636:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1637:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1638:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1639:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1640:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1641:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1642:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1643:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1644:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1645:13
			reg_val_2_80001008[(27 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1646:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1647:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1648:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1649:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1650:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1651:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1652:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1653:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1654:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1655:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1656:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1657:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1658:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1659:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1660:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1661:13
			reg_val_2_80001008[(28 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1662:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1663:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1664:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1665:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1666:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1667:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1668:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1669:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1670:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1671:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1672:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1673:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1674:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1675:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1676:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1677:13
			reg_val_2_80001008[(29 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1678:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1679:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1680:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1681:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1682:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1683:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1684:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1685:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1686:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1687:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1688:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1689:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1690:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1691:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1692:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1693:13
			reg_val_2_80001008[(30 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1694:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 31-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1695:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 63-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1696:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 95-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1697:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 127-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1698:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 159-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1699:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 191-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1700:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 223-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1701:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 255-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1702:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 287-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1703:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 319-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1704:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 351-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1705:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 383-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1706:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 415-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1707:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 447-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1708:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 479-:32] <= 32'h00000000;
			// Trace: ../../rtl/local_mem.sv:1709:13
			reg_val_2_80001008[(31 * ((0 || 0 ? 16 : 64) * 8)) + 511-:32] <= 32'h00000000;
		end
		else
			// Trace: ../../rtl/local_mem.sv:1713:13
			reg_val_2_80001008 = next_reg_val_2_80001008;
	end
	// Trace: ../../rtl/local_mem.sv:1717:5
	always @(*) begin : WRITE_LOGIC_2_80001008
		// Trace: ../../rtl/local_mem.sv:1719:9
		begin : sv2v_autoblock_3
			// Trace: ../../rtl/local_mem.sv:1719:14
			reg signed [31:0] i;
			// Trace: ../../rtl/local_mem.sv:1719:14
			for (i = 0; i < 32; i = i + 1)
				begin
					// Trace: ../../rtl/local_mem.sv:1721:13
					next_reg_val_2_80001008[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8] = reg_val_2_80001008[i * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8];
				end
		end
		if (wen_2_80001008)
			// Trace: ../../rtl/local_mem.sv:1726:13
			next_reg_val_2_80001008[wsel_2_80001008 * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8] = wdata_2_80001008;
	end
	// Trace: ../../rtl/local_mem.sv:1730:5
	always @(*) begin : READ_LOGIC_2_80001008
		// Trace: ../../rtl/local_mem.sv:1732:9
		rdata_2_80001008 = reg_val_2_80001008[rsel_2_80001008 * ((0 || 0 ? 16 : 64) * 8)+:(0 || 0 ? 16 : 64) * 8];
	end
	// Trace: ../../rtl/local_mem.sv:1736:5
	reg [1:0] chunk_sel;
	// Trace: ../../rtl/local_mem.sv:1739:5
	always @(*) begin : ADDR_HASHING_LOGIC
		// Trace: ../../rtl/local_mem.sv:1741:9
		tb_addr_out_of_bounds = 1'b0;
		// Trace: ../../rtl/local_mem.sv:1744:9
		if (mem_req_addr[(32 - $clog2((0 || 0 ? 16 : 64))) - 20] == 1'b1) begin
			begin
				// Trace: ../../rtl/local_mem.sv:1756:13
				if (mem_req_addr[(32 - $clog2((0 || 0 ? 16 : 64))) - 26] == 1'b0)
					// Trace: ../../rtl/local_mem.sv:1759:17
					chunk_sel = 1;
				else if (mem_req_addr[(32 - $clog2((0 || 0 ? 16 : 64))) - 26] == 1'b0)
					// Trace: ../../rtl/local_mem.sv:1764:17
					chunk_sel = 2;
			end
		end
		else if (mem_req_addr[(32 - $clog2((0 || 0 ? 16 : 64))) - 20] == 1'b0)
			// Trace: ../../rtl/local_mem.sv:1771:13
			chunk_sel = 0;
		else
			// Trace: ../../rtl/local_mem.sv:1776:13
			tb_addr_out_of_bounds = 1'b1;
		// Trace: ../../rtl/local_mem.sv:1781:9
		wsel_0_80000000 = mem_req_addr[5:0];
		// Trace: ../../rtl/local_mem.sv:1782:9
		wdata_0_80000000 = mem_req_data;
		// Trace: ../../rtl/local_mem.sv:1783:9
		rsel_0_80000000 = mem_req_addr[5:0];
		// Trace: ../../rtl/local_mem.sv:1785:9
		wsel_1_80001000 = mem_req_addr[0:0];
		// Trace: ../../rtl/local_mem.sv:1786:9
		wdata_1_80001000 = mem_req_data;
		// Trace: ../../rtl/local_mem.sv:1787:9
		rsel_1_80001000 = mem_req_addr[0:0];
		// Trace: ../../rtl/local_mem.sv:1789:9
		wsel_2_80001008 = mem_req_addr[4:0];
		// Trace: ../../rtl/local_mem.sv:1790:9
		wdata_2_80001008 = mem_req_data;
		// Trace: ../../rtl/local_mem.sv:1791:9
		rsel_2_80001008 = mem_req_addr[4:0];
		// Trace: ../../rtl/local_mem.sv:1794:9
		mem_rsp_data = {16 {32'hdeadbeef}};
		// Trace: ../../rtl/local_mem.sv:1796:9
		wen_0_80000000 = 1'b0;
		// Trace: ../../rtl/local_mem.sv:1797:9
		wen_1_80001000 = 1'b0;
		// Trace: ../../rtl/local_mem.sv:1798:9
		wen_2_80001008 = 1'b0;
		casez (chunk_sel)
			0: begin
				// Trace: ../../rtl/local_mem.sv:1807:17
				wen_0_80000000 = mem_req_rw;
				// Trace: ../../rtl/local_mem.sv:1809:17
				mem_rsp_data = rdata_0_80000000;
			end
			1: begin
				// Trace: ../../rtl/local_mem.sv:1816:17
				wen_1_80001000 = mem_req_rw;
				// Trace: ../../rtl/local_mem.sv:1818:17
				mem_rsp_data = rdata_1_80001000;
			end
			2: begin
				// Trace: ../../rtl/local_mem.sv:1825:17
				wen_2_80001008 = mem_req_rw;
				// Trace: ../../rtl/local_mem.sv:1827:17
				mem_rsp_data = rdata_2_80001008;
			end
			default: begin
				// Trace: ../../rtl/local_mem.sv:1834:17
				mem_rsp_data = {16 {32'hdeadbeef}};
				// Trace: ../../rtl/local_mem.sv:1835:17
				tb_addr_out_of_bounds = 1'b1;
			end
		endcase
	end
	// Trace: ../../rtl/local_mem.sv:1841:5
	always @(*) begin : OTHER_MEM_COMB_LOGIC
		// Trace: ../../rtl/local_mem.sv:1844:9
		mem_rsp_valid = mem_req_valid;
		// Trace: ../../rtl/local_mem.sv:1848:9
		mem_rsp_tag = mem_req_tag;
	end
	// Trace: ../../rtl/local_mem.sv:1852:5
	parameter MEM_REQ_READY_DELAY = 15;
	// Trace: ../../rtl/local_mem.sv:1853:5
	reg [MEM_REQ_READY_DELAY - 1:0] mem_req_ready_reg;
	reg [MEM_REQ_READY_DELAY - 1:0] next_mem_req_ready_reg;
	// Trace: ../../rtl/local_mem.sv:1856:5
	always @(posedge clk) begin : MEM_REQ_READY_REG_LOGIC
		// Trace: ../../rtl/local_mem.sv:1858:9
		if (reset)
			// Trace: ../../rtl/local_mem.sv:1860:13
			mem_req_ready_reg = 1'sb0;
		else
			// Trace: ../../rtl/local_mem.sv:1864:13
			mem_req_ready_reg = next_mem_req_ready_reg;
	end
	// Trace: ../../rtl/local_mem.sv:1869:5
	always @(*) begin : MEM_REQ_READY_DELAY_NEXT_STATE_LOGIC
		// Trace: ../../rtl/local_mem.sv:1871:9
		next_mem_req_ready_reg = {mem_req_ready_reg[MEM_REQ_READY_DELAY - 2:0], 1'b1};
		// Trace: ../../rtl/local_mem.sv:1872:9
		mem_req_ready = mem_req_ready_reg[MEM_REQ_READY_DELAY - 1];
	end
endmodule
module VX_axi_adapter (
	clk,
	reset,
	mem_req_valid,
	mem_req_rw,
	mem_req_byteen,
	mem_req_addr,
	mem_req_data,
	mem_req_tag,
	mem_rsp_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_req_ready,
	m_axi_awid,
	m_axi_awaddr,
	m_axi_awlen,
	m_axi_awsize,
	m_axi_awburst,
	m_axi_awlock,
	m_axi_awcache,
	m_axi_awprot,
	m_axi_awqos,
	m_axi_awvalid,
	m_axi_awready,
	m_axi_wdata,
	m_axi_wstrb,
	m_axi_wlast,
	m_axi_wvalid,
	m_axi_wready,
	m_axi_bid,
	m_axi_bresp,
	m_axi_bvalid,
	m_axi_bready,
	m_axi_arid,
	m_axi_araddr,
	m_axi_arlen,
	m_axi_arsize,
	m_axi_arburst,
	m_axi_arlock,
	m_axi_arcache,
	m_axi_arprot,
	m_axi_arqos,
	m_axi_arvalid,
	m_axi_arready,
	m_axi_rid,
	m_axi_rdata,
	m_axi_rresp,
	m_axi_rlast,
	m_axi_rvalid,
	m_axi_rready
);
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:4:15
	parameter VX_DATA_WIDTH = 512;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:5:15
	parameter VX_ADDR_WIDTH = 32 - $clog2(VX_DATA_WIDTH / 8);
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:6:15
	parameter VX_TAG_WIDTH = 8;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:7:15
	parameter AXI_DATA_WIDTH = VX_DATA_WIDTH;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:8:15
	parameter AXI_ADDR_WIDTH = 32;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:9:15
	parameter AXI_TID_WIDTH = VX_TAG_WIDTH;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:11:15
	parameter VX_BYTEEN_WIDTH = VX_DATA_WIDTH / 8;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:12:15
	parameter AXI_STROBE_WIDTH = AXI_DATA_WIDTH / 8;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:14:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:15:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:18:5
	input wire mem_req_valid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:19:5
	input wire mem_req_rw;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:20:5
	input wire [VX_BYTEEN_WIDTH - 1:0] mem_req_byteen;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:21:5
	input wire [VX_ADDR_WIDTH - 1:0] mem_req_addr;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:22:5
	input wire [VX_DATA_WIDTH - 1:0] mem_req_data;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:23:5
	input wire [VX_TAG_WIDTH - 1:0] mem_req_tag;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:26:5
	input wire mem_rsp_ready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:27:5
	output wire mem_rsp_valid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:28:5
	output wire [VX_DATA_WIDTH - 1:0] mem_rsp_data;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:29:5
	output wire [VX_TAG_WIDTH - 1:0] mem_rsp_tag;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:30:5
	output wire mem_req_ready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:33:5
	output wire [AXI_TID_WIDTH - 1:0] m_axi_awid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:34:5
	output wire [AXI_ADDR_WIDTH - 1:0] m_axi_awaddr;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:35:5
	output wire [7:0] m_axi_awlen;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:36:5
	output wire [2:0] m_axi_awsize;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:37:5
	output wire [1:0] m_axi_awburst;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:38:5
	output wire m_axi_awlock;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:39:5
	output wire [3:0] m_axi_awcache;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:40:5
	output wire [2:0] m_axi_awprot;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:41:5
	output wire [3:0] m_axi_awqos;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:42:5
	output wire m_axi_awvalid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:43:5
	input wire m_axi_awready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:46:5
	output wire [AXI_DATA_WIDTH - 1:0] m_axi_wdata;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:47:5
	output wire [AXI_STROBE_WIDTH - 1:0] m_axi_wstrb;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:48:5
	output wire m_axi_wlast;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:49:5
	output wire m_axi_wvalid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:50:5
	input wire m_axi_wready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:53:5
	input wire [AXI_TID_WIDTH - 1:0] m_axi_bid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:54:5
	input wire [1:0] m_axi_bresp;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:55:5
	input wire m_axi_bvalid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:56:5
	output wire m_axi_bready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:59:5
	output wire [AXI_TID_WIDTH - 1:0] m_axi_arid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:60:5
	output wire [AXI_ADDR_WIDTH - 1:0] m_axi_araddr;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:61:5
	output wire [7:0] m_axi_arlen;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:62:5
	output wire [2:0] m_axi_arsize;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:63:5
	output wire [1:0] m_axi_arburst;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:64:5
	output wire m_axi_arlock;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:65:5
	output wire [3:0] m_axi_arcache;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:66:5
	output wire [2:0] m_axi_arprot;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:67:5
	output wire [3:0] m_axi_arqos;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:68:5
	output wire m_axi_arvalid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:69:5
	input wire m_axi_arready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:72:5
	input wire [AXI_TID_WIDTH - 1:0] m_axi_rid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:73:5
	input wire [AXI_DATA_WIDTH - 1:0] m_axi_rdata;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:74:5
	input wire [1:0] m_axi_rresp;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:75:5
	input wire m_axi_rlast;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:76:5
	input wire m_axi_rvalid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:77:5
	output wire m_axi_rready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:79:5
	localparam AXSIZE = $clog2(VX_DATA_WIDTH / 8);
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:86:5
	reg awvalid_ack;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:87:5
	reg wvalid_ack;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:89:5
	wire mem_req_fire = mem_req_valid && mem_req_ready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:91:5
	always @(posedge clk)
		// Trace: ../../rtl/libs/VX_axi_adapter.sv:92:3
		if (reset) begin
			// Trace: ../../rtl/libs/VX_axi_adapter.sv:93:4
			awvalid_ack <= 0;
			// Trace: ../../rtl/libs/VX_axi_adapter.sv:94:13
			wvalid_ack <= 0;
		end
		else
			// Trace: ../../rtl/libs/VX_axi_adapter.sv:96:13
			if (mem_req_fire) begin
				// Trace: ../../rtl/libs/VX_axi_adapter.sv:97:17
				awvalid_ack <= 0;
				// Trace: ../../rtl/libs/VX_axi_adapter.sv:98:17
				wvalid_ack <= 0;
			end
			else begin
				// Trace: ../../rtl/libs/VX_axi_adapter.sv:100:17
				awvalid_ack <= m_axi_awvalid && m_axi_awready;
				// Trace: ../../rtl/libs/VX_axi_adapter.sv:101:17
				wvalid_ack <= m_axi_wvalid && m_axi_wready;
			end
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:106:5
	wire axi_write_ready = (m_axi_awready || awvalid_ack) && (m_axi_wready || wvalid_ack);
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:109:5
	assign m_axi_awvalid = (mem_req_valid && mem_req_rw) && !awvalid_ack;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:110:5
	assign m_axi_awid = mem_req_tag;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:111:5
	function automatic [AXI_ADDR_WIDTH - 1:0] sv2v_cast_DC0A3;
		input reg [AXI_ADDR_WIDTH - 1:0] inp;
		sv2v_cast_DC0A3 = inp;
	endfunction
	assign m_axi_awaddr = sv2v_cast_DC0A3(mem_req_addr) << AXSIZE;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:112:5
	assign m_axi_awlen = 8'b00000000;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:113:5
	function automatic signed [2:0] sv2v_cast_3_signed;
		input reg signed [2:0] inp;
		sv2v_cast_3_signed = inp;
	endfunction
	assign m_axi_awsize = sv2v_cast_3_signed(AXSIZE);
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:114:5
	assign m_axi_awburst = 2'b00;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:115:5
	assign m_axi_awlock = 1'b0;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:116:5
	assign m_axi_awcache = 4'b0000;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:117:5
	assign m_axi_awprot = 3'b000;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:118:5
	assign m_axi_awqos = 4'b0000;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:121:5
	assign m_axi_wvalid = (mem_req_valid && mem_req_rw) && !wvalid_ack;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:122:5
	assign m_axi_wdata = mem_req_data;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:123:5
	assign m_axi_wstrb = mem_req_byteen;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:124:5
	assign m_axi_wlast = 1'b1;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:129:5
	assign m_axi_bready = 1'b1;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:132:5
	assign m_axi_arvalid = mem_req_valid && !mem_req_rw;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:133:5
	assign m_axi_arid = mem_req_tag;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:134:5
	assign m_axi_araddr = sv2v_cast_DC0A3(mem_req_addr) << AXSIZE;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:135:5
	assign m_axi_arlen = 8'b00000000;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:136:5
	assign m_axi_arsize = sv2v_cast_3_signed(AXSIZE);
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:137:5
	assign m_axi_arburst = 2'b00;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:138:5
	assign m_axi_arlock = 1'b0;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:139:5
	assign m_axi_arcache = 4'b0000;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:140:5
	assign m_axi_arprot = 3'b000;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:141:5
	assign m_axi_arqos = 4'b0000;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:144:5
	assign mem_rsp_valid = m_axi_rvalid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:145:5
	assign mem_rsp_tag = m_axi_rid;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:146:5
	assign mem_rsp_data = m_axi_rdata;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:149:5
	assign m_axi_rready = mem_rsp_ready;
	// Trace: ../../rtl/libs/VX_axi_adapter.sv:152:2
	assign mem_req_ready = (mem_req_rw ? axi_write_ready : m_axi_arready);
endmodule
module VX_bits_insert (
	data_in,
	sel_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_bits_insert.sv:4:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_bits_insert.sv:5:15
	parameter S = 1;
	// Trace: ../../rtl/libs/VX_bits_insert.sv:6:15
	parameter POS = 0;
	// Trace: ../../rtl/libs/VX_bits_insert.sv:8:5
	input wire [N - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_bits_insert.sv:9:5
	input wire [S - 1:0] sel_in;
	// Trace: ../../rtl/libs/VX_bits_insert.sv:10:5
	output wire [(N + S) - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_bits_insert.sv:12:5
	generate
		if (POS == 0) begin : genblk1
			// Trace: ../../rtl/libs/VX_bits_insert.sv:13:9
			assign data_out = {data_in, sel_in};
		end
		else if (POS == N) begin : genblk1
			// Trace: ../../rtl/libs/VX_bits_insert.sv:15:9
			assign data_out = {sel_in, data_in};
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_bits_insert.sv:17:9
			assign data_out = {data_in[N - 1:POS], sel_in, data_in[POS - 1:0]};
		end
	endgenerate
endmodule
module VX_bits_remove (
	data_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_bits_remove.sv:4:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_bits_remove.sv:5:15
	parameter S = 1;
	// Trace: ../../rtl/libs/VX_bits_remove.sv:6:15
	parameter POS = 0;
	// Trace: ../../rtl/libs/VX_bits_remove.sv:8:5
	input wire [N - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_bits_remove.sv:9:5
	output wire [(N - S) - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_bits_remove.sv:13:5
	generate
		if (POS == 0) begin : genblk1
			// Trace: ../../rtl/libs/VX_bits_remove.sv:14:9
			assign data_out = data_in[N - 1:S];
		end
		else if (POS == N) begin : genblk1
			// Trace: ../../rtl/libs/VX_bits_remove.sv:16:9
			assign data_out = data_in[(N - S) - 1:0];
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_bits_remove.sv:18:9
			assign data_out = {data_in[N - 1:POS + S], data_in[POS - 1:0]};
		end
	endgenerate
endmodule
module VX_bypass_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:4:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:5:15
	parameter PASSTHRU = 0;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:7:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:8:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:9:5
	input wire valid_in;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:10:5
	output wire ready_in;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:11:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:12:5
	output wire [DATAW - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:13:5
	input wire ready_out;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:14:5
	output wire valid_out;
	// Trace: ../../rtl/libs/VX_bypass_buffer.sv:16:5
	generate
		if (PASSTHRU) begin : genblk1
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:19:9
			assign ready_in = ready_out;
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:20:9
			assign valid_out = valid_in;
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:21:9
			assign data_out = data_in;
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:23:9
			reg [DATAW - 1:0] buffer;
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:24:9
			reg buffer_valid;
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:26:9
			always @(posedge clk) begin
				// Trace: ../../rtl/libs/VX_bypass_buffer.sv:27:13
				if (reset)
					// Trace: ../../rtl/libs/VX_bypass_buffer.sv:28:17
					buffer_valid <= 0;
				else begin
					// Trace: ../../rtl/libs/VX_bypass_buffer.sv:30:17
					if (ready_out)
						// Trace: ../../rtl/libs/VX_bypass_buffer.sv:31:21
						buffer_valid <= 0;
					if (valid_in && ~ready_out) begin
						// Trace: macro expansion of ASSERT at ../../rtl/libs/VX_bypass_buffer.sv:34:55
						if (!buffer_valid)
							;
						// Trace: ../../rtl/libs/VX_bypass_buffer.sv:35:21
						buffer_valid <= 1;
					end
				end
				if (valid_in && ~ready_out)
					// Trace: ../../rtl/libs/VX_bypass_buffer.sv:40:17
					buffer <= data_in;
			end
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:44:9
			assign ready_in = ready_out || !buffer_valid;
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:45:9
			assign data_out = (buffer_valid ? buffer : data_in);
			// Trace: ../../rtl/libs/VX_bypass_buffer.sv:46:9
			assign valid_out = valid_in || buffer_valid;
		end
	endgenerate
endmodule
module VX_divider (
	clk,
	enable,
	numer,
	denom,
	quotient,
	remainder
);
	// Trace: ../../rtl/libs/VX_divider.sv:5:15
	parameter WIDTHN = 1;
	// Trace: ../../rtl/libs/VX_divider.sv:6:15
	parameter WIDTHD = 1;
	// Trace: ../../rtl/libs/VX_divider.sv:7:15
	parameter WIDTHQ = 1;
	// Trace: ../../rtl/libs/VX_divider.sv:8:15
	parameter WIDTHR = 1;
	// Trace: ../../rtl/libs/VX_divider.sv:9:15
	parameter NSIGNED = 0;
	// Trace: ../../rtl/libs/VX_divider.sv:10:15
	parameter DSIGNED = 0;
	// Trace: ../../rtl/libs/VX_divider.sv:11:15
	parameter LATENCY = 0;
	// Trace: ../../rtl/libs/VX_divider.sv:13:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_divider.sv:14:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_divider.sv:15:5
	input wire [WIDTHN - 1:0] numer;
	// Trace: ../../rtl/libs/VX_divider.sv:16:5
	input wire [WIDTHD - 1:0] denom;
	// Trace: ../../rtl/libs/VX_divider.sv:17:5
	output wire [WIDTHQ - 1:0] quotient;
	// Trace: ../../rtl/libs/VX_divider.sv:18:5
	output wire [WIDTHR - 1:0] remainder;
	// Trace: ../../rtl/libs/VX_divider.sv:49:5
	reg [WIDTHN - 1:0] quotient_unqual;
	// Trace: ../../rtl/libs/VX_divider.sv:50:5
	reg [WIDTHD - 1:0] remainder_unqual;
	// Trace: ../../rtl/libs/VX_divider.sv:52:5
	always @(*) begin
		// Trace: ../../rtl/libs/VX_divider.sv:53:9
		// Trace: ../../rtl/libs/VX_divider.sv:54:13
		if (NSIGNED && DSIGNED) begin
			// Trace: ../../rtl/libs/VX_divider.sv:55:17
			quotient_unqual = $signed(numer) / $signed(denom);
			// Trace: ../../rtl/libs/VX_divider.sv:56:17
			remainder_unqual = $signed(numer) % $signed(denom);
		end
		else if (NSIGNED && !DSIGNED) begin
			// Trace: ../../rtl/libs/VX_divider.sv:59:17
			quotient_unqual = $signed(numer) / denom;
			// Trace: ../../rtl/libs/VX_divider.sv:60:17
			remainder_unqual = $signed(numer) % denom;
		end
		else if (!NSIGNED && DSIGNED) begin
			// Trace: ../../rtl/libs/VX_divider.sv:63:17
			quotient_unqual = numer / $signed(denom);
			// Trace: ../../rtl/libs/VX_divider.sv:64:17
			remainder_unqual = numer % $signed(denom);
		end
		else begin
			// Trace: ../../rtl/libs/VX_divider.sv:67:17
			quotient_unqual = numer / denom;
			// Trace: ../../rtl/libs/VX_divider.sv:68:17
			remainder_unqual = numer % denom;
		end
	end
	// Trace: ../../rtl/libs/VX_divider.sv:73:5
	generate
		if (LATENCY == 0) begin : genblk1
			// Trace: ../../rtl/libs/VX_divider.sv:74:9
			assign quotient = quotient_unqual[WIDTHQ - 1:0];
			// Trace: ../../rtl/libs/VX_divider.sv:75:9
			assign remainder = remainder_unqual[WIDTHR - 1:0];
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_divider.sv:77:9
			reg [WIDTHN - 1:0] quotient_pipe [LATENCY - 1:0];
			// Trace: ../../rtl/libs/VX_divider.sv:78:9
			reg [WIDTHD - 1:0] remainder_pipe [LATENCY - 1:0];
			genvar i;
			for (i = 0; i < LATENCY; i = i + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_divider.sv:81:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_divider.sv:82:17
					if (enable) begin
						// Trace: ../../rtl/libs/VX_divider.sv:83:21
						quotient_pipe[i] <= (0 == i ? quotient_unqual : quotient_pipe[i - 1]);
						// Trace: ../../rtl/libs/VX_divider.sv:84:21
						remainder_pipe[i] <= (0 == i ? remainder_unqual : remainder_pipe[i - 1]);
					end
			end
			// Trace: ../../rtl/libs/VX_divider.sv:89:9
			assign quotient = quotient_pipe[LATENCY - 1][WIDTHQ - 1:0];
			// Trace: ../../rtl/libs/VX_divider.sv:90:9
			assign remainder = remainder_pipe[LATENCY - 1][WIDTHR - 1:0];
		end
	endgenerate
endmodule
module VX_dp_ram (
	clk,
	wren,
	waddr,
	wdata,
	raddr,
	rdata
);
	// Trace: ../../rtl/libs/VX_dp_ram.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:6:15
	parameter SIZE = 1;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:7:15
	parameter BYTEENW = 1;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:8:15
	parameter OUT_REG = 0;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:9:15
	parameter NO_RWCHECK = 0;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:10:15
	parameter LUTRAM = 0;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:11:15
	parameter ADDRW = $clog2(SIZE);
	// Trace: ../../rtl/libs/VX_dp_ram.sv:12:15
	parameter INIT_ENABLE = 0;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:13:15
	parameter INIT_FILE = "";
	// Trace: ../../rtl/libs/VX_dp_ram.sv:14:15
	parameter [DATAW - 1:0] INIT_VALUE = 0;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:16:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:17:5
	input wire [BYTEENW - 1:0] wren;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:18:5
	input wire [ADDRW - 1:0] waddr;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:19:5
	input wire [DATAW - 1:0] wdata;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:20:5
	input wire [ADDRW - 1:0] raddr;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:21:5
	output wire [DATAW - 1:0] rdata;
	// Trace: ../../rtl/libs/VX_dp_ram.sv:38:5
	generate
		if (LUTRAM) begin : genblk1
			if (OUT_REG) begin : genblk1
				// Trace: ../../rtl/libs/VX_dp_ram.sv:40:13
				reg [DATAW - 1:0] rdata_r;
				if (BYTEENW > 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_dp_ram.sv:42:32
					reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:44:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:44:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:44:234
							initial begin : sv2v_autoblock_1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:44:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:44:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:44:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_dp_ram.sv:46:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_dp_ram.sv:47:21
						begin : sv2v_autoblock_2
							// Trace: ../../rtl/libs/VX_dp_ram.sv:47:26
							integer i;
							// Trace: ../../rtl/libs/VX_dp_ram.sv:47:26
							for (i = 0; i < BYTEENW; i = i + 1)
								begin
									// Trace: ../../rtl/libs/VX_dp_ram.sv:48:25
									if (wren[i])
										// Trace: ../../rtl/libs/VX_dp_ram.sv:49:29
										ram[waddr][i * 8+:8] <= wdata[i * 8+:8];
								end
						end
						// Trace: ../../rtl/libs/VX_dp_ram.sv:51:21
						rdata_r <= ram[raddr];
					end
				end
				else begin : genblk1
					// Trace: ../../rtl/libs/VX_dp_ram.sv:54:32
					reg [DATAW - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:56:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:56:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:56:234
							initial begin : sv2v_autoblock_3
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:56:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:56:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:56:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_dp_ram.sv:58:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_dp_ram.sv:59:21
						if (wren)
							// Trace: ../../rtl/libs/VX_dp_ram.sv:60:25
							ram[waddr] <= wdata;
						// Trace: ../../rtl/libs/VX_dp_ram.sv:61:21
						rdata_r <= ram[raddr];
					end
				end
				// Trace: ../../rtl/libs/VX_dp_ram.sv:64:13
				assign rdata = rdata_r;
			end
			else begin : genblk1
				if (BYTEENW > 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_dp_ram.sv:67:32
					reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:69:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:69:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:69:234
							initial begin : sv2v_autoblock_4
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:69:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:69:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:69:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_dp_ram.sv:71:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_dp_ram.sv:72:21
						begin : sv2v_autoblock_5
							// Trace: ../../rtl/libs/VX_dp_ram.sv:72:26
							integer i;
							// Trace: ../../rtl/libs/VX_dp_ram.sv:72:26
							for (i = 0; i < BYTEENW; i = i + 1)
								begin
									// Trace: ../../rtl/libs/VX_dp_ram.sv:73:25
									if (wren[i])
										// Trace: ../../rtl/libs/VX_dp_ram.sv:74:29
										ram[waddr][i * 8+:8] <= wdata[i * 8+:8];
								end
						end
					// Trace: ../../rtl/libs/VX_dp_ram.sv:77:17
					assign rdata = ram[raddr];
				end
				else begin : genblk1
					// Trace: ../../rtl/libs/VX_dp_ram.sv:79:32
					reg [DATAW - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:81:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:81:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:81:234
							initial begin : sv2v_autoblock_6
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:81:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:81:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:81:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_dp_ram.sv:83:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_dp_ram.sv:84:21
						if (wren)
							// Trace: ../../rtl/libs/VX_dp_ram.sv:85:25
							ram[waddr] <= wdata;
					// Trace: ../../rtl/libs/VX_dp_ram.sv:87:17
					assign rdata = ram[raddr];
				end
			end
		end
		else begin : genblk1
			if (OUT_REG) begin : genblk1
				// Trace: ../../rtl/libs/VX_dp_ram.sv:92:13
				reg [DATAW - 1:0] rdata_r;
				if (BYTEENW > 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_dp_ram.sv:95:17
					reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:97:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:97:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:97:234
							initial begin : sv2v_autoblock_7
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:97:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:97:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:97:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_dp_ram.sv:99:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_dp_ram.sv:100:21
						begin : sv2v_autoblock_8
							// Trace: ../../rtl/libs/VX_dp_ram.sv:100:26
							integer i;
							// Trace: ../../rtl/libs/VX_dp_ram.sv:100:26
							for (i = 0; i < BYTEENW; i = i + 1)
								begin
									// Trace: ../../rtl/libs/VX_dp_ram.sv:101:25
									if (wren[i])
										// Trace: ../../rtl/libs/VX_dp_ram.sv:102:29
										ram[waddr][i * 8+:8] <= wdata[i * 8+:8];
								end
						end
						// Trace: ../../rtl/libs/VX_dp_ram.sv:104:21
						rdata_r <= ram[raddr];
					end
				end
				else begin : genblk1
					// Trace: ../../rtl/libs/VX_dp_ram.sv:107:17
					reg [DATAW - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:109:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:109:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:109:234
							initial begin : sv2v_autoblock_9
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:109:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:109:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:109:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_dp_ram.sv:111:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_dp_ram.sv:112:21
						if (wren)
							// Trace: ../../rtl/libs/VX_dp_ram.sv:113:25
							ram[waddr] <= wdata;
						// Trace: ../../rtl/libs/VX_dp_ram.sv:114:21
						rdata_r <= ram[raddr];
					end
				end
				// Trace: ../../rtl/libs/VX_dp_ram.sv:117:13
				assign rdata = rdata_r;
			end
			else begin : genblk1
				if (NO_RWCHECK) begin : genblk1
					if (BYTEENW > 1) begin : genblk1
						// Trace: ../../rtl/libs/VX_dp_ram.sv:121:38
						reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
						if (INIT_ENABLE) begin : genblk1
							if (INIT_FILE != "") begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:123:136
								initial begin
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:123:144
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:123:238
								initial begin : sv2v_autoblock_10
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:123:298
									integer i;
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:123:298
									for (i = 0; i < SIZE; i = i + 1)
										begin
											// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:123:348
											ram[i] = INIT_VALUE;
										end
								end
							end
						end
						// Trace: ../../rtl/libs/VX_dp_ram.sv:125:21
						always @(posedge clk)
							// Trace: ../../rtl/libs/VX_dp_ram.sv:126:25
							begin : sv2v_autoblock_11
								// Trace: ../../rtl/libs/VX_dp_ram.sv:126:30
								integer i;
								// Trace: ../../rtl/libs/VX_dp_ram.sv:126:30
								for (i = 0; i < BYTEENW; i = i + 1)
									begin
										// Trace: ../../rtl/libs/VX_dp_ram.sv:127:29
										if (wren[i])
											// Trace: ../../rtl/libs/VX_dp_ram.sv:128:33
											ram[waddr][i * 8+:8] <= wdata[i * 8+:8];
									end
							end
						// Trace: ../../rtl/libs/VX_dp_ram.sv:131:21
						assign rdata = ram[raddr];
					end
					else begin : genblk1
						// Trace: ../../rtl/libs/VX_dp_ram.sv:133:38
						reg [DATAW - 1:0] ram [SIZE - 1:0];
						if (INIT_ENABLE) begin : genblk1
							if (INIT_FILE != "") begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:135:136
								initial begin
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:135:144
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:135:238
								initial begin : sv2v_autoblock_12
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:135:298
									integer i;
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:135:298
									for (i = 0; i < SIZE; i = i + 1)
										begin
											// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:135:348
											ram[i] = INIT_VALUE;
										end
								end
							end
						end
						// Trace: ../../rtl/libs/VX_dp_ram.sv:137:21
						always @(posedge clk)
							// Trace: ../../rtl/libs/VX_dp_ram.sv:138:25
							if (wren)
								// Trace: ../../rtl/libs/VX_dp_ram.sv:139:29
								ram[waddr] <= wdata;
						// Trace: ../../rtl/libs/VX_dp_ram.sv:141:21
						assign rdata = ram[raddr];
					end
				end
				else begin : genblk1
					if (BYTEENW > 1) begin : genblk1
						// Trace: ../../rtl/libs/VX_dp_ram.sv:145:21
						reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
						if (INIT_ENABLE) begin : genblk1
							if (INIT_FILE != "") begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:147:136
								initial begin
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:147:144
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:147:238
								initial begin : sv2v_autoblock_13
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:147:298
									integer i;
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:147:298
									for (i = 0; i < SIZE; i = i + 1)
										begin
											// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:147:348
											ram[i] = INIT_VALUE;
										end
								end
							end
						end
						// Trace: ../../rtl/libs/VX_dp_ram.sv:149:21
						always @(posedge clk)
							// Trace: ../../rtl/libs/VX_dp_ram.sv:150:25
							begin : sv2v_autoblock_14
								// Trace: ../../rtl/libs/VX_dp_ram.sv:150:30
								integer i;
								// Trace: ../../rtl/libs/VX_dp_ram.sv:150:30
								for (i = 0; i < BYTEENW; i = i + 1)
									begin
										// Trace: ../../rtl/libs/VX_dp_ram.sv:151:29
										if (wren[i])
											// Trace: ../../rtl/libs/VX_dp_ram.sv:152:33
											ram[waddr][i * 8+:8] <= wdata[i * 8+:8];
									end
							end
						// Trace: ../../rtl/libs/VX_dp_ram.sv:155:21
						assign rdata = ram[raddr];
					end
					else begin : genblk1
						// Trace: ../../rtl/libs/VX_dp_ram.sv:157:21
						reg [DATAW - 1:0] ram [SIZE - 1:0];
						if (INIT_ENABLE) begin : genblk1
							if (INIT_FILE != "") begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:159:136
								initial begin
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:159:144
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:159:238
								initial begin : sv2v_autoblock_15
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:159:298
									integer i;
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:159:298
									for (i = 0; i < SIZE; i = i + 1)
										begin
											// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_dp_ram.sv:159:348
											ram[i] = INIT_VALUE;
										end
								end
							end
						end
						// Trace: ../../rtl/libs/VX_dp_ram.sv:161:21
						always @(posedge clk)
							// Trace: ../../rtl/libs/VX_dp_ram.sv:162:25
							if (wren)
								// Trace: ../../rtl/libs/VX_dp_ram.sv:163:29
								ram[waddr] <= wdata;
						// Trace: ../../rtl/libs/VX_dp_ram.sv:165:21
						assign rdata = ram[raddr];
					end
				end
			end
		end
	endgenerate
endmodule
module VX_elastic_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:6:15
	parameter SIZE = 2;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:7:15
	parameter OUT_REG = 0;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:8:15
	parameter LUTRAM = 0;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:10:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:11:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:13:5
	input wire valid_in;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:14:5
	output wire ready_in;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:15:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:17:5
	output wire [DATAW - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:18:5
	input wire ready_out;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:19:5
	output wire valid_out;
	// Trace: ../../rtl/libs/VX_elastic_buffer.sv:23:5
	generate
		if (SIZE == 0) begin : genblk1
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:28:9
			assign valid_out = valid_in;
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:29:9
			assign data_out = data_in;
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:30:9
			assign ready_in = ready_out;
		end
		else if (SIZE == 2) begin : genblk1
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:34:9
			VX_skid_buffer #(
				.DATAW(DATAW),
				.OUT_REG(OUT_REG)
			) queue(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.data_in(data_in),
				.ready_in(ready_in),
				.valid_out(valid_out),
				.data_out(data_out),
				.ready_out(ready_out)
			);
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:50:9
			wire empty;
			wire full;
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:52:9
			wire push = valid_in && ready_in;
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:53:9
			wire pop = valid_out && ready_out;
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:55:9
			VX_fifo_queue #(
				.DATAW(DATAW),
				.SIZE(SIZE),
				.OUT_REG(OUT_REG),
				.LUTRAM(LUTRAM)
			) queue(
				.clk(clk),
				.reset(reset),
				.push(push),
				.pop(pop),
				.data_in(data_in),
				.data_out(data_out),
				.empty(empty),
				.full(full)
			);
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:74:9
			assign ready_in = ~full;
			// Trace: ../../rtl/libs/VX_elastic_buffer.sv:75:9
			assign valid_out = ~empty;
		end
	endgenerate
endmodule
module VX_fair_arbiter (
	clk,
	reset,
	enable,
	requests,
	grant_index,
	grant_onehot,
	grant_valid
);
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:5:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:6:15
	parameter LOCK_ENABLE = 0;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:7:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:9:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:10:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:11:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:12:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:13:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:14:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:15:5
	output wire grant_valid;
	// Trace: ../../rtl/libs/VX_fair_arbiter.sv:18:5
	generate
		if (NUM_REQS == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:22:9
			assign grant_index = 0;
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:23:9
			assign grant_onehot = requests;
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:24:9
			assign grant_valid = requests[0];
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:28:9
			reg [NUM_REQS - 1:0] buffer;
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:29:9
			reg use_buffer;
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:31:9
			wire [NUM_REQS - 1:0] requests_qual = (use_buffer ? buffer : requests);
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:32:9
			wire [NUM_REQS - 1:0] buffer_n = requests_qual & ~grant_onehot;
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:34:9
			always @(posedge clk) begin
				// Trace: ../../rtl/libs/VX_fair_arbiter.sv:35:13
				if (reset)
					// Trace: ../../rtl/libs/VX_fair_arbiter.sv:36:17
					use_buffer <= 0;
				else if (!LOCK_ENABLE || enable)
					// Trace: ../../rtl/libs/VX_fair_arbiter.sv:38:17
					use_buffer <= buffer_n != 0;
				if (!LOCK_ENABLE || enable)
					// Trace: ../../rtl/libs/VX_fair_arbiter.sv:41:17
					buffer <= buffer_n;
			end
			// Trace: ../../rtl/libs/VX_fair_arbiter.sv:45:9
			VX_fixed_arbiter #(
				.NUM_REQS(NUM_REQS),
				.LOCK_ENABLE(LOCK_ENABLE)
			) fixed_arbiter(
				.clk(clk),
				.reset(reset),
				.enable(enable),
				.requests(requests_qual),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot),
				.grant_valid(grant_valid)
			);
		end
	endgenerate
endmodule
module VX_fifo_queue (
	clk,
	reset,
	push,
	pop,
	data_in,
	data_out,
	empty,
	alm_empty,
	full,
	alm_full,
	size
);
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:6:15
	parameter SIZE = 2;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:7:15
	parameter ALM_FULL = SIZE - 1;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:8:15
	parameter ALM_EMPTY = 1;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:9:15
	parameter ADDRW = $clog2(SIZE);
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:10:15
	parameter SIZEW = $clog2(SIZE + 1);
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:11:15
	parameter OUT_REG = 0;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:12:15
	parameter LUTRAM = 1;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:14:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:15:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:16:5
	input wire push;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:17:5
	input wire pop;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:18:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:19:5
	output wire [DATAW - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:20:5
	output wire empty;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:21:5
	output wire alm_empty;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:22:5
	output wire full;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:23:5
	output wire alm_full;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:24:5
	output wire [SIZEW - 1:0] size;
	// Trace: ../../rtl/libs/VX_fifo_queue.sv:28:5
	function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
		input reg signed [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D_signed = inp;
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	function automatic [ADDRW - 1:0] sv2v_cast_8BB5D;
		input reg [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D = inp;
	endfunction
	generate
		if (SIZE == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:30:9
			reg [DATAW - 1:0] head_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:31:9
			reg size_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:33:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_fifo_queue.sv:34:13
				if (reset) begin
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:35:17
					head_r <= 0;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:36:17
					size_r <= 0;
				end
				else begin
					// Trace: macro expansion of ASSERT at ../../rtl/libs/VX_fifo_queue.sv:38:52
					if (!push || !full)
						;
					if (!pop || !empty)
						;
					if (push) begin
						begin
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:41:21
							if (!pop)
								// Trace: ../../rtl/libs/VX_fifo_queue.sv:42:25
								size_r <= 1;
						end
					end
					else if (pop)
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:45:21
						size_r <= 0;
					if (push)
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:48:21
						head_r <= data_in;
				end
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:53:9
			assign data_out = head_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:54:9
			assign empty = size_r == 0;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:55:9
			assign alm_empty = 1'b1;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:56:9
			assign full = size_r != 0;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:57:9
			assign alm_full = 1'b1;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:58:9
			assign size = size_r;
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:62:9
			reg empty_r;
			reg alm_empty_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:63:9
			reg full_r;
			reg alm_full_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:64:9
			reg [ADDRW - 1:0] used_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:66:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_fifo_queue.sv:67:13
				if (reset) begin
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:68:17
					empty_r <= 1;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:69:17
					alm_empty_r <= 1;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:70:17
					full_r <= 0;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:71:17
					alm_full_r <= 0;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:72:17
					used_r <= 0;
				end
				else begin
					// Trace: macro expansion of ASSERT at ../../rtl/libs/VX_fifo_queue.sv:74:52
					if (!push || !full)
						;
					if (!pop || !empty)
						;
					if (push) begin
						begin
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:77:21
							if (!pop) begin
								// Trace: ../../rtl/libs/VX_fifo_queue.sv:78:25
								empty_r <= 0;
								// Trace: ../../rtl/libs/VX_fifo_queue.sv:79:25
								if (used_r == sv2v_cast_8BB5D_signed(ALM_EMPTY))
									// Trace: ../../rtl/libs/VX_fifo_queue.sv:80:29
									alm_empty_r <= 0;
								if (used_r == sv2v_cast_8BB5D_signed(SIZE - 1))
									// Trace: ../../rtl/libs/VX_fifo_queue.sv:82:29
									full_r <= 1;
								if (used_r == sv2v_cast_8BB5D_signed(ALM_FULL - 1))
									// Trace: ../../rtl/libs/VX_fifo_queue.sv:84:29
									alm_full_r <= 1;
							end
						end
					end
					else if (pop) begin
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:87:21
						full_r <= 0;
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:88:21
						if (used_r == sv2v_cast_8BB5D_signed(ALM_FULL))
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:89:25
							alm_full_r <= 0;
						if (used_r == sv2v_cast_8BB5D_signed(1))
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:91:25
							empty_r <= 1;
						if (used_r == sv2v_cast_8BB5D_signed(ALM_EMPTY + 1))
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:93:25
							alm_empty_r <= 1;
					end
					if (SIZE > 2)
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:96:21
						used_r <= used_r + sv2v_cast_8BB5D_signed($signed(sv2v_cast_2(push) - sv2v_cast_2(pop)));
					else
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:99:21
						used_r[0] <= used_r[0] ^ (push ^ pop);
				end
			if (SIZE == 2) begin : genblk1
				if (0 == OUT_REG) begin : genblk1
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:108:17
					reg [DATAW - 1:0] shift_reg [1:0];
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:110:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:111:21
						if (push) begin
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:112:25
							shift_reg[1] <= shift_reg[0];
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:113:25
							shift_reg[0] <= data_in;
						end
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:117:17
					assign data_out = shift_reg[!used_r[0]];
				end
				else begin : genblk1
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:121:17
					reg [DATAW - 1:0] data_out_r;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:122:17
					reg [DATAW - 1:0] buffer;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:124:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:125:21
						if (push)
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:126:25
							buffer <= data_in;
						if (push && (empty_r || (used_r && pop)))
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:129:25
							data_out_r <= data_in;
						else if (pop)
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:131:25
							data_out_r <= buffer;
					end
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:135:17
					assign data_out = data_out_r;
				end
			end
			else begin : genblk1
				if (0 == OUT_REG) begin : genblk1
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:143:17
					reg [ADDRW - 1:0] rd_ptr_r;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:144:17
					reg [ADDRW - 1:0] wr_ptr_r;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:146:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:147:21
						if (reset) begin
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:148:25
							rd_ptr_r <= 0;
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:149:25
							wr_ptr_r <= 0;
						end
						else begin
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:151:25
							wr_ptr_r <= wr_ptr_r + sv2v_cast_8BB5D(push);
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:152:25
							rd_ptr_r <= rd_ptr_r + sv2v_cast_8BB5D(pop);
						end
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:156:17
					VX_dp_ram #(
						.DATAW(DATAW),
						.SIZE(SIZE),
						.OUT_REG(0),
						.LUTRAM(LUTRAM)
					) dp_ram(
						.clk(clk),
						.wren(push),
						.waddr(wr_ptr_r),
						.wdata(data_in),
						.raddr(rd_ptr_r),
						.rdata(data_out)
					);
				end
				else begin : genblk1
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:172:17
					wire [DATAW - 1:0] dout;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:173:17
					reg [DATAW - 1:0] dout_r;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:174:17
					reg [ADDRW - 1:0] wr_ptr_r;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:175:17
					reg [ADDRW - 1:0] rd_ptr_r;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:176:17
					reg [ADDRW - 1:0] rd_ptr_n_r;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:178:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:179:21
						if (reset) begin
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:180:25
							wr_ptr_r <= 0;
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:181:25
							rd_ptr_r <= 0;
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:182:25
							rd_ptr_n_r <= 1;
						end
						else begin
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:184:25
							if (push)
								// Trace: ../../rtl/libs/VX_fifo_queue.sv:185:29
								wr_ptr_r <= wr_ptr_r + sv2v_cast_8BB5D_signed(1);
							if (pop) begin
								// Trace: ../../rtl/libs/VX_fifo_queue.sv:188:29
								rd_ptr_r <= rd_ptr_n_r;
								// Trace: ../../rtl/libs/VX_fifo_queue.sv:189:29
								if (SIZE > 2)
									// Trace: ../../rtl/libs/VX_fifo_queue.sv:190:33
									rd_ptr_n_r <= rd_ptr_r + sv2v_cast_8BB5D_signed(2);
								else
									// Trace: ../../rtl/libs/VX_fifo_queue.sv:192:33
									rd_ptr_n_r <= ~rd_ptr_n_r;
							end
						end
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:198:17
					VX_dp_ram #(
						.DATAW(DATAW),
						.SIZE(SIZE),
						.OUT_REG(0),
						.LUTRAM(LUTRAM)
					) dp_ram(
						.clk(clk),
						.wren(push),
						.waddr(wr_ptr_r),
						.wdata(data_in),
						.raddr(rd_ptr_n_r),
						.rdata(dout)
					);
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:212:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_fifo_queue.sv:213:21
						if (push && (empty_r || ((used_r == sv2v_cast_8BB5D_signed(1)) && pop)))
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:214:25
							dout_r <= data_in;
						else if (pop)
							// Trace: ../../rtl/libs/VX_fifo_queue.sv:216:25
							dout_r <= dout;
					// Trace: ../../rtl/libs/VX_fifo_queue.sv:220:17
					assign data_out = dout_r;
				end
			end
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:224:9
			assign empty = empty_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:225:9
			assign alm_empty = alm_empty_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:226:9
			assign full = full_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:227:9
			assign alm_full = alm_full_r;
			// Trace: ../../rtl/libs/VX_fifo_queue.sv:228:9
			assign size = {full_r, used_r};
		end
	endgenerate
endmodule
module VX_find_first (
	data_i,
	valid_i,
	data_o,
	valid_o
);
	// Trace: ../../rtl/libs/VX_find_first.sv:5:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_find_first.sv:6:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_find_first.sv:7:15
	parameter REVERSE = 0;
	// Trace: ../../rtl/libs/VX_find_first.sv:8:15
	parameter LOGN = $clog2(N);
	// Trace: ../../rtl/libs/VX_find_first.sv:10:5
	input wire [(N * DATAW) - 1:0] data_i;
	// Trace: ../../rtl/libs/VX_find_first.sv:11:5
	input wire [N - 1:0] valid_i;
	// Trace: ../../rtl/libs/VX_find_first.sv:12:5
	output wire [DATAW - 1:0] data_o;
	// Trace: ../../rtl/libs/VX_find_first.sv:13:5
	output wire valid_o;
	// Trace: ../../rtl/libs/VX_find_first.sv:15:5
	localparam TL = (1 << LOGN) - 1;
	// Trace: ../../rtl/libs/VX_find_first.sv:16:5
	localparam TN = (1 << (LOGN + 1)) - 1;
	// Trace: ../../rtl/libs/VX_find_first.sv:19:5
	wire [TN - 1:0] s_n;
	// Trace: ../../rtl/libs/VX_find_first.sv:20:5
	wire [(TN * DATAW) - 1:0] d_n;
	// Trace: ../../rtl/libs/VX_find_first.sv:23:5
	genvar i;
	generate
		for (i = 0; i < N; i = i + 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_find_first.sv:24:9
			assign s_n[TL + i] = (REVERSE ? valid_i[(N - 1) - i] : valid_i[i]);
			// Trace: ../../rtl/libs/VX_find_first.sv:25:9
			assign d_n[(TL + i) * DATAW+:DATAW] = (REVERSE ? data_i[((N - 1) - i) * DATAW+:DATAW] : data_i[i * DATAW+:DATAW]);
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_find_first.sv:28:5
	generate
		for (i = TL + N; i < TN; i = i + 1) begin : genblk2
			// Trace: ../../rtl/libs/VX_find_first.sv:29:9
			assign s_n[i] = 0;
			// Trace: ../../rtl/libs/VX_find_first.sv:30:9
			assign d_n[i * DATAW+:DATAW] = 1'sbx;
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_find_first.sv:33:5
	genvar j;
	generate
		for (j = 0; j < LOGN; j = j + 1) begin : genblk3
			genvar i;
			for (i = 0; i < (2 ** j); i = i + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_find_first.sv:35:13
				assign s_n[((2 ** j) - 1) + i] = s_n[((2 ** (j + 1)) - 1) + (i * 2)] | s_n[(((2 ** (j + 1)) - 1) + (i * 2)) + 1];
				// Trace: ../../rtl/libs/VX_find_first.sv:36:13
				assign d_n[(((2 ** j) - 1) + i) * DATAW+:DATAW] = (s_n[((2 ** (j + 1)) - 1) + (i * 2)] ? d_n[(((2 ** (j + 1)) - 1) + (i * 2)) * DATAW+:DATAW] : d_n[((((2 ** (j + 1)) - 1) + (i * 2)) + 1) * DATAW+:DATAW]);
			end
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_find_first.sv:40:5
	assign valid_o = s_n[0];
	// Trace: ../../rtl/libs/VX_find_first.sv:41:5
	assign data_o = d_n[0+:DATAW];
endmodule
module VX_fixed_arbiter (
	clk,
	reset,
	requests,
	enable,
	grant_index,
	grant_onehot,
	grant_valid
);
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:5:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:6:15
	parameter LOCK_ENABLE = 0;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:7:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:9:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:10:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:11:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:12:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:13:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:14:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:15:5
	output wire grant_valid;
	// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:23:5
	generate
		if (NUM_REQS == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:25:9
			assign grant_index = 0;
			// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:26:9
			assign grant_onehot = requests;
			// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:27:9
			assign grant_valid = requests[0];
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_fixed_arbiter.sv:31:9
			VX_priority_encoder #(.N(NUM_REQS)) tid_select(
				.data_in(requests),
				.index(grant_index),
				.onehot(grant_onehot),
				.valid_out(grant_valid)
			);
		end
	endgenerate
endmodule
module VX_index_buffer (
	clk,
	reset,
	write_addr,
	write_data,
	acquire_slot,
	read_addr,
	read_data,
	release_addr,
	release_slot,
	empty,
	full
);
	// Trace: ../../rtl/libs/VX_index_buffer.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:6:15
	parameter SIZE = 1;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:7:15
	parameter LUTRAM = 1;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:8:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: ../../rtl/libs/VX_index_buffer.sv:10:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:11:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:13:5
	output wire [ADDRW - 1:0] write_addr;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:14:5
	input wire [DATAW - 1:0] write_data;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:15:5
	input wire acquire_slot;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:17:5
	input wire [ADDRW - 1:0] read_addr;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:18:5
	output wire [DATAW - 1:0] read_data;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:19:5
	input wire [ADDRW - 1:0] release_addr;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:20:5
	input wire release_slot;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:22:5
	output wire empty;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:23:5
	output wire full;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:25:5
	reg [SIZE - 1:0] free_slots;
	reg [SIZE - 1:0] free_slots_n;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:26:5
	reg [ADDRW - 1:0] write_addr_r;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:27:5
	reg empty_r;
	reg full_r;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:29:5
	wire free_valid;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:30:5
	wire [ADDRW - 1:0] free_index;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:32:5
	VX_lzc #(.N(SIZE)) free_slots_sel(
		.in_i(free_slots_n),
		.cnt_o(free_index),
		.valid_o(free_valid)
	);
	// Trace: ../../rtl/libs/VX_index_buffer.sv:40:5
	always @(*) begin
		// Trace: ../../rtl/libs/VX_index_buffer.sv:41:9
		free_slots_n = free_slots;
		// Trace: ../../rtl/libs/VX_index_buffer.sv:42:9
		if (release_slot)
			// Trace: ../../rtl/libs/VX_index_buffer.sv:43:13
			free_slots_n[release_addr] = 1;
		if (acquire_slot)
			// Trace: ../../rtl/libs/VX_index_buffer.sv:46:13
			free_slots_n[write_addr_r] = 0;
	end
	// Trace: ../../rtl/libs/VX_index_buffer.sv:50:5
	function automatic [ADDRW - 1:0] sv2v_cast_8BB5D;
		input reg [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D = inp;
	endfunction
	always @(posedge clk)
		// Trace: ../../rtl/libs/VX_index_buffer.sv:51:9
		if (reset) begin
			// Trace: ../../rtl/libs/VX_index_buffer.sv:52:13
			write_addr_r <= sv2v_cast_8BB5D(1'b0);
			// Trace: ../../rtl/libs/VX_index_buffer.sv:53:13
			free_slots <= {SIZE {1'b1}};
			// Trace: ../../rtl/libs/VX_index_buffer.sv:54:13
			empty_r <= 1'b1;
			// Trace: ../../rtl/libs/VX_index_buffer.sv:55:13
			full_r <= 1'b0;
		end
		else begin
			// Trace: ../../rtl/libs/VX_index_buffer.sv:57:13
			if (release_slot)
				// Trace: macro expansion of ASSERT at ../../rtl/libs/VX_index_buffer.sv:58:112
				if (0 == free_slots[release_addr])
					;
			if (acquire_slot)
				// Trace: macro expansion of ASSERT at ../../rtl/libs/VX_index_buffer.sv:61:105
				if (1 == free_slots[write_addr])
					;
			// Trace: ../../rtl/libs/VX_index_buffer.sv:63:13
			write_addr_r <= free_index;
			// Trace: ../../rtl/libs/VX_index_buffer.sv:64:13
			free_slots <= free_slots_n;
			// Trace: ../../rtl/libs/VX_index_buffer.sv:65:13
			empty_r <= &free_slots_n;
			// Trace: ../../rtl/libs/VX_index_buffer.sv:66:13
			full_r <= ~free_valid;
		end
	// Trace: ../../rtl/libs/VX_index_buffer.sv:70:5
	VX_dp_ram #(
		.DATAW(DATAW),
		.SIZE(SIZE),
		.LUTRAM(LUTRAM)
	) data_table(
		.clk(clk),
		.wren(acquire_slot),
		.waddr(write_addr_r),
		.wdata(write_data),
		.raddr(read_addr),
		.rdata(read_data)
	);
	// Trace: ../../rtl/libs/VX_index_buffer.sv:83:5
	assign write_addr = write_addr_r;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:84:5
	assign empty = empty_r;
	// Trace: ../../rtl/libs/VX_index_buffer.sv:85:5
	assign full = full_r;
endmodule
module VX_index_queue (
	clk,
	reset,
	write_data,
	write_addr,
	push,
	pop,
	full,
	empty,
	read_addr,
	read_data
);
	// Trace: ../../rtl/libs/VX_index_queue.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_index_queue.sv:6:15
	parameter SIZE = 1;
	// Trace: ../../rtl/libs/VX_index_queue.sv:8:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_index_queue.sv:9:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_index_queue.sv:10:5
	input wire [DATAW - 1:0] write_data;
	// Trace: ../../rtl/libs/VX_index_queue.sv:11:5
	output wire [(SIZE > 1 ? $clog2(SIZE) : 1) - 1:0] write_addr;
	// Trace: ../../rtl/libs/VX_index_queue.sv:12:5
	input wire push;
	// Trace: ../../rtl/libs/VX_index_queue.sv:13:5
	input wire pop;
	// Trace: ../../rtl/libs/VX_index_queue.sv:14:5
	output wire full;
	// Trace: ../../rtl/libs/VX_index_queue.sv:15:5
	output wire empty;
	// Trace: ../../rtl/libs/VX_index_queue.sv:16:5
	input wire [(SIZE > 1 ? $clog2(SIZE) : 1) - 1:0] read_addr;
	// Trace: ../../rtl/libs/VX_index_queue.sv:17:5
	output wire [DATAW - 1:0] read_data;
	// Trace: ../../rtl/libs/VX_index_queue.sv:19:5
	reg [DATAW - 1:0] entries [SIZE - 1:0];
	// Trace: ../../rtl/libs/VX_index_queue.sv:20:5
	reg [SIZE - 1:0] valid;
	// Trace: ../../rtl/libs/VX_index_queue.sv:21:5
	reg [(SIZE > 1 ? $clog2(SIZE) : 1):0] rd_ptr;
	reg [(SIZE > 1 ? $clog2(SIZE) : 1):0] wr_ptr;
	// Trace: ../../rtl/libs/VX_index_queue.sv:23:5
	wire [(SIZE > 1 ? $clog2(SIZE) : 1) - 1:0] rd_a;
	wire [(SIZE > 1 ? $clog2(SIZE) : 1) - 1:0] wr_a;
	// Trace: ../../rtl/libs/VX_index_queue.sv:24:5
	wire enqueue;
	wire dequeue;
	// Trace: ../../rtl/libs/VX_index_queue.sv:26:5
	assign rd_a = rd_ptr[(SIZE > 1 ? $clog2(SIZE) : 1) - 1:0];
	// Trace: ../../rtl/libs/VX_index_queue.sv:27:5
	assign wr_a = wr_ptr[(SIZE > 1 ? $clog2(SIZE) : 1) - 1:0];
	// Trace: ../../rtl/libs/VX_index_queue.sv:29:5
	assign empty = wr_ptr == rd_ptr;
	// Trace: ../../rtl/libs/VX_index_queue.sv:30:5
	assign full = (wr_a == rd_a) && (wr_ptr[(SIZE > 1 ? $clog2(SIZE) : 1)] != rd_ptr[(SIZE > 1 ? $clog2(SIZE) : 1)]);
	// Trace: ../../rtl/libs/VX_index_queue.sv:32:5
	assign enqueue = push;
	// Trace: ../../rtl/libs/VX_index_queue.sv:33:5
	assign dequeue = !empty && !valid[rd_a];
	// Trace: ../../rtl/libs/VX_index_queue.sv:37:5
	always @(posedge clk) begin
		// Trace: ../../rtl/libs/VX_index_queue.sv:38:9
		if (reset) begin
			// Trace: ../../rtl/libs/VX_index_queue.sv:39:13
			rd_ptr <= 0;
			// Trace: ../../rtl/libs/VX_index_queue.sv:40:13
			wr_ptr <= 0;
			// Trace: ../../rtl/libs/VX_index_queue.sv:41:13
			valid <= 0;
		end
		else begin
			// Trace: ../../rtl/libs/VX_index_queue.sv:43:13
			if (enqueue) begin
				// Trace: ../../rtl/libs/VX_index_queue.sv:44:17
				valid[wr_a] <= 1;
				// Trace: ../../rtl/libs/VX_index_queue.sv:45:17
				wr_ptr <= wr_ptr + 1;
			end
			if (dequeue)
				// Trace: ../../rtl/libs/VX_index_queue.sv:48:17
				rd_ptr <= rd_ptr + 1;
			if (pop)
				// Trace: ../../rtl/libs/VX_index_queue.sv:51:17
				valid[read_addr] <= 0;
		end
		if (enqueue)
			// Trace: ../../rtl/libs/VX_index_queue.sv:56:13
			entries[wr_a] <= write_data;
	end
	// Trace: ../../rtl/libs/VX_index_queue.sv:60:5
	assign write_addr = wr_a;
	// Trace: ../../rtl/libs/VX_index_queue.sv:61:5
	assign read_data = entries[read_addr];
endmodule
module VX_lzc (
	in_i,
	cnt_o,
	valid_o
);
	// Trace: ../../rtl/libs/VX_lzc.sv:5:15
	parameter N = 2;
	// Trace: ../../rtl/libs/VX_lzc.sv:6:15
	parameter MODE = 0;
	// Trace: ../../rtl/libs/VX_lzc.sv:7:15
	parameter LOGN = $clog2(N);
	// Trace: ../../rtl/libs/VX_lzc.sv:9:5
	input wire [N - 1:0] in_i;
	// Trace: ../../rtl/libs/VX_lzc.sv:10:5
	output wire [LOGN - 1:0] cnt_o;
	// Trace: ../../rtl/libs/VX_lzc.sv:11:5
	output wire valid_o;
	// Trace: ../../rtl/libs/VX_lzc.sv:13:5
	wire [(N * LOGN) - 1:0] indices;
	// Trace: ../../rtl/libs/VX_lzc.sv:15:5
	genvar i;
	function automatic signed [LOGN - 1:0] sv2v_cast_B9644_signed;
		input reg signed [LOGN - 1:0] inp;
		sv2v_cast_B9644_signed = inp;
	endfunction
	generate
		for (i = 0; i < N; i = i + 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_lzc.sv:16:9
			assign indices[i * LOGN+:LOGN] = (MODE ? sv2v_cast_B9644_signed((N - 1) - i) : sv2v_cast_B9644_signed(i));
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_lzc.sv:19:5
	VX_find_first #(
		.N(N),
		.DATAW(LOGN),
		.REVERSE(MODE)
	) find_first(
		.data_i(indices),
		.valid_i(in_i),
		.data_o(cnt_o),
		.valid_o(valid_o)
	);
endmodule
module VX_matrix_arbiter (
	clk,
	reset,
	enable,
	requests,
	grant_index,
	grant_onehot,
	grant_valid
);
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:5:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:6:15
	parameter LOCK_ENABLE = 0;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:7:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:9:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:10:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:11:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:12:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:13:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:14:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:15:5
	output wire grant_valid;
	// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:18:5
	generate
		if (NUM_REQS == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:23:9
			assign grant_index = 0;
			// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:24:9
			assign grant_onehot = requests;
			// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:25:9
			assign grant_valid = requests[0];
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:29:9
			reg [NUM_REQS - 1:1] state [NUM_REQS - 1:0];
			// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:30:9
			wire [NUM_REQS - 1:0] pri [NUM_REQS - 1:0];
			// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:31:9
			wire [NUM_REQS - 1:0] grant_unqual;
			genvar i;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
				genvar j;
				for (j = 0; j < NUM_REQS; j = j + 1) begin : genblk1
					if (j > i) begin : genblk1
						// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:36:21
						assign pri[j][i] = requests[i] && state[i][j];
					end
					else if (j < i) begin : genblk1
						// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:39:21
						assign pri[j][i] = requests[i] && !state[j][i];
					end
					else begin : genblk1
						// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:42:21
						assign pri[j][i] = 0;
					end
				end
				// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:45:13
				assign grant_unqual[i] = requests[i] && !(|pri[i]);
			end
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk2
				genvar j;
				for (j = i + 1; j < NUM_REQS; j = j + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:50:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:51:21
						if (reset)
							// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:52:25
							state[i][j] <= 0;
						else
							// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:54:25
							state[i][j] <= (state[i][j] || grant_unqual[j]) && !grant_unqual[i];
				end
			end
			if (LOCK_ENABLE == 0) begin : genblk3
				// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:62:13
				assign grant_onehot = grant_unqual;
			end
			else begin : genblk3
				// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:64:13
				reg [NUM_REQS - 1:0] grant_unqual_prev;
				// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:65:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:66:17
					if (reset)
						// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:67:21
						grant_unqual_prev <= 0;
					else if (enable)
						// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:69:21
						grant_unqual_prev <= grant_unqual;
				// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:72:13
				assign grant_onehot = (enable ? grant_unqual : grant_unqual_prev);
			end
			// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:75:9
			VX_onehot_encoder #(.N(NUM_REQS)) encoder(
				.data_in(grant_unqual),
				.data_out(grant_index)
			);
			// Trace: ../../rtl/libs/VX_matrix_arbiter.sv:83:9
			assign grant_valid = |requests;
		end
	endgenerate
endmodule
module VX_multiplier (
	clk,
	enable,
	dataa,
	datab,
	result
);
	// Trace: ../../rtl/libs/VX_multiplier.sv:5:15
	parameter WIDTHA = 1;
	// Trace: ../../rtl/libs/VX_multiplier.sv:6:15
	parameter WIDTHB = 1;
	// Trace: ../../rtl/libs/VX_multiplier.sv:7:15
	parameter WIDTHP = 1;
	// Trace: ../../rtl/libs/VX_multiplier.sv:8:15
	parameter SIGNED = 0;
	// Trace: ../../rtl/libs/VX_multiplier.sv:9:15
	parameter LATENCY = 0;
	// Trace: ../../rtl/libs/VX_multiplier.sv:11:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_multiplier.sv:12:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_multiplier.sv:13:5
	input wire [WIDTHA - 1:0] dataa;
	// Trace: ../../rtl/libs/VX_multiplier.sv:14:5
	input wire [WIDTHB - 1:0] datab;
	// Trace: ../../rtl/libs/VX_multiplier.sv:15:5
	output wire [WIDTHP - 1:0] result;
	// Trace: ../../rtl/libs/VX_multiplier.sv:40:5
	wire [WIDTHP - 1:0] result_unqual;
	// Trace: ../../rtl/libs/VX_multiplier.sv:42:5
	generate
		if (SIGNED) begin : genblk1
			// Trace: ../../rtl/libs/VX_multiplier.sv:43:9
			assign result_unqual = $signed(dataa) * $signed(datab);
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_multiplier.sv:45:9
			assign result_unqual = dataa * datab;
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_multiplier.sv:48:5
	generate
		if (LATENCY == 0) begin : genblk2
			// Trace: ../../rtl/libs/VX_multiplier.sv:49:9
			assign result = result_unqual;
		end
		else begin : genblk2
			// Trace: ../../rtl/libs/VX_multiplier.sv:51:9
			reg [WIDTHP - 1:0] result_pipe [LATENCY - 1:0];
			// Trace: ../../rtl/libs/VX_multiplier.sv:52:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_multiplier.sv:53:13
				if (enable)
					// Trace: ../../rtl/libs/VX_multiplier.sv:54:17
					result_pipe[0] <= result_unqual;
			genvar i;
			for (i = 1; i < LATENCY; i = i + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_multiplier.sv:58:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_multiplier.sv:59:17
					if (enable)
						// Trace: ../../rtl/libs/VX_multiplier.sv:60:21
						result_pipe[i] <= result_pipe[i - 1];
			end
			// Trace: ../../rtl/libs/VX_multiplier.sv:64:9
			assign result = result_pipe[LATENCY - 1];
		end
	endgenerate
endmodule
module VX_mux (
	data_in,
	sel_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_mux.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_mux.sv:6:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_mux.sv:7:15
	parameter LN = $clog2(N);
	// Trace: ../../rtl/libs/VX_mux.sv:9:5
	input wire [(N * DATAW) - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_mux.sv:10:5
	input wire [LN - 1:0] sel_in;
	// Trace: ../../rtl/libs/VX_mux.sv:11:5
	output wire [DATAW - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_mux.sv:13:5
	generate
		if (N > 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_mux.sv:14:9
			assign data_out = data_in[sel_in * DATAW+:DATAW];
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_mux.sv:17:9
			assign data_out = data_in;
		end
	endgenerate
endmodule
module VX_onehot_encoder (
	data_in,
	data_out,
	valid_out
);
	// Trace: ../../rtl/libs/VX_onehot_encoder.sv:8:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_onehot_encoder.sv:9:15
	parameter REVERSE = 0;
	// Trace: ../../rtl/libs/VX_onehot_encoder.sv:10:15
	parameter MODEL = 1;
	// Trace: ../../rtl/libs/VX_onehot_encoder.sv:11:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: ../../rtl/libs/VX_onehot_encoder.sv:13:5
	input wire [N - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_onehot_encoder.sv:14:5
	output wire [LN - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_onehot_encoder.sv:15:5
	output wire valid_out;
	// Trace: ../../rtl/libs/VX_onehot_encoder.sv:17:5
	function automatic signed [(N > 1 ? $clog2(N) : 1) - 1:0] sv2v_cast_374F3_signed;
		input reg signed [(N > 1 ? $clog2(N) : 1) - 1:0] inp;
		sv2v_cast_374F3_signed = inp;
	endfunction
	generate
		if (N == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:19:9
			assign data_out = data_in;
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:20:9
			assign valid_out = data_in;
		end
		else if (N == 2) begin : genblk1
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:24:9
			assign data_out = data_in[!REVERSE];
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:25:9
			assign valid_out = |data_in;
		end
		else if (MODEL == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:29:9
			localparam levels_lp = $clog2(N);
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:30:9
			localparam aligned_width_lp = 1 << $clog2(N);
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:32:9
			wire [(levels_lp >= 0 ? ((levels_lp + 1) * aligned_width_lp) - 1 : ((1 - levels_lp) * aligned_width_lp) + ((levels_lp * aligned_width_lp) - 1)):(levels_lp >= 0 ? 0 : levels_lp * aligned_width_lp)] addr;
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:33:9
			wire [(levels_lp >= 0 ? ((levels_lp + 1) * aligned_width_lp) - 1 : ((1 - levels_lp) * aligned_width_lp) + ((levels_lp * aligned_width_lp) - 1)):(levels_lp >= 0 ? 0 : levels_lp * aligned_width_lp)] v;
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:36:9
			function automatic [aligned_width_lp - 1:0] sv2v_cast_65C44;
				input reg [aligned_width_lp - 1:0] inp;
				sv2v_cast_65C44 = inp;
			endfunction
			assign v[(levels_lp >= 0 ? 0 : levels_lp) * aligned_width_lp+:aligned_width_lp] = (REVERSE ? data_in << (aligned_width_lp - N) : sv2v_cast_65C44(data_in));
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:37:9
			assign addr[(levels_lp >= 0 ? 0 : levels_lp) * aligned_width_lp+:aligned_width_lp] = 1'sbx;
			genvar level;
			for (level = 1; level < (levels_lp + 1); level = level + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_onehot_encoder.sv:40:13
				localparam segments_lp = 2 ** (levels_lp - level);
				// Trace: ../../rtl/libs/VX_onehot_encoder.sv:41:13
				localparam segment_slot_lp = aligned_width_lp / segments_lp;
				// Trace: ../../rtl/libs/VX_onehot_encoder.sv:42:13
				localparam segment_width_lp = level;
				genvar segment;
				for (segment = 0; segment < segments_lp; segment = segment + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_onehot_encoder.sv:45:17
					wire [1:0] vs = {v[((levels_lp >= 0 ? level - 1 : levels_lp - (level - 1)) * aligned_width_lp) + ((segment * segment_slot_lp) + (segment_slot_lp >> 1))], v[((levels_lp >= 0 ? level - 1 : levels_lp - (level - 1)) * aligned_width_lp) + (segment * segment_slot_lp)]};
					// Trace: ../../rtl/libs/VX_onehot_encoder.sv:50:17
					assign v[((levels_lp >= 0 ? level : levels_lp - level) * aligned_width_lp) + (segment * segment_slot_lp)] = |vs;
					if (level == 1) begin : genblk1
						// Trace: ../../rtl/libs/VX_onehot_encoder.sv:53:21
						assign addr[((levels_lp >= 0 ? level : levels_lp - level) * aligned_width_lp) + (segment * segment_slot_lp)+:segment_width_lp] = vs[!REVERSE];
					end
					else begin : genblk1
						// Trace: ../../rtl/libs/VX_onehot_encoder.sv:55:21
						assign addr[((levels_lp >= 0 ? level : levels_lp - level) * aligned_width_lp) + (segment * segment_slot_lp)+:segment_width_lp] = {vs[!REVERSE], addr[((levels_lp >= 0 ? level - 1 : levels_lp - (level - 1)) * aligned_width_lp) + (segment * segment_slot_lp)+:segment_width_lp - 1] | addr[((levels_lp >= 0 ? level - 1 : levels_lp - (level - 1)) * aligned_width_lp) + ((segment * segment_slot_lp) + (segment_slot_lp >> 1))+:segment_width_lp - 1]};
					end
				end
			end
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:63:9
			assign data_out = addr[((levels_lp >= 0 ? levels_lp : levels_lp - levels_lp) * aligned_width_lp) + ((N > 1 ? $clog2(N) : 1) - 1)-:(N > 1 ? $clog2(N) : 1)];
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:64:9
			assign valid_out = v[(levels_lp >= 0 ? levels_lp : levels_lp - levels_lp) * aligned_width_lp];
		end
		else if (MODEL == 2) begin : genblk1
			genvar j;
			for (j = 0; j < LN; j = j + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_onehot_encoder.sv:69:13
				wire [N - 1:0] mask;
				genvar i;
				for (i = 0; i < N; i = i + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_onehot_encoder.sv:71:17
					assign mask[i] = i[j];
				end
				// Trace: ../../rtl/libs/VX_onehot_encoder.sv:73:13
				assign data_out[j] = |(mask & data_in);
			end
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:76:9
			assign valid_out = |data_in;
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:80:9
			reg [LN - 1:0] index_r;
			if (REVERSE) begin : genblk1
				// Trace: ../../rtl/libs/VX_onehot_encoder.sv:83:13
				always @(*) begin
					// Trace: ../../rtl/libs/VX_onehot_encoder.sv:84:17
					index_r = 1'sbx;
					// Trace: ../../rtl/libs/VX_onehot_encoder.sv:85:17
					begin : sv2v_autoblock_1
						// Trace: ../../rtl/libs/VX_onehot_encoder.sv:85:22
						integer i;
						// Trace: ../../rtl/libs/VX_onehot_encoder.sv:85:22
						for (i = N - 1; i >= 0; i = i - 1)
							begin
								// Trace: ../../rtl/libs/VX_onehot_encoder.sv:86:21
								if (data_in[i])
									// Trace: ../../rtl/libs/VX_onehot_encoder.sv:87:25
									index_r = sv2v_cast_374F3_signed(i);
							end
					end
				end
			end
			else begin : genblk1
				// Trace: ../../rtl/libs/VX_onehot_encoder.sv:92:13
				always @(*) begin
					// Trace: ../../rtl/libs/VX_onehot_encoder.sv:93:17
					index_r = 1'sbx;
					// Trace: ../../rtl/libs/VX_onehot_encoder.sv:94:17
					begin : sv2v_autoblock_2
						// Trace: ../../rtl/libs/VX_onehot_encoder.sv:94:22
						integer i;
						// Trace: ../../rtl/libs/VX_onehot_encoder.sv:94:22
						for (i = 0; i < N; i = i + 1)
							begin
								// Trace: ../../rtl/libs/VX_onehot_encoder.sv:95:21
								if (data_in[i])
									// Trace: ../../rtl/libs/VX_onehot_encoder.sv:96:25
									index_r = sv2v_cast_374F3_signed(i);
							end
					end
				end
			end
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:102:9
			assign data_out = index_r;
			// Trace: ../../rtl/libs/VX_onehot_encoder.sv:103:9
			assign valid_out = |data_in;
		end
	endgenerate
endmodule
module VX_onehot_mux (
	data_in,
	sel_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_onehot_mux.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_onehot_mux.sv:6:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_onehot_mux.sv:7:15
	parameter MODEL = 1;
	// Trace: ../../rtl/libs/VX_onehot_mux.sv:9:5
	input wire [(N * DATAW) - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_onehot_mux.sv:10:5
	input wire [N - 1:0] sel_in;
	// Trace: ../../rtl/libs/VX_onehot_mux.sv:11:5
	output wire [DATAW - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_onehot_mux.sv:13:5
	generate
		if (N > 1) begin : genblk1
			if (MODEL == 1) begin : genblk1
				genvar i;
				for (i = 0; i < N; i = i + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_onehot_mux.sv:16:17
					assign data_out = (sel_in[i] ? data_in[i * DATAW+:DATAW] : {DATAW {1'sbz}});
				end
			end
			else if (MODEL == 2) begin : genblk1
				// Trace: ../../rtl/libs/VX_onehot_mux.sv:19:13
				reg [DATAW - 1:0] data_out_r;
				// Trace: ../../rtl/libs/VX_onehot_mux.sv:20:13
				always @(*) begin
					// Trace: ../../rtl/libs/VX_onehot_mux.sv:21:17
					data_out_r = 1'sb0;
					// Trace: ../../rtl/libs/VX_onehot_mux.sv:22:17
					begin : sv2v_autoblock_1
						// Trace: ../../rtl/libs/VX_onehot_mux.sv:22:22
						integer i;
						// Trace: ../../rtl/libs/VX_onehot_mux.sv:22:22
						for (i = 0; i < N; i = i + 1)
							begin
								// Trace: ../../rtl/libs/VX_onehot_mux.sv:23:21
								data_out_r = data_out_r | ({DATAW {sel_in[i]}} & data_in[i * DATAW+:DATAW]);
							end
					end
				end
				// Trace: ../../rtl/libs/VX_onehot_mux.sv:26:13
				assign data_out = data_out_r;
			end
			else if (MODEL == 3) begin : genblk1
				// Trace: ../../rtl/libs/VX_onehot_mux.sv:28:13
				wire [(N * DATAW) - 1:0] mask;
				genvar i;
				for (i = 0; i < N; i = i + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_onehot_mux.sv:30:17
					assign mask[i * DATAW+:DATAW] = {DATAW {sel_in[i]}} & data_in[i * DATAW+:DATAW];
				end
				for (i = 0; i < DATAW; i = i + 1) begin : genblk2
					// Trace: ../../rtl/libs/VX_onehot_mux.sv:33:17
					wire [N - 1:0] gather;
					genvar j;
					for (j = 0; j < N; j = j + 1) begin : genblk1
						// Trace: ../../rtl/libs/VX_onehot_mux.sv:35:21
						assign gather[j] = mask[(j * DATAW) + i];
					end
					// Trace: ../../rtl/libs/VX_onehot_mux.sv:37:17
					assign data_out[i] = |gather;
				end
			end
			else begin : genblk1
				// Trace: ../../rtl/libs/VX_onehot_mux.sv:40:13
				reg [DATAW - 1:0] data_out_r;
				// Trace: ../../rtl/libs/VX_onehot_mux.sv:41:13
				always @(*) begin
					// Trace: ../../rtl/libs/VX_onehot_mux.sv:42:17
					data_out_r = 1'sbx;
					// Trace: ../../rtl/libs/VX_onehot_mux.sv:43:17
					begin : sv2v_autoblock_2
						// Trace: ../../rtl/libs/VX_onehot_mux.sv:43:22
						integer i;
						// Trace: ../../rtl/libs/VX_onehot_mux.sv:43:22
						for (i = N - 1; i >= 0; i = i - 1)
							begin
								// Trace: ../../rtl/libs/VX_onehot_mux.sv:44:21
								if (sel_in[i])
									// Trace: ../../rtl/libs/VX_onehot_mux.sv:45:25
									data_out_r = data_in[i * DATAW+:DATAW];
							end
					end
				end
				// Trace: ../../rtl/libs/VX_onehot_mux.sv:49:13
				assign data_out = data_out_r;
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_onehot_mux.sv:53:9
			assign data_out = data_in;
		end
	endgenerate
endmodule
module VX_pending_size (
	clk,
	reset,
	incr,
	decr,
	empty,
	full,
	size
);
	// Trace: ../../rtl/libs/VX_pending_size.sv:5:15
	parameter SIZE = 1;
	// Trace: ../../rtl/libs/VX_pending_size.sv:6:15
	parameter SIZEW = $clog2(SIZE + 1);
	// Trace: ../../rtl/libs/VX_pending_size.sv:8:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_pending_size.sv:9:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_pending_size.sv:10:5
	input wire incr;
	// Trace: ../../rtl/libs/VX_pending_size.sv:11:5
	input wire decr;
	// Trace: ../../rtl/libs/VX_pending_size.sv:12:5
	output wire empty;
	// Trace: ../../rtl/libs/VX_pending_size.sv:13:5
	output wire full;
	// Trace: ../../rtl/libs/VX_pending_size.sv:14:5
	output wire [SIZEW - 1:0] size;
	// Trace: ../../rtl/libs/VX_pending_size.sv:16:5
	localparam ADDRW = $clog2(SIZE);
	// Trace: ../../rtl/libs/VX_pending_size.sv:18:5
	reg [ADDRW - 1:0] used_r;
	// Trace: ../../rtl/libs/VX_pending_size.sv:19:5
	reg empty_r;
	// Trace: ../../rtl/libs/VX_pending_size.sv:20:5
	reg full_r;
	// Trace: ../../rtl/libs/VX_pending_size.sv:22:5
	function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
		input reg signed [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D_signed = inp;
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	always @(posedge clk)
		// Trace: ../../rtl/libs/VX_pending_size.sv:23:9
		if (reset) begin
			// Trace: ../../rtl/libs/VX_pending_size.sv:24:13
			used_r <= 0;
			// Trace: ../../rtl/libs/VX_pending_size.sv:25:13
			empty_r <= 1;
			// Trace: ../../rtl/libs/VX_pending_size.sv:26:13
			full_r <= 0;
		end
		else begin
			// Trace: macro expansion of ASSERT at ../../rtl/libs/VX_pending_size.sv:28:48
			if (!incr || !full)
				;
			if (incr) begin
				begin
					// Trace: ../../rtl/libs/VX_pending_size.sv:30:17
					if (!decr) begin
						// Trace: ../../rtl/libs/VX_pending_size.sv:31:21
						empty_r <= 0;
						// Trace: ../../rtl/libs/VX_pending_size.sv:32:21
						if (used_r == sv2v_cast_8BB5D_signed(SIZE - 1))
							// Trace: ../../rtl/libs/VX_pending_size.sv:33:25
							full_r <= 1;
					end
				end
			end
			else if (decr) begin
				// Trace: ../../rtl/libs/VX_pending_size.sv:36:17
				full_r <= 0;
				// Trace: ../../rtl/libs/VX_pending_size.sv:37:17
				if (used_r == sv2v_cast_8BB5D_signed(1))
					// Trace: ../../rtl/libs/VX_pending_size.sv:38:21
					empty_r <= 1;
			end
			// Trace: ../../rtl/libs/VX_pending_size.sv:40:13
			used_r <= used_r + sv2v_cast_8BB5D_signed($signed(sv2v_cast_2(incr && !decr) - sv2v_cast_2(decr && !incr)));
		end
	// Trace: ../../rtl/libs/VX_pending_size.sv:44:5
	assign empty = empty_r;
	// Trace: ../../rtl/libs/VX_pending_size.sv:45:5
	assign full = full_r;
	// Trace: ../../rtl/libs/VX_pending_size.sv:46:5
	assign size = {full_r, used_r};
endmodule
module VX_pipe_register (
	clk,
	reset,
	enable,
	data_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_pipe_register.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_pipe_register.sv:6:15
	parameter RESETW = DATAW;
	// Trace: ../../rtl/libs/VX_pipe_register.sv:7:15
	parameter DEPTH = 1;
	// Trace: ../../rtl/libs/VX_pipe_register.sv:9:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_pipe_register.sv:10:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_pipe_register.sv:11:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_pipe_register.sv:12:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_pipe_register.sv:13:5
	output wire [DATAW - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_pipe_register.sv:16:5
	function automatic signed [RESETW - 1:0] sv2v_cast_5A382_signed;
		input reg signed [RESETW - 1:0] inp;
		sv2v_cast_5A382_signed = inp;
	endfunction
	generate
		if (DEPTH == 0) begin : genblk1
			// Trace: ../../rtl/libs/VX_pipe_register.sv:20:9
			assign data_out = data_in;
		end
		else if (DEPTH == 1) begin : genblk1
			if (RESETW == 0) begin : genblk1
				// Trace: ../../rtl/libs/VX_pipe_register.sv:24:13
				reg [DATAW - 1:0] value;
				// Trace: ../../rtl/libs/VX_pipe_register.sv:26:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_pipe_register.sv:27:17
					if (enable)
						// Trace: ../../rtl/libs/VX_pipe_register.sv:28:21
						value <= data_in;
				// Trace: ../../rtl/libs/VX_pipe_register.sv:31:13
				assign data_out = value;
			end
			else if (RESETW == DATAW) begin : genblk1
				// Trace: ../../rtl/libs/VX_pipe_register.sv:33:13
				reg [DATAW - 1:0] value;
				// Trace: ../../rtl/libs/VX_pipe_register.sv:35:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_pipe_register.sv:36:17
					if (reset)
						// Trace: ../../rtl/libs/VX_pipe_register.sv:37:21
						value <= sv2v_cast_5A382_signed(0);
					else if (enable)
						// Trace: ../../rtl/libs/VX_pipe_register.sv:39:21
						value <= data_in;
				// Trace: ../../rtl/libs/VX_pipe_register.sv:42:13
				assign data_out = value;
			end
			else begin : genblk1
				// Trace: ../../rtl/libs/VX_pipe_register.sv:44:13
				reg [(DATAW - RESETW) - 1:0] value_d;
				// Trace: ../../rtl/libs/VX_pipe_register.sv:45:13
				reg [RESETW - 1:0] value_r;
				// Trace: ../../rtl/libs/VX_pipe_register.sv:47:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_pipe_register.sv:48:17
					if (reset)
						// Trace: ../../rtl/libs/VX_pipe_register.sv:49:21
						value_r <= sv2v_cast_5A382_signed(0);
					else if (enable)
						// Trace: ../../rtl/libs/VX_pipe_register.sv:51:21
						value_r <= data_in[DATAW - 1:DATAW - RESETW];
				// Trace: ../../rtl/libs/VX_pipe_register.sv:55:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_pipe_register.sv:56:17
					if (enable)
						// Trace: ../../rtl/libs/VX_pipe_register.sv:57:21
						value_d <= data_in[(DATAW - RESETW) - 1:0];
				// Trace: ../../rtl/libs/VX_pipe_register.sv:60:13
				assign data_out = {value_r, value_d};
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_pipe_register.sv:63:9
			VX_shift_register #(
				.DATAW(DATAW),
				.RESETW(RESETW),
				.DEPTH(DEPTH)
			) shift_reg(
				.clk(clk),
				.reset(reset),
				.enable(enable),
				.data_in(data_in),
				.data_out(data_out)
			);
		end
	endgenerate
endmodule
module VX_popcount (
	in_i,
	cnt_o
);
	// Trace: ../../rtl/libs/VX_popcount.sv:5:15
	parameter MODEL = 1;
	// Trace: ../../rtl/libs/VX_popcount.sv:6:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_popcount.sv:7:15
	parameter M = $clog2(N + 1);
	// Trace: ../../rtl/libs/VX_popcount.sv:9:5
	input wire [N - 1:0] in_i;
	// Trace: ../../rtl/libs/VX_popcount.sv:10:5
	output wire [M - 1:0] cnt_o;
	// Trace: ../../rtl/libs/VX_popcount.sv:20:5
	generate
		if (N == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_popcount.sv:22:9
			assign cnt_o = in_i;
		end
		else if (MODEL == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_popcount.sv:26:9
			localparam PN = 1 << $clog2(N);
			// Trace: ../../rtl/libs/VX_popcount.sv:27:9
			localparam LOGPN = $clog2(PN);
			// Trace: ../../rtl/libs/VX_popcount.sv:29:9
			wire [M - 1:0] tmp [0:PN - 1][0:PN - 1];
			genvar i;
			for (i = 0; i < N; i = i + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_popcount.sv:32:13
				assign tmp[0][i] = in_i[i];
			end
			for (i = N; i < PN; i = i + 1) begin : genblk2
				// Trace: ../../rtl/libs/VX_popcount.sv:36:13
				assign tmp[0][i] = 1'sb0;
			end
			genvar j;
			for (j = 0; j < LOGPN; j = j + 1) begin : genblk3
				genvar i;
				for (i = 0; i < (1 << ((LOGPN - j) - 1)); i = i + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_popcount.sv:41:17
					assign tmp[j + 1][i] = tmp[j][i * 2] + tmp[j][(i * 2) + 1];
				end
			end
			// Trace: ../../rtl/libs/VX_popcount.sv:45:9
			assign cnt_o = tmp[LOGPN][0];
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_popcount.sv:49:9
			reg [M - 1:0] cnt_r;
			// Trace: ../../rtl/libs/VX_popcount.sv:51:9
			always @(*) begin
				// Trace: ../../rtl/libs/VX_popcount.sv:52:13
				cnt_r = 1'sb0;
				// Trace: ../../rtl/libs/VX_popcount.sv:53:13
				begin : sv2v_autoblock_1
					// Trace: ../../rtl/libs/VX_popcount.sv:53:18
					integer i;
					// Trace: ../../rtl/libs/VX_popcount.sv:53:18
					for (i = 0; i < N; i = i + 1)
						begin
							// Trace: ../../rtl/libs/VX_popcount.sv:55:17
							cnt_r = cnt_r + in_i[i];
						end
				end
			end
			// Trace: ../../rtl/libs/VX_popcount.sv:60:9
			assign cnt_o = cnt_r;
		end
	endgenerate
endmodule
module VX_priority_encoder (
	data_in,
	onehot,
	index,
	valid_out
);
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:5:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:6:15
	parameter REVERSE = 0;
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:7:15
	parameter MODEL = 1;
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:8:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:10:5
	input wire [N - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:11:5
	output wire [N - 1:0] onehot;
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:12:5
	output wire [LN - 1:0] index;
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:13:5
	output wire valid_out;
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:15:5
	wire [N - 1:0] reversed;
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:17:5
	generate
		if (REVERSE) begin : genblk1
			genvar i;
			for (i = 0; i < N; i = i + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_priority_encoder.sv:19:13
				assign reversed[(N - i) - 1] = data_in[i];
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:22:9
			assign reversed = data_in;
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_priority_encoder.sv:25:5
	function automatic signed [LN - 1:0] sv2v_cast_83428_signed;
		input reg signed [LN - 1:0] inp;
		sv2v_cast_83428_signed = inp;
	endfunction
	generate
		if (N == 1) begin : genblk2
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:27:9
			assign onehot = reversed;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:28:9
			assign index = 0;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:29:9
			assign valid_out = reversed;
		end
		else if (N == 2) begin : genblk2
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:33:9
			assign onehot = {~reversed[0], reversed[0]};
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:34:9
			assign index = ~reversed[0];
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:35:9
			assign valid_out = |reversed;
		end
		else if (MODEL == 1) begin : genblk2
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:39:9
			wire [N - 1:0] scan_lo;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:41:9
			VX_scan #(
				.N(N),
				.OP(2)
			) scan(
				.data_in(reversed),
				.data_out(scan_lo)
			);
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:49:9
			VX_lzc #(.N(N)) lzc(
				.in_i(reversed),
				.cnt_o(index)
			);
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:57:9
			assign onehot = scan_lo & {~scan_lo[N - 2:0], 1'b1};
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:58:9
			assign valid_out = scan_lo[N - 1];
		end
		else if (MODEL == 2) begin : genblk2
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:63:9
			wire [N - 1:0] higher_pri_regs;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:65:9
			assign higher_pri_regs[N - 1:1] = higher_pri_regs[N - 2:0] | reversed[N - 2:0];
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:66:9
			assign higher_pri_regs[0] = 1'b0;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:67:9
			assign onehot[N - 1:0] = reversed[N - 1:0] & ~higher_pri_regs[N - 1:0];
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:69:9
			VX_lzc #(.N(N)) lzc(
				.in_i(reversed),
				.cnt_o(index),
				.valid_o(valid_out)
			);
		end
		else if (MODEL == 3) begin : genblk2
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:79:9
			assign onehot = reversed & ~(reversed - 1);
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:81:9
			VX_lzc #(.N(N)) lzc(
				.in_i(reversed),
				.cnt_o(index),
				.valid_o(valid_out)
			);
		end
		else begin : genblk2
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:91:9
			reg [LN - 1:0] index_r;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:92:9
			reg [N - 1:0] onehot_r;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:94:9
			always @(*) begin
				// Trace: ../../rtl/libs/VX_priority_encoder.sv:95:13
				index_r = 1'sbx;
				// Trace: ../../rtl/libs/VX_priority_encoder.sv:96:13
				onehot_r = 1'sbx;
				// Trace: ../../rtl/libs/VX_priority_encoder.sv:97:13
				begin : sv2v_autoblock_1
					// Trace: ../../rtl/libs/VX_priority_encoder.sv:97:18
					integer i;
					// Trace: ../../rtl/libs/VX_priority_encoder.sv:97:18
					for (i = N - 1; i >= 0; i = i - 1)
						begin
							// Trace: ../../rtl/libs/VX_priority_encoder.sv:98:17
							if (reversed[i]) begin
								// Trace: ../../rtl/libs/VX_priority_encoder.sv:99:21
								index_r = sv2v_cast_83428_signed(i);
								// Trace: ../../rtl/libs/VX_priority_encoder.sv:100:21
								onehot_r = 0;
								// Trace: ../../rtl/libs/VX_priority_encoder.sv:101:21
								onehot_r[i] = 1'b1;
							end
						end
				end
			end
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:106:9
			assign index = index_r;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:107:9
			assign onehot = onehot_r;
			// Trace: ../../rtl/libs/VX_priority_encoder.sv:108:9
			assign valid_out = |reversed;
		end
	endgenerate
endmodule
module VX_reset_relay (
	clk,
	reset,
	reset_o
);
	// Trace: ../../rtl/libs/VX_reset_relay.sv:4:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_reset_relay.sv:5:15
	parameter DEPTH = 1;
	// Trace: ../../rtl/libs/VX_reset_relay.sv:7:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_reset_relay.sv:8:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_reset_relay.sv:9:5
	output wire [N - 1:0] reset_o;
	// Trace: ../../rtl/libs/VX_reset_relay.sv:12:5
	generate
		if (DEPTH > 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_reset_relay.sv:13:37
			reg [N - 1:0] reset_r [DEPTH - 1:0];
			// Trace: ../../rtl/libs/VX_reset_relay.sv:14:9
			always @(posedge clk) begin
				// Trace: ../../rtl/libs/VX_reset_relay.sv:15:13
				begin : sv2v_autoblock_1
					// Trace: ../../rtl/libs/VX_reset_relay.sv:15:18
					integer i;
					// Trace: ../../rtl/libs/VX_reset_relay.sv:15:18
					for (i = DEPTH - 1; i > 0; i = i - 1)
						begin
							// Trace: ../../rtl/libs/VX_reset_relay.sv:16:17
							reset_r[i] <= reset_r[i - 1];
						end
				end
				// Trace: ../../rtl/libs/VX_reset_relay.sv:17:13
				reset_r[0] <= {N {reset}};
			end
			// Trace: ../../rtl/libs/VX_reset_relay.sv:19:9
			assign reset_o = reset_r[DEPTH - 1];
		end
		else if (DEPTH == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_reset_relay.sv:21:23
			reg [N - 1:0] reset_r;
			// Trace: ../../rtl/libs/VX_reset_relay.sv:22:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_reset_relay.sv:23:13
				reset_r <= {N {reset}};
			// Trace: ../../rtl/libs/VX_reset_relay.sv:25:9
			assign reset_o = reset_r;
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_reset_relay.sv:28:9
			assign reset_o = {N {reset}};
		end
	endgenerate
endmodule
module VX_rr_arbiter (
	clk,
	reset,
	enable,
	requests,
	grant_index,
	grant_onehot,
	grant_valid
);
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:5:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:6:15
	parameter LOCK_ENABLE = 0;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:7:15
	parameter MODEL = 1;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:8:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:10:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:11:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:12:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:13:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:14:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:15:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:16:5
	output wire grant_valid;
	// Trace: ../../rtl/libs/VX_rr_arbiter.sv:19:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_REQS == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:24:9
			assign grant_index = 0;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:25:9
			assign grant_onehot = requests;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:26:9
			assign grant_valid = requests[0];
		end
		else if (NUM_REQS == 2) begin : genblk1
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:30:9
			reg [LOG_NUM_REQS - 1:0] grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:31:9
			reg [NUM_REQS - 1:0] grant_onehot_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:32:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:34:9
			always @(*)
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:35:13
				casez ({state, requests})
					3'b001, 3'b1z1: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:37:28
						grant_onehot_r = 2'b01;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:37:52
						grant_index_r = sv2v_cast_76B5F_signed(0);
					end
					default: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:38:28
						grant_onehot_r = 2'b10;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:38:52
						grant_index_r = sv2v_cast_76B5F_signed(1);
					end
				endcase
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:42:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:43:13
				if (reset)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:44:17
					state <= 0;
				else if (!LOCK_ENABLE || enable)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:46:17
					state <= grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:50:9
			assign grant_index = grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:51:9
			assign grant_onehot = grant_onehot_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:52:9
			assign grant_valid = |requests;
		end
		else if (NUM_REQS == 4) begin : genblk1
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:56:9
			reg [LOG_NUM_REQS - 1:0] grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:57:9
			reg [NUM_REQS - 1:0] grant_onehot_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:58:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:60:9
			always @(*)
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:61:13
				casez ({state, requests})
					6'b000001, 6'b0100z1, 6'b100zz1, 6'b11zzz1: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:65:31
						grant_onehot_r = 4'b0001;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:65:57
						grant_index_r = sv2v_cast_76B5F_signed(0);
					end
					6'b00zz1z, 6'b010010, 6'b100z10, 6'b11zz10: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:69:31
						grant_onehot_r = 4'b0010;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:69:57
						grant_index_r = sv2v_cast_76B5F_signed(1);
					end
					6'b00z10z, 6'b01z1zz, 6'b100100, 6'b11z100: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:73:31
						grant_onehot_r = 4'b0100;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:73:57
						grant_index_r = sv2v_cast_76B5F_signed(2);
					end
					default: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:74:31
						grant_onehot_r = 4'b1000;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:74:57
						grant_index_r = sv2v_cast_76B5F_signed(3);
					end
				endcase
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:78:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:79:13
				if (reset)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:80:17
					state <= 0;
				else if (!LOCK_ENABLE || enable)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:82:17
					state <= grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:86:9
			assign grant_index = grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:87:9
			assign grant_onehot = grant_onehot_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:88:9
			assign grant_valid = |requests;
		end
		else if (NUM_REQS == 8) begin : genblk1
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:92:9
			reg [LOG_NUM_REQS - 1:0] grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:93:9
			reg [NUM_REQS - 1:0] grant_onehot_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:94:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:96:9
			always @(*)
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:97:13
				casez ({state, requests})
					11'b00000000001, 11'b001000000z1, 11'b01000000zz1, 11'b0110000zzz1, 11'b100000zzzz1, 11'b10100zzzzz1, 11'b1100zzzzzz1, 11'b111zzzzzzz1: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:105:37
						grant_onehot_r = 8'b00000001;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:105:67
						grant_index_r = sv2v_cast_76B5F_signed(0);
					end
					11'b000zzzzzz1z, 11'b00100000010, 11'b01000000z10, 11'b0110000zz10, 11'b100000zzz10, 11'b10100zzzz10, 11'b1100zzzzz10, 11'b111zzzzzz10: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:113:37
						grant_onehot_r = 8'b00000010;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:113:67
						grant_index_r = sv2v_cast_76B5F_signed(1);
					end
					11'b000zzzzz10z, 11'b001zzzzz1zz, 11'b01000000100, 11'b0110000z100, 11'b100000zz100, 11'b10100zzz100, 11'b1100zzzz100, 11'b111zzzzz100: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:121:37
						grant_onehot_r = 8'b00000100;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:121:67
						grant_index_r = sv2v_cast_76B5F_signed(2);
					end
					11'b000zzzz100z, 11'b001zzzz10zz, 11'b010zzzz1zzz, 11'b01100001000, 11'b100000z1000, 11'b10100zz1000, 11'b1100zzz1000, 11'b111zzzz1000: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:129:37
						grant_onehot_r = 8'b00001000;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:129:67
						grant_index_r = sv2v_cast_76B5F_signed(3);
					end
					11'b000zzz1000z, 11'b001zzz100zz, 11'b010zzz10zzz, 11'b011zzz1zzzz, 11'b10000010000, 11'b10100z10000, 11'b1100zz10000, 11'b111zzz10000: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:137:37
						grant_onehot_r = 8'b00010000;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:137:67
						grant_index_r = sv2v_cast_76B5F_signed(4);
					end
					11'b000zz10000z, 11'b001zz1000zz, 11'b010zz100zzz, 11'b011zz10zzzz, 11'b100zz1zzzzz, 11'b10100100000, 11'b1100z100000, 11'b111zz100000: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:145:37
						grant_onehot_r = 8'b00100000;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:145:67
						grant_index_r = sv2v_cast_76B5F_signed(5);
					end
					11'b000z100000z, 11'b001z10000zz, 11'b010z1000zzz, 11'b011z100zzzz, 11'b100z10zzzzz, 11'b101z1zzzzzz, 11'b11001000000, 11'b111z1000000: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:153:37
						grant_onehot_r = 8'b01000000;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:153:67
						grant_index_r = sv2v_cast_76B5F_signed(6);
					end
					default: begin
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:154:37
						grant_onehot_r = 8'b10000000;
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:154:67
						grant_index_r = sv2v_cast_76B5F_signed(7);
					end
				endcase
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:158:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:159:13
				if (reset)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:160:17
					state <= 0;
				else if (!LOCK_ENABLE || enable)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:162:17
					state <= grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:166:9
			assign grant_index = grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:167:9
			assign grant_onehot = grant_onehot_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:168:9
			assign grant_valid = |requests;
		end
		else if (MODEL == 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:173:9
			wire [NUM_REQS - 1:0] mask_higher_pri_regs;
			wire [NUM_REQS - 1:0] unmask_higher_pri_regs;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:175:9
			wire [NUM_REQS - 1:0] grant_masked;
			wire [NUM_REQS - 1:0] grant_unmasked;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:177:9
			reg [NUM_REQS - 1:0] pointer_reg;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:179:9
			wire [NUM_REQS - 1:0] req_masked = requests & pointer_reg;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:181:9
			assign mask_higher_pri_regs[NUM_REQS - 1:1] = mask_higher_pri_regs[NUM_REQS - 2:0] | req_masked[NUM_REQS - 2:0];
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:182:9
			assign mask_higher_pri_regs[0] = 1'b0;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:183:9
			assign grant_masked[NUM_REQS - 1:0] = req_masked[NUM_REQS - 1:0] & ~mask_higher_pri_regs[NUM_REQS - 1:0];
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:185:9
			assign unmask_higher_pri_regs[NUM_REQS - 1:1] = unmask_higher_pri_regs[NUM_REQS - 2:0] | requests[NUM_REQS - 2:0];
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:186:9
			assign unmask_higher_pri_regs[0] = 1'b0;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:187:9
			assign grant_unmasked[NUM_REQS - 1:0] = requests[NUM_REQS - 1:0] & ~unmask_higher_pri_regs[NUM_REQS - 1:0];
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:189:9
			wire no_req_masked = ~(|req_masked);
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:190:9
			assign grant_onehot = ({NUM_REQS {no_req_masked}} & grant_unmasked) | grant_masked;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:192:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:193:7
				if (reset)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:194:5
					pointer_reg <= {NUM_REQS {1'b1}};
				else if (!LOCK_ENABLE || enable)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:196:5
					if (|req_masked)
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:197:21
						pointer_reg <= mask_higher_pri_regs;
					else if (|requests)
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:199:21
						pointer_reg <= unmask_higher_pri_regs;
					else
						// Trace: ../../rtl/libs/VX_rr_arbiter.sv:201:21
						pointer_reg <= pointer_reg;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:206:9
			assign grant_valid = |requests;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:208:9
			VX_onehot_encoder #(.N(NUM_REQS)) onehot_encoder(
				.data_in(grant_onehot),
				.data_out(grant_index)
			);
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:218:9
			reg [LOG_NUM_REQS - 1:0] grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:219:9
			reg [NUM_REQS - 1:0] grant_onehot_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:220:9
			reg [NUM_REQS - 1:0] state;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:222:9
			always @(*) begin
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:223:13
				grant_index_r = 1'sbx;
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:224:13
				grant_onehot_r = 1'sbx;
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:225:13
				begin : sv2v_autoblock_1
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:225:18
					integer i;
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:225:18
					for (i = 0; i < NUM_REQS; i = i + 1)
						begin
							// Trace: ../../rtl/libs/VX_rr_arbiter.sv:226:17
							begin : sv2v_autoblock_2
								// Trace: ../../rtl/libs/VX_rr_arbiter.sv:226:22
								integer j;
								// Trace: ../../rtl/libs/VX_rr_arbiter.sv:226:22
								for (j = 0; j < NUM_REQS; j = j + 1)
									begin
										// Trace: ../../rtl/libs/VX_rr_arbiter.sv:227:21
										if (state[i] && requests[(j + 1) % NUM_REQS]) begin
											// Trace: ../../rtl/libs/VX_rr_arbiter.sv:228:25
											grant_index_r = sv2v_cast_76B5F_signed((j + 1) % NUM_REQS);
											// Trace: ../../rtl/libs/VX_rr_arbiter.sv:229:25
											grant_onehot_r = 1'sb0;
											// Trace: ../../rtl/libs/VX_rr_arbiter.sv:230:25
											grant_onehot_r[(j + 1) % NUM_REQS] = 1;
										end
									end
							end
						end
				end
			end
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:236:9
			always @(posedge clk)
				// Trace: ../../rtl/libs/VX_rr_arbiter.sv:237:13
				if (reset)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:238:17
					state <= 0;
				else if (!LOCK_ENABLE || enable)
					// Trace: ../../rtl/libs/VX_rr_arbiter.sv:240:17
					state <= grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:244:9
			assign grant_index = grant_index_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:245:9
			assign grant_onehot = grant_onehot_r;
			// Trace: ../../rtl/libs/VX_rr_arbiter.sv:246:9
			assign grant_valid = |requests;
		end
	endgenerate
endmodule
module VX_scan (
	data_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_scan.sv:8:15
	parameter N = 1;
	// Trace: ../../rtl/libs/VX_scan.sv:9:15
	parameter OP = 0;
	// Trace: ../../rtl/libs/VX_scan.sv:10:15
	parameter REVERSE = 0;
	// Trace: ../../rtl/libs/VX_scan.sv:12:5
	input wire [N - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_scan.sv:13:5
	output wire [N - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_scan.sv:17:5
	localparam LOGN = $clog2(N);
	// Trace: ../../rtl/libs/VX_scan.sv:19:5
	wire [(LOGN >= 0 ? ((LOGN + 1) * N) - 1 : ((1 - LOGN) * N) + ((LOGN * N) - 1)):(LOGN >= 0 ? 0 : LOGN * N)] t;
	// Trace: ../../rtl/libs/VX_scan.sv:22:5
	generate
		if (REVERSE) begin : genblk1
			// Trace: ../../rtl/libs/VX_scan.sv:23:9
			assign t[(LOGN >= 0 ? 0 : LOGN) * N+:N] = data_in;
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_scan.sv:25:9
			function automatic [N - 1:0] _sv2v_strm_F2A76;
				input reg [(0 + N) - 1:0] inp;
				reg [(0 + N) - 1:0] _sv2v_strm_55E18_inp;
				reg [(0 + N) - 1:0] _sv2v_strm_55E18_out;
				integer _sv2v_strm_55E18_idx;
				begin
					_sv2v_strm_55E18_inp = {inp};
					for (_sv2v_strm_55E18_idx = 0; _sv2v_strm_55E18_idx <= ((0 + N) - 1); _sv2v_strm_55E18_idx = _sv2v_strm_55E18_idx + 1)
						_sv2v_strm_55E18_out[((0 + N) - 1) - _sv2v_strm_55E18_idx-:1] = _sv2v_strm_55E18_inp[_sv2v_strm_55E18_idx+:1];
					_sv2v_strm_F2A76 = ((0 + N) <= N ? _sv2v_strm_55E18_out << (N - (0 + N)) : _sv2v_strm_55E18_out >> ((0 + N) - N));
				end
			endfunction
			assign t[(LOGN >= 0 ? 0 : LOGN) * N+:N] = _sv2v_strm_F2A76({data_in});
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_scan.sv:29:5
	function automatic [N - 1:0] sv2v_cast_AC047;
		input reg [N - 1:0] inp;
		sv2v_cast_AC047 = inp;
	endfunction
	generate
		if ((N == 2) && (OP == 1)) begin : genblk2
			// Trace: ../../rtl/libs/VX_scan.sv:30:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 1], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 1-:2]};
		end
		else if ((N == 3) && (OP == 1)) begin : genblk2
			// Trace: ../../rtl/libs/VX_scan.sv:32:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 2-:2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 2-:3]};
		end
		else if ((N == 4) && (OP == 1)) begin : genblk2
			// Trace: ../../rtl/libs/VX_scan.sv:34:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 3], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:3], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:4]};
		end
		else begin : genblk2
			// Trace: ../../rtl/libs/VX_scan.sv:37:9
			wire [N - 1:0] fill;
			genvar i;
			for (i = 0; i < LOGN; i = i + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_scan.sv:39:13
				wire [N - 1:0] shifted = sv2v_cast_AC047({fill, t[(LOGN >= 0 ? i : LOGN - i) * N+:N]} >> (1 << i));
				if (OP == 0) begin : genblk1
					// Trace: ../../rtl/libs/VX_scan.sv:41:11
					assign fill = {N {1'b0}};
					// Trace: ../../rtl/libs/VX_scan.sv:42:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] ^ shifted;
				end
				else if (OP == 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_scan.sv:44:11
					assign fill = {N {1'b1}};
					// Trace: ../../rtl/libs/VX_scan.sv:45:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] & shifted;
				end
				else if (OP == 2) begin : genblk1
					// Trace: ../../rtl/libs/VX_scan.sv:47:11
					assign fill = {N {1'b0}};
					// Trace: ../../rtl/libs/VX_scan.sv:48:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] | shifted;
				end
			end
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_scan.sv:54:5
	generate
		if (REVERSE) begin : genblk3
			// Trace: ../../rtl/libs/VX_scan.sv:55:9
			assign data_out = t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N];
		end
		else begin : genblk3
			genvar i;
			for (i = 0; i < N; i = i + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_scan.sv:58:13
				assign data_out[i] = t[((LOGN >= 0 ? LOGN : LOGN - LOGN) * N) + ((N - 1) - i)];
			end
		end
	endgenerate
endmodule
module VX_scope (
	clk,
	reset,
	start,
	stop,
	changed,
	data_in,
	bus_in,
	bus_out,
	bus_write,
	bus_read
);
	// Trace: ../../rtl/libs/VX_scope.sv:5:15
	parameter DATAW = 64;
	// Trace: ../../rtl/libs/VX_scope.sv:6:15
	parameter BUSW = 64;
	// Trace: ../../rtl/libs/VX_scope.sv:7:15
	parameter SIZE = 16;
	// Trace: ../../rtl/libs/VX_scope.sv:8:15
	parameter UPDW = 1;
	// Trace: ../../rtl/libs/VX_scope.sv:9:15
	parameter DELTAW = 16;
	// Trace: ../../rtl/libs/VX_scope.sv:11:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_scope.sv:12:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_scope.sv:13:5
	input wire start;
	// Trace: ../../rtl/libs/VX_scope.sv:14:5
	input wire stop;
	// Trace: ../../rtl/libs/VX_scope.sv:15:5
	input wire changed;
	// Trace: ../../rtl/libs/VX_scope.sv:16:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_scope.sv:17:5
	input wire [BUSW - 1:0] bus_in;
	// Trace: ../../rtl/libs/VX_scope.sv:18:5
	output wire [BUSW - 1:0] bus_out;
	// Trace: ../../rtl/libs/VX_scope.sv:19:5
	input wire bus_write;
	// Trace: ../../rtl/libs/VX_scope.sv:20:5
	input wire bus_read;
	// Trace: ../../rtl/libs/VX_scope.sv:22:5
	localparam UPDW_ENABLE = UPDW != 0;
	// Trace: ../../rtl/libs/VX_scope.sv:23:5
	localparam MAX_DELTA = (2 ** DELTAW) - 1;
	// Trace: ../../rtl/libs/VX_scope.sv:25:5
	localparam CMD_GET_VALID = 3'd0;
	// Trace: ../../rtl/libs/VX_scope.sv:26:5
	localparam CMD_GET_DATA = 3'd1;
	// Trace: ../../rtl/libs/VX_scope.sv:27:5
	localparam CMD_GET_WIDTH = 3'd2;
	// Trace: ../../rtl/libs/VX_scope.sv:28:5
	localparam CMD_GET_COUNT = 3'd3;
	// Trace: ../../rtl/libs/VX_scope.sv:29:5
	localparam CMD_SET_START = 3'd4;
	// Trace: ../../rtl/libs/VX_scope.sv:30:5
	localparam CMD_SET_STOP = 3'd5;
	// Trace: ../../rtl/libs/VX_scope.sv:31:5
	localparam CMD_GET_OFFSET = 3'd6;
	// Trace: ../../rtl/libs/VX_scope.sv:33:5
	localparam GET_VALID = 3'd0;
	// Trace: ../../rtl/libs/VX_scope.sv:34:5
	localparam GET_DATA = 3'd1;
	// Trace: ../../rtl/libs/VX_scope.sv:35:5
	localparam GET_WIDTH = 3'd2;
	// Trace: ../../rtl/libs/VX_scope.sv:36:5
	localparam GET_COUNT = 3'd3;
	// Trace: ../../rtl/libs/VX_scope.sv:37:5
	localparam GET_OFFSET = 3'd6;
	// Trace: ../../rtl/libs/VX_scope.sv:39:22
	reg [DATAW - 1:0] data_store [SIZE - 1:0];
	// Trace: ../../rtl/libs/VX_scope.sv:40:22
	reg [DELTAW - 1:0] delta_store [SIZE - 1:0];
	// Trace: ../../rtl/libs/VX_scope.sv:42:5
	reg [UPDW - 1:0] prev_trigger_id;
	// Trace: ../../rtl/libs/VX_scope.sv:43:5
	reg [DELTAW - 1:0] delta;
	// Trace: ../../rtl/libs/VX_scope.sv:44:5
	reg [BUSW - 1:0] bus_out_r;
	// Trace: ../../rtl/libs/VX_scope.sv:45:5
	reg [63:0] timestamp;
	reg [63:0] start_time;
	// Trace: ../../rtl/libs/VX_scope.sv:47:5
	reg [$clog2(SIZE) - 1:0] raddr;
	reg [$clog2(SIZE) - 1:0] waddr;
	reg [$clog2(SIZE) - 1:0] waddr_end;
	// Trace: ../../rtl/libs/VX_scope.sv:49:5
	reg [(DATAW > 1 ? $clog2(DATAW) : 1) - 1:0] read_offset;
	// Trace: ../../rtl/libs/VX_scope.sv:51:5
	reg cmd_start;
	reg started;
	reg start_wait;
	reg recording;
	reg data_valid;
	reg read_delta;
	reg delta_flush;
	// Trace: ../../rtl/libs/VX_scope.sv:53:5
	reg [BUSW - 3:0] delay_val;
	reg [BUSW - 3:0] delay_cntr;
	// Trace: ../../rtl/libs/VX_scope.sv:55:5
	reg [2:0] get_cmd;
	// Trace: ../../rtl/libs/VX_scope.sv:56:5
	wire [2:0] cmd_type;
	// Trace: ../../rtl/libs/VX_scope.sv:57:5
	wire [BUSW - 4:0] cmd_data;
	// Trace: ../../rtl/libs/VX_scope.sv:58:5
	assign {cmd_data, cmd_type} = bus_in;
	// Trace: ../../rtl/libs/VX_scope.sv:60:5
	wire [UPDW - 1:0] trigger_id = data_in[UPDW - 1:0];
	// Trace: ../../rtl/libs/VX_scope.sv:62:5
	function automatic [2:0] sv2v_cast_796CB;
		input reg [2:0] inp;
		sv2v_cast_796CB = inp;
	endfunction
	function automatic signed [$clog2(SIZE) - 1:0] sv2v_cast_088D1_signed;
		input reg signed [$clog2(SIZE) - 1:0] inp;
		sv2v_cast_088D1_signed = inp;
	endfunction
	function automatic [((BUSW - 3) >= 0 ? BUSW - 2 : 4 - BUSW) - 1:0] sv2v_cast_E8B95;
		input reg [((BUSW - 3) >= 0 ? BUSW - 2 : 4 - BUSW) - 1:0] inp;
		sv2v_cast_E8B95 = inp;
	endfunction
	function automatic [$clog2(SIZE) - 1:0] sv2v_cast_088D1;
		input reg [$clog2(SIZE) - 1:0] inp;
		sv2v_cast_088D1 = inp;
	endfunction
	function automatic signed [DELTAW - 1:0] sv2v_cast_B4011_signed;
		input reg signed [DELTAW - 1:0] inp;
		sv2v_cast_B4011_signed = inp;
	endfunction
	function automatic signed [(DATAW > 1 ? $clog2(DATAW) : 1) - 1:0] sv2v_cast_11141_signed;
		input reg signed [(DATAW > 1 ? $clog2(DATAW) : 1) - 1:0] inp;
		sv2v_cast_11141_signed = inp;
	endfunction
	always @(posedge clk) begin
		// Trace: ../../rtl/libs/VX_scope.sv:63:9
		if (reset) begin
			// Trace: ../../rtl/libs/VX_scope.sv:64:13
			get_cmd <= sv2v_cast_796CB(CMD_GET_VALID);
			// Trace: ../../rtl/libs/VX_scope.sv:65:13
			raddr <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:66:13
			waddr <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:67:13
			waddr_end <= sv2v_cast_088D1_signed(SIZE - 1);
			// Trace: ../../rtl/libs/VX_scope.sv:68:13
			cmd_start <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:69:13
			started <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:70:13
			start_wait <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:71:13
			recording <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:72:13
			delay_val <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:73:13
			delay_cntr <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:74:13
			delta <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:75:13
			delta_flush <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:76:13
			prev_trigger_id <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:77:13
			read_offset <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:78:13
			read_delta <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:79:13
			data_valid <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:80:13
			timestamp <= 0;
			// Trace: ../../rtl/libs/VX_scope.sv:81:13
			start_time <= 0;
		end
		else begin
			// Trace: ../../rtl/libs/VX_scope.sv:84:13
			timestamp <= timestamp + 1;
			// Trace: ../../rtl/libs/VX_scope.sv:86:13
			if (bus_write)
				// Trace: ../../rtl/libs/VX_scope.sv:87:17
				case (cmd_type)
					CMD_GET_VALID, CMD_GET_DATA, CMD_GET_WIDTH, CMD_GET_OFFSET, CMD_GET_COUNT:
						// Trace: ../../rtl/libs/VX_scope.sv:92:36
						get_cmd <= sv2v_cast_796CB(cmd_type);
					CMD_SET_START: begin
						// Trace: ../../rtl/libs/VX_scope.sv:94:25
						delay_val <= sv2v_cast_E8B95(cmd_data);
						// Trace: ../../rtl/libs/VX_scope.sv:95:25
						cmd_start <= 1;
					end
					CMD_SET_STOP:
						// Trace: ../../rtl/libs/VX_scope.sv:101:25
						waddr_end <= sv2v_cast_088D1(cmd_data);
					default:
						;
				endcase
			if (!started && (start || cmd_start)) begin
				// Trace: ../../rtl/libs/VX_scope.sv:111:17
				started <= 1;
				// Trace: ../../rtl/libs/VX_scope.sv:112:17
				delta_flush <= 1;
				// Trace: ../../rtl/libs/VX_scope.sv:113:17
				if (0 == delay_val) begin
					// Trace: ../../rtl/libs/VX_scope.sv:114:21
					start_wait <= 0;
					// Trace: ../../rtl/libs/VX_scope.sv:115:21
					recording <= 1;
					// Trace: ../../rtl/libs/VX_scope.sv:116:21
					delta <= 0;
					// Trace: ../../rtl/libs/VX_scope.sv:117:21
					delay_cntr <= 0;
					// Trace: ../../rtl/libs/VX_scope.sv:118:21
					start_time <= timestamp;
				end
				else begin
					// Trace: ../../rtl/libs/VX_scope.sv:123:21
					start_wait <= 1;
					// Trace: ../../rtl/libs/VX_scope.sv:124:21
					delay_cntr <= delay_val;
				end
			end
			if (start_wait) begin
				// Trace: ../../rtl/libs/VX_scope.sv:129:17
				delay_cntr <= delay_cntr - 1;
				// Trace: ../../rtl/libs/VX_scope.sv:130:17
				if (1 == delay_cntr) begin
					// Trace: ../../rtl/libs/VX_scope.sv:131:21
					start_wait <= 0;
					// Trace: ../../rtl/libs/VX_scope.sv:132:21
					recording <= 1;
					// Trace: ../../rtl/libs/VX_scope.sv:133:21
					delta <= 0;
					// Trace: ../../rtl/libs/VX_scope.sv:134:21
					start_time <= timestamp;
				end
			end
			if (recording) begin
				// Trace: ../../rtl/libs/VX_scope.sv:142:17
				if (UPDW_ENABLE) begin
					// Trace: ../../rtl/libs/VX_scope.sv:143:21
					if ((delta_flush || changed) || (trigger_id != prev_trigger_id)) begin
						// Trace: ../../rtl/libs/VX_scope.sv:146:25
						delta_store[waddr] <= delta;
						// Trace: ../../rtl/libs/VX_scope.sv:147:25
						data_store[waddr] <= data_in;
						// Trace: ../../rtl/libs/VX_scope.sv:148:25
						waddr <= waddr + sv2v_cast_088D1_signed(1);
						// Trace: ../../rtl/libs/VX_scope.sv:149:25
						delta <= 0;
						// Trace: ../../rtl/libs/VX_scope.sv:150:25
						delta_flush <= 0;
					end
					else begin
						// Trace: ../../rtl/libs/VX_scope.sv:152:25
						delta <= delta + sv2v_cast_B4011_signed(1);
						// Trace: ../../rtl/libs/VX_scope.sv:153:25
						delta_flush <= delta == (MAX_DELTA - 1);
					end
					// Trace: ../../rtl/libs/VX_scope.sv:155:21
					prev_trigger_id <= trigger_id;
				end
				else begin
					// Trace: ../../rtl/libs/VX_scope.sv:157:21
					delta_store[waddr] <= 0;
					// Trace: ../../rtl/libs/VX_scope.sv:158:21
					data_store[waddr] <= data_in;
					// Trace: ../../rtl/libs/VX_scope.sv:159:21
					waddr <= waddr + 1;
				end
				if (stop || (waddr >= waddr_end)) begin
					// Trace: ../../rtl/libs/VX_scope.sv:167:21
					waddr <= waddr;
					// Trace: ../../rtl/libs/VX_scope.sv:168:21
					recording <= 0;
					// Trace: ../../rtl/libs/VX_scope.sv:169:21
					data_valid <= 1;
					// Trace: ../../rtl/libs/VX_scope.sv:170:21
					read_delta <= 1;
				end
			end
			if ((bus_read && (get_cmd == GET_DATA)) && data_valid)
				// Trace: ../../rtl/libs/VX_scope.sv:177:17
				if (read_delta)
					// Trace: ../../rtl/libs/VX_scope.sv:178:21
					read_delta <= 0;
				else
					// Trace: ../../rtl/libs/VX_scope.sv:180:21
					if (DATAW > BUSW) begin
						begin
							// Trace: ../../rtl/libs/VX_scope.sv:181:25
							if (read_offset < sv2v_cast_11141_signed(DATAW - BUSW))
								// Trace: ../../rtl/libs/VX_scope.sv:182:29
								read_offset <= read_offset + sv2v_cast_11141_signed(BUSW);
							else begin
								// Trace: ../../rtl/libs/VX_scope.sv:184:29
								raddr <= raddr + sv2v_cast_088D1_signed(1);
								// Trace: ../../rtl/libs/VX_scope.sv:185:29
								read_offset <= 0;
								// Trace: ../../rtl/libs/VX_scope.sv:186:29
								read_delta <= 1;
								// Trace: ../../rtl/libs/VX_scope.sv:187:29
								if (raddr == waddr)
									// Trace: ../../rtl/libs/VX_scope.sv:188:33
									data_valid <= 0;
							end
						end
					end
					else begin
						// Trace: ../../rtl/libs/VX_scope.sv:192:25
						raddr <= raddr + 1;
						// Trace: ../../rtl/libs/VX_scope.sv:193:25
						read_delta <= 1;
						// Trace: ../../rtl/libs/VX_scope.sv:194:25
						if (raddr == waddr)
							// Trace: ../../rtl/libs/VX_scope.sv:195:29
							data_valid <= 0;
					end
		end
		if (recording)
			// Trace: ../../rtl/libs/VX_scope.sv:203:13
			if (UPDW_ENABLE) begin
				begin
					// Trace: ../../rtl/libs/VX_scope.sv:204:17
					if ((delta_flush || changed) || (trigger_id != prev_trigger_id)) begin
						// Trace: ../../rtl/libs/VX_scope.sv:207:21
						delta_store[waddr] <= delta;
						// Trace: ../../rtl/libs/VX_scope.sv:208:21
						data_store[waddr] <= data_in;
					end
				end
			end
			else begin
				// Trace: ../../rtl/libs/VX_scope.sv:211:17
				delta_store[waddr] <= 0;
				// Trace: ../../rtl/libs/VX_scope.sv:212:17
				data_store[waddr] <= data_in;
			end
	end
	// Trace: ../../rtl/libs/VX_scope.sv:217:5
	function automatic [BUSW - 1:0] sv2v_cast_39A33;
		input reg [BUSW - 1:0] inp;
		sv2v_cast_39A33 = inp;
	endfunction
	function automatic signed [BUSW - 1:0] sv2v_cast_39A33_signed;
		input reg signed [BUSW - 1:0] inp;
		sv2v_cast_39A33_signed = inp;
	endfunction
	always @(*)
		// Trace: ../../rtl/libs/VX_scope.sv:218:9
		case (get_cmd)
			GET_VALID:
				// Trace: ../../rtl/libs/VX_scope.sv:219:25
				bus_out_r = sv2v_cast_39A33(data_valid);
			GET_WIDTH:
				// Trace: ../../rtl/libs/VX_scope.sv:220:25
				bus_out_r = sv2v_cast_39A33_signed(DATAW);
			GET_COUNT:
				// Trace: ../../rtl/libs/VX_scope.sv:221:25
				bus_out_r = sv2v_cast_39A33(waddr) + sv2v_cast_39A33_signed(1);
			GET_OFFSET:
				// Trace: ../../rtl/libs/VX_scope.sv:222:25
				bus_out_r = sv2v_cast_39A33(start_time);
			GET_DATA:
				// Trace: ../../rtl/libs/VX_scope.sv:224:25
				bus_out_r = (read_delta ? sv2v_cast_39A33(delta_store[raddr]) : sv2v_cast_39A33(data_store[raddr] >> read_offset));
			default:
				// Trace: ../../rtl/libs/VX_scope.sv:226:25
				bus_out_r = 0;
		endcase
	// Trace: ../../rtl/libs/VX_scope.sv:230:5
	assign bus_out = bus_out_r;
endmodule
module VX_serial_div (
	clk,
	reset,
	valid_in,
	ready_in,
	numer,
	denom,
	signed_mode,
	tag_in,
	quotient,
	remainder,
	ready_out,
	valid_out,
	tag_out
);
	// Trace: ../../rtl/libs/VX_serial_div.sv:5:15
	parameter WIDTHN = 1;
	// Trace: ../../rtl/libs/VX_serial_div.sv:6:15
	parameter WIDTHD = 1;
	// Trace: ../../rtl/libs/VX_serial_div.sv:7:15
	parameter WIDTHQ = 1;
	// Trace: ../../rtl/libs/VX_serial_div.sv:8:15
	parameter WIDTHR = 1;
	// Trace: ../../rtl/libs/VX_serial_div.sv:9:15
	parameter LANES = 1;
	// Trace: ../../rtl/libs/VX_serial_div.sv:10:15
	parameter TAGW = 1;
	// Trace: ../../rtl/libs/VX_serial_div.sv:12:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_serial_div.sv:13:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_serial_div.sv:15:5
	input wire valid_in;
	// Trace: ../../rtl/libs/VX_serial_div.sv:16:5
	output wire ready_in;
	// Trace: ../../rtl/libs/VX_serial_div.sv:17:5
	input wire [(LANES * WIDTHN) - 1:0] numer;
	// Trace: ../../rtl/libs/VX_serial_div.sv:18:5
	input wire [(LANES * WIDTHD) - 1:0] denom;
	// Trace: ../../rtl/libs/VX_serial_div.sv:19:5
	input wire signed_mode;
	// Trace: ../../rtl/libs/VX_serial_div.sv:20:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/libs/VX_serial_div.sv:22:5
	output wire [(LANES * WIDTHQ) - 1:0] quotient;
	// Trace: ../../rtl/libs/VX_serial_div.sv:23:5
	output wire [(LANES * WIDTHR) - 1:0] remainder;
	// Trace: ../../rtl/libs/VX_serial_div.sv:24:5
	input wire ready_out;
	// Trace: ../../rtl/libs/VX_serial_div.sv:25:5
	output wire valid_out;
	// Trace: ../../rtl/libs/VX_serial_div.sv:26:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/libs/VX_serial_div.sv:28:5
	localparam MIN_ND = (WIDTHN < WIDTHD ? WIDTHN : WIDTHD);
	// Trace: ../../rtl/libs/VX_serial_div.sv:29:5
	localparam CNTRW = $clog2(WIDTHN + 1);
	// Trace: ../../rtl/libs/VX_serial_div.sv:31:5
	reg [((WIDTHN + MIN_ND) >= 0 ? (LANES * ((WIDTHN + MIN_ND) + 1)) - 1 : (LANES * (1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) - 1)):((WIDTHN + MIN_ND) >= 0 ? 0 : (WIDTHN + MIN_ND) + 0)] working;
	// Trace: ../../rtl/libs/VX_serial_div.sv:32:5
	reg [(LANES * WIDTHD) - 1:0] denom_r;
	// Trace: ../../rtl/libs/VX_serial_div.sv:34:5
	wire [(LANES * WIDTHN) - 1:0] numer_qual;
	// Trace: ../../rtl/libs/VX_serial_div.sv:35:5
	wire [(LANES * WIDTHD) - 1:0] denom_qual;
	// Trace: ../../rtl/libs/VX_serial_div.sv:36:5
	wire [(WIDTHD >= 0 ? (LANES * (WIDTHD + 1)) - 1 : (LANES * (1 - WIDTHD)) + (WIDTHD - 1)):(WIDTHD >= 0 ? 0 : WIDTHD + 0)] sub_result;
	// Trace: ../../rtl/libs/VX_serial_div.sv:38:5
	reg [LANES - 1:0] inv_quot;
	reg [LANES - 1:0] inv_rem;
	// Trace: ../../rtl/libs/VX_serial_div.sv:40:5
	reg [CNTRW - 1:0] cntr;
	// Trace: ../../rtl/libs/VX_serial_div.sv:41:5
	reg is_busy;
	// Trace: ../../rtl/libs/VX_serial_div.sv:43:5
	reg [TAGW - 1:0] tag_r;
	// Trace: ../../rtl/libs/VX_serial_div.sv:45:5
	wire done = ~(|cntr);
	// Trace: ../../rtl/libs/VX_serial_div.sv:47:5
	wire push = valid_in && ready_in;
	// Trace: ../../rtl/libs/VX_serial_div.sv:48:5
	wire pop = valid_out && ready_out;
	// Trace: ../../rtl/libs/VX_serial_div.sv:50:5
	genvar i;
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_serial_div.sv:51:9
			wire negate_numer = signed_mode && numer[(i * WIDTHN) + (WIDTHN - 1)];
			// Trace: ../../rtl/libs/VX_serial_div.sv:52:9
			wire negate_denom = signed_mode && denom[(i * WIDTHD) + (WIDTHD - 1)];
			// Trace: ../../rtl/libs/VX_serial_div.sv:53:9
			assign numer_qual[i * WIDTHN+:WIDTHN] = (negate_numer ? -$signed(numer[i * WIDTHN+:WIDTHN]) : numer[i * WIDTHN+:WIDTHN]);
			// Trace: ../../rtl/libs/VX_serial_div.sv:54:9
			assign denom_qual[i * WIDTHD+:WIDTHD] = (negate_denom ? -$signed(denom[i * WIDTHD+:WIDTHD]) : denom[i * WIDTHD+:WIDTHD]);
			// Trace: ../../rtl/libs/VX_serial_div.sv:55:9
			assign sub_result[(WIDTHD >= 0 ? 0 : WIDTHD) + (i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD))+:(WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)] = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1))) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1)-:((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)] - denom_r[i * WIDTHD+:WIDTHD];
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_serial_div.sv:58:5
	function automatic signed [CNTRW - 1:0] sv2v_cast_A86AD_signed;
		input reg signed [CNTRW - 1:0] inp;
		sv2v_cast_A86AD_signed = inp;
	endfunction
	always @(posedge clk) begin
		// Trace: ../../rtl/libs/VX_serial_div.sv:59:9
		if (reset) begin
			// Trace: ../../rtl/libs/VX_serial_div.sv:60:13
			cntr <= 0;
			// Trace: ../../rtl/libs/VX_serial_div.sv:61:13
			is_busy <= 0;
		end
		else begin
			// Trace: ../../rtl/libs/VX_serial_div.sv:63:13
			if (push) begin
				// Trace: ../../rtl/libs/VX_serial_div.sv:64:17
				cntr <= WIDTHN;
				// Trace: ../../rtl/libs/VX_serial_div.sv:65:17
				is_busy <= 1;
			end
			else if (!done)
				// Trace: ../../rtl/libs/VX_serial_div.sv:67:17
				cntr <= cntr - sv2v_cast_A86AD_signed(1);
			if (pop)
				// Trace: ../../rtl/libs/VX_serial_div.sv:70:17
				is_busy <= 0;
		end
		if (push) begin
			// Trace: ../../rtl/libs/VX_serial_div.sv:75:13
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/libs/VX_serial_div.sv:75:18
				integer i;
				// Trace: ../../rtl/libs/VX_serial_div.sv:75:18
				for (i = 0; i < LANES; i = i + 1)
					begin
						// Trace: ../../rtl/libs/VX_serial_div.sv:76:17
						working[((WIDTHN + MIN_ND) >= 0 ? 0 : WIDTHN + MIN_ND) + (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND)))+:((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))] <= {{WIDTHD {1'b0}}, numer_qual[i * WIDTHN+:WIDTHN], 1'b0};
						// Trace: ../../rtl/libs/VX_serial_div.sv:77:17
						denom_r[i * WIDTHD+:WIDTHD] <= denom_qual[i * WIDTHD+:WIDTHD];
						// Trace: ../../rtl/libs/VX_serial_div.sv:78:17
						inv_quot[i] <= ((denom[i * WIDTHD+:WIDTHD] != 0) && signed_mode) && (numer[(i * WIDTHN) + 31] ^ denom[(i * WIDTHD) + 31]);
						// Trace: ../../rtl/libs/VX_serial_div.sv:79:17
						inv_rem[i] <= signed_mode && numer[(i * WIDTHN) + 31];
					end
			end
			// Trace: ../../rtl/libs/VX_serial_div.sv:81:13
			tag_r <= tag_in;
		end
		else if (!done)
			// Trace: ../../rtl/libs/VX_serial_div.sv:83:13
			begin : sv2v_autoblock_2
				// Trace: ../../rtl/libs/VX_serial_div.sv:83:18
				integer i;
				// Trace: ../../rtl/libs/VX_serial_div.sv:83:18
				for (i = 0; i < LANES; i = i + 1)
					begin
						// Trace: ../../rtl/libs/VX_serial_div.sv:84:17
						working[((WIDTHN + MIN_ND) >= 0 ? 0 : WIDTHN + MIN_ND) + (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND)))+:((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))] <= (sub_result[(i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD : WIDTHD - WIDTHD)] ? {working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) - 1 : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) - 1 : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) - 1))) + (WIDTHN + MIN_ND)) - 1)-:WIDTHN + MIN_ND], 1'b0} : {sub_result[(WIDTHD >= 0 ? (i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD - 1 : WIDTHD - (WIDTHD - 1)) : (((i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD - 1 : WIDTHD - (WIDTHD - 1))) + WIDTHD) - 1)-:WIDTHD], working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHN - 1 : (WIDTHN + MIN_ND) - (WIDTHN - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHN - 1 : (WIDTHN + MIN_ND) - (WIDTHN - 1))) + WIDTHN) - 1)-:WIDTHN], 1'b1});
					end
			end
	end
	// Trace: ../../rtl/libs/VX_serial_div.sv:90:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk2
			// Trace: ../../rtl/libs/VX_serial_div.sv:91:9
			wire [WIDTHQ - 1:0] q = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHQ - 1 : (WIDTHN + MIN_ND) - (WIDTHQ - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHQ - 1 : (WIDTHN + MIN_ND) - (WIDTHQ - 1))) + WIDTHQ) - 1)-:WIDTHQ];
			// Trace: ../../rtl/libs/VX_serial_div.sv:92:9
			wire [WIDTHR - 1:0] r = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1))) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1)-:((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)];
			// Trace: ../../rtl/libs/VX_serial_div.sv:93:9
			assign quotient[i * WIDTHQ+:WIDTHQ] = (inv_quot[i] ? -$signed(q) : q);
			// Trace: ../../rtl/libs/VX_serial_div.sv:94:9
			assign remainder[i * WIDTHR+:WIDTHR] = (inv_rem[i] ? -$signed(r) : r);
		end
	endgenerate
	// Trace: ../../rtl/libs/VX_serial_div.sv:97:5
	assign ready_in = !is_busy;
	// Trace: ../../rtl/libs/VX_serial_div.sv:98:5
	assign tag_out = tag_r;
	// Trace: ../../rtl/libs/VX_serial_div.sv:99:5
	assign valid_out = is_busy && done;
endmodule
module VX_shift_register_nr (
	clk,
	enable,
	data_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_shift_register.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:6:15
	parameter DEPTH = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:7:15
	parameter NTAPS = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:8:15
	parameter DEPTHW = $clog2(DEPTH);
	// Trace: ../../rtl/libs/VX_shift_register.sv:9:15
	function automatic signed [DEPTHW - 1:0] sv2v_cast_5F7C4_signed;
		input reg signed [DEPTHW - 1:0] inp;
		sv2v_cast_5F7C4_signed = inp;
	endfunction
	parameter [(DEPTHW * NTAPS) - 1:0] TAPS = {NTAPS {sv2v_cast_5F7C4_signed(DEPTH - 1)}};
	// Trace: ../../rtl/libs/VX_shift_register.sv:11:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_shift_register.sv:12:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_shift_register.sv:13:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_shift_register.sv:14:5
	output wire [(NTAPS * DATAW) - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_shift_register.sv:16:5
	reg [(DEPTH * DATAW) - 1:0] entries;
	// Trace: ../../rtl/libs/VX_shift_register.sv:18:5
	always @(posedge clk)
		// Trace: ../../rtl/libs/VX_shift_register.sv:19:9
		if (enable) begin
			// Trace: ../../rtl/libs/VX_shift_register.sv:20:13
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/libs/VX_shift_register.sv:20:18
				integer i;
				// Trace: ../../rtl/libs/VX_shift_register.sv:20:18
				for (i = DEPTH - 1; i > 0; i = i - 1)
					begin
						// Trace: ../../rtl/libs/VX_shift_register.sv:21:17
						entries[i * DATAW+:DATAW] <= entries[(i - 1) * DATAW+:DATAW];
					end
			end
			// Trace: ../../rtl/libs/VX_shift_register.sv:22:13
			entries[0+:DATAW] <= data_in;
		end
	// Trace: ../../rtl/libs/VX_shift_register.sv:26:5
	genvar i;
	generate
		for (i = 0; i < NTAPS; i = i + 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_shift_register.sv:27:9
			assign data_out[i * DATAW+:DATAW] = entries[TAPS[i * DEPTHW+:DEPTHW] * DATAW+:DATAW];
		end
	endgenerate
endmodule
module VX_shift_register_wr (
	clk,
	reset,
	enable,
	data_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_shift_register.sv:33:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:34:15
	parameter DEPTH = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:35:15
	parameter NTAPS = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:36:15
	parameter DEPTHW = $clog2(DEPTH);
	// Trace: ../../rtl/libs/VX_shift_register.sv:37:15
	function automatic signed [DEPTHW - 1:0] sv2v_cast_5F7C4_signed;
		input reg signed [DEPTHW - 1:0] inp;
		sv2v_cast_5F7C4_signed = inp;
	endfunction
	parameter [(DEPTHW * NTAPS) - 1:0] TAPS = {NTAPS {sv2v_cast_5F7C4_signed(DEPTH - 1)}};
	// Trace: ../../rtl/libs/VX_shift_register.sv:39:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_shift_register.sv:40:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_shift_register.sv:41:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_shift_register.sv:42:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_shift_register.sv:43:5
	output wire [(NTAPS * DATAW) - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_shift_register.sv:45:5
	reg [(DEPTH * DATAW) - 1:0] entries;
	// Trace: ../../rtl/libs/VX_shift_register.sv:47:5
	always @(posedge clk)
		// Trace: ../../rtl/libs/VX_shift_register.sv:48:9
		if (reset)
			// Trace: ../../rtl/libs/VX_shift_register.sv:49:13
			entries <= 1'sb0;
		else if (enable) begin
			// Trace: ../../rtl/libs/VX_shift_register.sv:51:13
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/libs/VX_shift_register.sv:51:18
				integer i;
				// Trace: ../../rtl/libs/VX_shift_register.sv:51:18
				for (i = DEPTH - 1; i > 0; i = i - 1)
					begin
						// Trace: ../../rtl/libs/VX_shift_register.sv:52:17
						entries[i * DATAW+:DATAW] <= entries[(i - 1) * DATAW+:DATAW];
					end
			end
			// Trace: ../../rtl/libs/VX_shift_register.sv:53:13
			entries[0+:DATAW] <= data_in;
		end
	// Trace: ../../rtl/libs/VX_shift_register.sv:57:5
	genvar i;
	generate
		for (i = 0; i < NTAPS; i = i + 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_shift_register.sv:58:9
			assign data_out[i * DATAW+:DATAW] = entries[TAPS[i * DEPTHW+:DEPTHW] * DATAW+:DATAW];
		end
	endgenerate
endmodule
module VX_shift_register (
	clk,
	reset,
	enable,
	data_in,
	data_out
);
	// Trace: ../../rtl/libs/VX_shift_register.sv:64:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:65:15
	parameter RESETW = 0;
	// Trace: ../../rtl/libs/VX_shift_register.sv:66:15
	parameter DEPTH = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:67:15
	parameter NTAPS = 1;
	// Trace: ../../rtl/libs/VX_shift_register.sv:68:15
	parameter DEPTHW = $clog2(DEPTH);
	// Trace: ../../rtl/libs/VX_shift_register.sv:69:15
	function automatic signed [DEPTHW - 1:0] sv2v_cast_5F7C4_signed;
		input reg signed [DEPTHW - 1:0] inp;
		sv2v_cast_5F7C4_signed = inp;
	endfunction
	parameter [(DEPTHW * NTAPS) - 1:0] TAPS = {NTAPS {sv2v_cast_5F7C4_signed(DEPTH - 1)}};
	// Trace: ../../rtl/libs/VX_shift_register.sv:71:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_shift_register.sv:72:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_shift_register.sv:73:5
	input wire enable;
	// Trace: ../../rtl/libs/VX_shift_register.sv:74:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_shift_register.sv:75:5
	output wire [(NTAPS * DATAW) - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_shift_register.sv:77:5
	generate
		if (RESETW != 0) begin : genblk1
			if (RESETW == DATAW) begin : genblk1
				// Trace: ../../rtl/libs/VX_shift_register.sv:80:13
				VX_shift_register_wr #(
					.DATAW(DATAW),
					.DEPTH(DEPTH),
					.NTAPS(NTAPS),
					.TAPS(TAPS)
				) sr(
					.clk(clk),
					.reset(reset),
					.enable(enable),
					.data_in(data_in),
					.data_out(data_out)
				);
			end
			else begin : genblk1
				// Trace: ../../rtl/libs/VX_shift_register.sv:95:13
				VX_shift_register_wr #(
					.DATAW(RESETW),
					.DEPTH(DEPTH),
					.NTAPS(NTAPS),
					.TAPS(TAPS)
				) sr_wr(
					.clk(clk),
					.reset(reset),
					.enable(enable),
					.data_in(data_in[DATAW - 1:DATAW - RESETW]),
					.data_out(data_out[DATAW - 1:DATAW - RESETW])
				);
				// Trace: ../../rtl/libs/VX_shift_register.sv:108:13
				VX_shift_register_nr #(
					.DATAW(DATAW - RESETW),
					.DEPTH(DEPTH),
					.NTAPS(NTAPS),
					.TAPS(TAPS)
				) sr_nr(
					.clk(clk),
					.enable(enable),
					.data_in(data_in[(DATAW - RESETW) - 1:0]),
					.data_out(data_out[(DATAW - RESETW) - 1:0])
				);
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_shift_register.sv:126:9
			VX_shift_register_nr #(
				.DATAW(DATAW),
				.DEPTH(DEPTH),
				.NTAPS(NTAPS),
				.TAPS(TAPS)
			) sr(
				.clk(clk),
				.enable(enable),
				.data_in(data_in),
				.data_out(data_out)
			);
		end
	endgenerate
endmodule
module VX_skid_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:6:15
	parameter PASSTHRU = 0;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:7:15
	parameter NOBACKPRESSURE = 0;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:8:15
	parameter OUT_REG = 0;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:10:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:11:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:13:5
	input wire valid_in;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:14:5
	output wire ready_in;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:15:5
	input wire [DATAW - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:17:5
	output wire [DATAW - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:18:5
	input wire ready_out;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:19:5
	output wire valid_out;
	// Trace: ../../rtl/libs/VX_skid_buffer.sv:22:5
	generate
		if (PASSTHRU) begin : genblk1
			// Trace: ../../rtl/libs/VX_skid_buffer.sv:27:9
			assign valid_out = valid_in;
			// Trace: ../../rtl/libs/VX_skid_buffer.sv:28:9
			assign data_out = data_in;
			// Trace: ../../rtl/libs/VX_skid_buffer.sv:29:9
			assign ready_in = ready_out;
		end
		else if (NOBACKPRESSURE) begin : genblk1
			// Trace: ../../rtl/libs/VX_skid_buffer.sv:35:9
			wire stall = valid_out && ~ready_out;
			// Trace: ../../rtl/libs/VX_skid_buffer.sv:37:9
			VX_pipe_register #(
				.DATAW(1 + DATAW),
				.RESETW(1)
			) pipe_reg(
				.clk(clk),
				.reset(reset),
				.enable(!stall),
				.data_in({valid_in, data_in}),
				.data_out({valid_out, data_out})
			);
			// Trace: ../../rtl/libs/VX_skid_buffer.sv:48:9
			assign ready_in = ~stall;
		end
		else begin : genblk1
			if (OUT_REG) begin : genblk1
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:54:13
				reg [DATAW - 1:0] data_out_r;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:55:13
				reg [DATAW - 1:0] buffer;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:56:13
				reg valid_out_r;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:57:13
				reg use_buffer;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:59:13
				wire push = valid_in && ready_in;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:60:13
				wire pop = !valid_out_r || ready_out;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:62:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_skid_buffer.sv:63:17
					if (reset) begin
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:64:21
						valid_out_r <= 0;
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:65:21
						use_buffer <= 0;
					end
					else begin
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:67:21
						if (ready_out)
							// Trace: ../../rtl/libs/VX_skid_buffer.sv:68:25
							use_buffer <= 0;
						else if (valid_in && valid_out_r)
							// Trace: ../../rtl/libs/VX_skid_buffer.sv:70:25
							use_buffer <= 1;
						if (pop)
							// Trace: ../../rtl/libs/VX_skid_buffer.sv:73:25
							valid_out_r <= valid_in || use_buffer;
					end
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:78:13
				always @(posedge clk) begin
					// Trace: ../../rtl/libs/VX_skid_buffer.sv:79:17
					if (push)
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:80:21
						buffer <= data_in;
					if (pop && !use_buffer)
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:83:21
						data_out_r <= data_in;
					else if (ready_out)
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:85:21
						data_out_r <= buffer;
				end
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:89:13
				assign ready_in = !use_buffer;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:90:13
				assign valid_out = valid_out_r;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:91:13
				assign data_out = data_out_r;
			end
			else begin : genblk1
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:95:13
				reg [DATAW - 1:0] shift_reg [1:0];
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:96:13
				reg valid_out_r;
				reg ready_in_r;
				reg rd_ptr_r;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:98:13
				wire push = valid_in && ready_in;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:99:13
				wire pop = valid_out_r && ready_out;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:101:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_skid_buffer.sv:102:17
					if (reset) begin
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:103:21
						valid_out_r <= 0;
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:104:21
						ready_in_r <= 1;
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:105:21
						rd_ptr_r <= 1;
					end
					else begin
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:107:21
						if (push) begin
							begin
								// Trace: ../../rtl/libs/VX_skid_buffer.sv:108:25
								if (!pop) begin
									// Trace: ../../rtl/libs/VX_skid_buffer.sv:109:29
									ready_in_r <= rd_ptr_r;
									// Trace: ../../rtl/libs/VX_skid_buffer.sv:110:29
									valid_out_r <= 1;
								end
							end
						end
						else if (pop) begin
							// Trace: ../../rtl/libs/VX_skid_buffer.sv:113:25
							ready_in_r <= 1;
							// Trace: ../../rtl/libs/VX_skid_buffer.sv:114:25
							valid_out_r <= rd_ptr_r;
						end
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:116:21
						rd_ptr_r <= rd_ptr_r ^ (push ^ pop);
					end
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:120:13
				always @(posedge clk)
					// Trace: ../../rtl/libs/VX_skid_buffer.sv:121:17
					if (push) begin
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:122:21
						shift_reg[1] <= shift_reg[0];
						// Trace: ../../rtl/libs/VX_skid_buffer.sv:123:21
						shift_reg[0] <= data_in;
					end
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:127:13
				assign ready_in = ready_in_r;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:128:13
				assign valid_out = valid_out_r;
				// Trace: ../../rtl/libs/VX_skid_buffer.sv:129:13
				assign data_out = shift_reg[rd_ptr_r];
			end
		end
	endgenerate
endmodule
module VX_sp_ram (
	clk,
	addr,
	wren,
	wdata,
	rdata
);
	// Trace: ../../rtl/libs/VX_sp_ram.sv:5:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:6:15
	parameter SIZE = 1;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:7:15
	parameter BYTEENW = 1;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:8:15
	parameter OUT_REG = 0;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:9:15
	parameter NO_RWCHECK = 0;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:10:15
	parameter LUTRAM = 0;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:11:15
	parameter ADDRW = $clog2(SIZE);
	// Trace: ../../rtl/libs/VX_sp_ram.sv:12:15
	parameter INIT_ENABLE = 0;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:13:15
	parameter INIT_FILE = "";
	// Trace: ../../rtl/libs/VX_sp_ram.sv:14:15
	parameter [DATAW - 1:0] INIT_VALUE = 0;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:16:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:17:5
	input wire [ADDRW - 1:0] addr;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:18:5
	input wire [BYTEENW - 1:0] wren;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:19:5
	input wire [DATAW - 1:0] wdata;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:20:5
	output wire [DATAW - 1:0] rdata;
	// Trace: ../../rtl/libs/VX_sp_ram.sv:37:5
	generate
		if (LUTRAM) begin : genblk1
			if (OUT_REG) begin : genblk1
				// Trace: ../../rtl/libs/VX_sp_ram.sv:39:13
				reg [DATAW - 1:0] rdata_r;
				if (BYTEENW > 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_sp_ram.sv:42:32
					reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:44:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:44:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:44:234
							initial begin : sv2v_autoblock_1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:44:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:44:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:44:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_sp_ram.sv:46:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_sp_ram.sv:47:21
						begin : sv2v_autoblock_2
							// Trace: ../../rtl/libs/VX_sp_ram.sv:47:26
							integer i;
							// Trace: ../../rtl/libs/VX_sp_ram.sv:47:26
							for (i = 0; i < BYTEENW; i = i + 1)
								begin
									// Trace: ../../rtl/libs/VX_sp_ram.sv:48:25
									if (wren[i])
										// Trace: ../../rtl/libs/VX_sp_ram.sv:49:29
										ram[addr][i * 8+:8] <= wdata[i * 8+:8];
								end
						end
						// Trace: ../../rtl/libs/VX_sp_ram.sv:51:21
						rdata_r <= ram[addr];
					end
				end
				else begin : genblk1
					// Trace: ../../rtl/libs/VX_sp_ram.sv:54:32
					reg [DATAW - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:56:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:56:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:56:234
							initial begin : sv2v_autoblock_3
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:56:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:56:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:56:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_sp_ram.sv:58:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_sp_ram.sv:59:21
						if (wren)
							// Trace: ../../rtl/libs/VX_sp_ram.sv:60:25
							ram[addr] <= wdata;
						// Trace: ../../rtl/libs/VX_sp_ram.sv:61:21
						rdata_r <= ram[addr];
					end
				end
				// Trace: ../../rtl/libs/VX_sp_ram.sv:64:13
				assign rdata = rdata_r;
			end
			else begin : genblk1
				if (BYTEENW > 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_sp_ram.sv:67:32
					reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:69:131
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:69:139
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:69:233
							initial begin : sv2v_autoblock_4
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:69:293
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:69:293
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:69:343
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_sp_ram.sv:71:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_sp_ram.sv:72:21
						begin : sv2v_autoblock_5
							// Trace: ../../rtl/libs/VX_sp_ram.sv:72:26
							integer i;
							// Trace: ../../rtl/libs/VX_sp_ram.sv:72:26
							for (i = 0; i < BYTEENW; i = i + 1)
								begin
									// Trace: ../../rtl/libs/VX_sp_ram.sv:73:25
									if (wren[i])
										// Trace: ../../rtl/libs/VX_sp_ram.sv:74:29
										ram[addr][i * 8+:8] <= wdata[i * 8+:8];
								end
						end
					// Trace: ../../rtl/libs/VX_sp_ram.sv:77:17
					assign rdata = ram[addr];
				end
				else begin : genblk1
					// Trace: ../../rtl/libs/VX_sp_ram.sv:79:32
					reg [DATAW - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:81:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:81:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:81:234
							initial begin : sv2v_autoblock_6
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:81:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:81:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:81:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_sp_ram.sv:83:17
					always @(posedge clk)
						// Trace: ../../rtl/libs/VX_sp_ram.sv:84:21
						if (wren)
							// Trace: ../../rtl/libs/VX_sp_ram.sv:85:25
							ram[addr] <= wdata;
					// Trace: ../../rtl/libs/VX_sp_ram.sv:87:17
					assign rdata = ram[addr];
				end
			end
		end
		else begin : genblk1
			if (OUT_REG) begin : genblk1
				// Trace: ../../rtl/libs/VX_sp_ram.sv:92:13
				reg [DATAW - 1:0] rdata_r;
				if (BYTEENW > 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_sp_ram.sv:95:17
					reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:97:132
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:97:140
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:97:234
							initial begin : sv2v_autoblock_7
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:97:294
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:97:294
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:97:344
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_sp_ram.sv:99:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_sp_ram.sv:100:21
						begin : sv2v_autoblock_8
							// Trace: ../../rtl/libs/VX_sp_ram.sv:100:26
							integer i;
							// Trace: ../../rtl/libs/VX_sp_ram.sv:100:26
							for (i = 0; i < BYTEENW; i = i + 1)
								begin
									// Trace: ../../rtl/libs/VX_sp_ram.sv:101:25
									if (wren[i])
										// Trace: ../../rtl/libs/VX_sp_ram.sv:102:29
										ram[addr][i * 8+:8] <= wdata[i * 8+:8];
								end
						end
						// Trace: ../../rtl/libs/VX_sp_ram.sv:104:21
						rdata_r <= ram[addr];
					end
				end
				else begin : genblk1
					// Trace: ../../rtl/libs/VX_sp_ram.sv:107:17
					reg [DATAW - 1:0] ram [SIZE - 1:0];
					if (INIT_ENABLE) begin : genblk1
						if (INIT_FILE != "") begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:109:131
							initial begin
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:109:139
								$readmemh(INIT_FILE, ram);
							end
						end
						else begin : genblk1
							// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:109:233
							initial begin : sv2v_autoblock_9
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:109:293
								integer i;
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:109:293
								for (i = 0; i < SIZE; i = i + 1)
									begin
										// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:109:343
										ram[i] = INIT_VALUE;
									end
							end
						end
					end
					// Trace: ../../rtl/libs/VX_sp_ram.sv:111:17
					always @(posedge clk) begin
						// Trace: ../../rtl/libs/VX_sp_ram.sv:112:21
						if (wren)
							// Trace: ../../rtl/libs/VX_sp_ram.sv:113:25
							ram[addr] <= wdata;
						// Trace: ../../rtl/libs/VX_sp_ram.sv:114:21
						rdata_r <= ram[addr];
					end
				end
				// Trace: ../../rtl/libs/VX_sp_ram.sv:117:13
				assign rdata = rdata_r;
			end
			else begin : genblk1
				if (NO_RWCHECK) begin : genblk1
					if (BYTEENW > 1) begin : genblk1
						// Trace: ../../rtl/libs/VX_sp_ram.sv:121:38
						reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
						if (INIT_ENABLE) begin : genblk1
							if (INIT_FILE != "") begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:123:136
								initial begin
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:123:144
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:123:238
								initial begin : sv2v_autoblock_10
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:123:298
									integer i;
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:123:298
									for (i = 0; i < SIZE; i = i + 1)
										begin
											// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:123:348
											ram[i] = INIT_VALUE;
										end
								end
							end
						end
						// Trace: ../../rtl/libs/VX_sp_ram.sv:125:21
						always @(posedge clk)
							// Trace: ../../rtl/libs/VX_sp_ram.sv:126:25
							begin : sv2v_autoblock_11
								// Trace: ../../rtl/libs/VX_sp_ram.sv:126:30
								integer i;
								// Trace: ../../rtl/libs/VX_sp_ram.sv:126:30
								for (i = 0; i < BYTEENW; i = i + 1)
									begin
										// Trace: ../../rtl/libs/VX_sp_ram.sv:127:29
										if (wren[i])
											// Trace: ../../rtl/libs/VX_sp_ram.sv:128:33
											ram[addr][i * 8+:8] <= wdata[i * 8+:8];
									end
							end
						// Trace: ../../rtl/libs/VX_sp_ram.sv:131:21
						assign rdata = ram[addr];
					end
					else begin : genblk1
						// Trace: ../../rtl/libs/VX_sp_ram.sv:133:38
						reg [DATAW - 1:0] ram [SIZE - 1:0];
						if (INIT_ENABLE) begin : genblk1
							if (INIT_FILE != "") begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:135:136
								initial begin
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:135:144
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:135:238
								initial begin : sv2v_autoblock_12
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:135:298
									integer i;
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:135:298
									for (i = 0; i < SIZE; i = i + 1)
										begin
											// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:135:348
											ram[i] = INIT_VALUE;
										end
								end
							end
						end
						// Trace: ../../rtl/libs/VX_sp_ram.sv:137:21
						always @(posedge clk)
							// Trace: ../../rtl/libs/VX_sp_ram.sv:138:25
							if (wren)
								// Trace: ../../rtl/libs/VX_sp_ram.sv:139:29
								ram[addr] <= wdata;
						// Trace: ../../rtl/libs/VX_sp_ram.sv:141:21
						assign rdata = ram[addr];
					end
				end
				else begin : genblk1
					if (BYTEENW > 1) begin : genblk1
						// Trace: ../../rtl/libs/VX_sp_ram.sv:145:21
						reg [(BYTEENW * 8) - 1:0] ram [SIZE - 1:0];
						if (INIT_ENABLE) begin : genblk1
							if (INIT_FILE != "") begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:147:136
								initial begin
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:147:144
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:147:238
								initial begin : sv2v_autoblock_13
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:147:298
									integer i;
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:147:298
									for (i = 0; i < SIZE; i = i + 1)
										begin
											// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:147:348
											ram[i] = INIT_VALUE;
										end
								end
							end
						end
						// Trace: ../../rtl/libs/VX_sp_ram.sv:149:21
						always @(posedge clk)
							// Trace: ../../rtl/libs/VX_sp_ram.sv:150:25
							begin : sv2v_autoblock_14
								// Trace: ../../rtl/libs/VX_sp_ram.sv:150:30
								integer i;
								// Trace: ../../rtl/libs/VX_sp_ram.sv:150:30
								for (i = 0; i < BYTEENW; i = i + 1)
									begin
										// Trace: ../../rtl/libs/VX_sp_ram.sv:151:29
										if (wren[i])
											// Trace: ../../rtl/libs/VX_sp_ram.sv:152:33
											ram[addr][i * 8+:8] <= wdata[i * 8+:8];
									end
							end
						// Trace: ../../rtl/libs/VX_sp_ram.sv:155:21
						assign rdata = ram[addr];
					end
					else begin : genblk1
						// Trace: ../../rtl/libs/VX_sp_ram.sv:157:21
						reg [DATAW - 1:0] ram [SIZE - 1:0];
						if (INIT_ENABLE) begin : genblk1
							if (INIT_FILE != "") begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:159:136
								initial begin
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:159:144
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : genblk1
								// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:159:238
								initial begin : sv2v_autoblock_15
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:159:298
									integer i;
									// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:159:298
									for (i = 0; i < SIZE; i = i + 1)
										begin
											// Trace: macro expansion of RAM_INITIALIZATION at ../../rtl/libs/VX_sp_ram.sv:159:348
											ram[i] = INIT_VALUE;
										end
								end
							end
						end
						// Trace: ../../rtl/libs/VX_sp_ram.sv:161:21
						always @(posedge clk)
							// Trace: ../../rtl/libs/VX_sp_ram.sv:162:25
							if (wren)
								// Trace: ../../rtl/libs/VX_sp_ram.sv:163:29
								ram[addr] <= wdata;
						// Trace: ../../rtl/libs/VX_sp_ram.sv:165:21
						assign rdata = ram[addr];
					end
				end
			end
		end
	endgenerate
endmodule
module VX_stream_arbiter (
	clk,
	reset,
	valid_in,
	data_in,
	ready_in,
	valid_out,
	data_out,
	ready_out
);
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:4:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:5:15
	parameter LANES = 1;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:6:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:7:15
	parameter TYPE = "P";
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:8:15
	parameter LOCK_ENABLE = 1;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:9:15
	parameter BUFFERED = 0;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:11:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:12:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:14:5
	input wire [(NUM_REQS * LANES) - 1:0] valid_in;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:15:5
	input wire [((NUM_REQS * LANES) * DATAW) - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:16:5
	output wire [(NUM_REQS * LANES) - 1:0] ready_in;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:18:5
	output wire [LANES - 1:0] valid_out;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:19:5
	output wire [(LANES * DATAW) - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:20:5
	input wire [LANES - 1:0] ready_out;
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:22:5
	localparam LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: ../../rtl/libs/VX_stream_arbiter.sv:24:5
	generate
		if (NUM_REQS > 1) begin : genblk1
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:25:9
			wire sel_valid;
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:26:9
			wire sel_ready;
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:27:9
			wire [LOG_NUM_REQS - 1:0] sel_index;
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:28:9
			wire [NUM_REQS - 1:0] sel_onehot;
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:30:9
			wire [NUM_REQS - 1:0] valid_in_any;
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:31:9
			wire [LANES - 1:0] ready_in_sel;
			if (LANES > 1) begin : genblk1
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_stream_arbiter.sv:35:17
					assign valid_in_any[i] = |valid_in[i * LANES+:LANES];
				end
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:37:13
				assign sel_ready = |ready_in_sel;
			end
			else begin : genblk1
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_stream_arbiter.sv:40:17
					assign valid_in_any[i] = valid_in[i * LANES+:LANES];
				end
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:42:13
				assign sel_ready = ready_in_sel;
			end
			if (TYPE == "P") begin : genblk2
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:46:13
				VX_fixed_arbiter #(
					.NUM_REQS(NUM_REQS),
					.LOCK_ENABLE(LOCK_ENABLE)
				) sel_arb(
					.clk(clk),
					.reset(reset),
					.requests(valid_in_any),
					.enable(sel_ready),
					.grant_valid(sel_valid),
					.grant_index(sel_index),
					.grant_onehot(sel_onehot)
				);
			end
			else if (TYPE == "R") begin : genblk2
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:59:13
				VX_rr_arbiter #(
					.NUM_REQS(NUM_REQS),
					.LOCK_ENABLE(LOCK_ENABLE)
				) sel_arb(
					.clk(clk),
					.reset(reset),
					.requests(valid_in_any),
					.enable(sel_ready),
					.grant_valid(sel_valid),
					.grant_index(sel_index),
					.grant_onehot(sel_onehot)
				);
			end
			else if (TYPE == "F") begin : genblk2
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:72:13
				VX_fair_arbiter #(
					.NUM_REQS(NUM_REQS),
					.LOCK_ENABLE(LOCK_ENABLE)
				) sel_arb(
					.clk(clk),
					.reset(reset),
					.requests(valid_in_any),
					.enable(sel_ready),
					.grant_valid(sel_valid),
					.grant_index(sel_index),
					.grant_onehot(sel_onehot)
				);
			end
			else if (TYPE == "M") begin : genblk2
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:85:13
				VX_matrix_arbiter #(
					.NUM_REQS(NUM_REQS),
					.LOCK_ENABLE(LOCK_ENABLE)
				) sel_arb(
					.clk(clk),
					.reset(reset),
					.requests(valid_in_any),
					.enable(sel_ready),
					.grant_valid(sel_valid),
					.grant_index(sel_index),
					.grant_onehot(sel_onehot)
				);
			end
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:101:9
			wire [LANES - 1:0] valid_in_sel;
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:102:9
			wire [(LANES * DATAW) - 1:0] data_in_sel;
			if (LANES > 1) begin : genblk3
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:105:13
				wire [(NUM_REQS * (LANES * (1 + DATAW))) - 1:0] valid_data_in;
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_stream_arbiter.sv:107:17
					assign valid_data_in[i * (LANES * (1 + DATAW))+:LANES * (1 + DATAW)] = {valid_in[i * LANES+:LANES], data_in[DATAW * (i * LANES)+:DATAW * LANES]};
				end
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:109:13
				assign {valid_in_sel, data_in_sel} = valid_data_in[sel_index * (LANES * (1 + DATAW))+:LANES * (1 + DATAW)];
			end
			else begin : genblk3
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:112:13
				assign data_in_sel = data_in[DATAW * (sel_index * LANES)+:DATAW * LANES];
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:113:13
				assign valid_in_sel = sel_valid;
			end
			genvar i;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk4
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:117:13
				assign ready_in[i * LANES+:LANES] = ready_in_sel & {LANES {sel_onehot[i]}};
			end
			for (i = 0; i < LANES; i = i + 1) begin : genblk5
				// Trace: ../../rtl/libs/VX_stream_arbiter.sv:121:13
				VX_skid_buffer #(
					.DATAW(DATAW),
					.PASSTHRU(0 == BUFFERED),
					.OUT_REG(2 == BUFFERED)
				) out_buffer(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in_sel[i]),
					.data_in(data_in_sel[i * DATAW+:DATAW]),
					.ready_in(ready_in_sel[i]),
					.valid_out(valid_out[i]),
					.data_out(data_out[i * DATAW+:DATAW]),
					.ready_out(ready_out[i])
				);
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:142:9
			assign valid_out = valid_in;
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:143:9
			assign data_out = data_in;
			// Trace: ../../rtl/libs/VX_stream_arbiter.sv:144:9
			assign ready_in = ready_out;
		end
	endgenerate
endmodule
module VX_stream_demux (
	clk,
	reset,
	sel_in,
	valid_in,
	data_in,
	ready_in,
	valid_out,
	data_out,
	ready_out
);
	// Trace: ../../rtl/libs/VX_stream_demux.sv:4:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:5:15
	parameter LANES = 1;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:6:15
	parameter DATAW = 1;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:7:15
	parameter BUFFERED = 0;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:8:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: ../../rtl/libs/VX_stream_demux.sv:10:5
	input wire clk;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:11:5
	input wire reset;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:13:5
	input wire [(LANES * LOG_NUM_REQS) - 1:0] sel_in;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:15:5
	input wire [LANES - 1:0] valid_in;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:16:5
	input wire [(LANES * DATAW) - 1:0] data_in;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:17:5
	output wire [LANES - 1:0] ready_in;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:19:5
	output wire [(NUM_REQS * LANES) - 1:0] valid_out;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:20:5
	output wire [((NUM_REQS * LANES) * DATAW) - 1:0] data_out;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:21:5
	input wire [(NUM_REQS * LANES) - 1:0] ready_out;
	// Trace: ../../rtl/libs/VX_stream_demux.sv:24:5
	generate
		if (NUM_REQS > 1) begin : genblk1
			genvar j;
			for (j = 0; j < LANES; j = j + 1) begin : genblk1
				// Trace: ../../rtl/libs/VX_stream_demux.sv:28:13
				reg [NUM_REQS - 1:0] valid_in_sel;
				// Trace: ../../rtl/libs/VX_stream_demux.sv:29:13
				wire [NUM_REQS - 1:0] ready_in_sel;
				// Trace: ../../rtl/libs/VX_stream_demux.sv:31:13
				always @(*) begin
					// Trace: ../../rtl/libs/VX_stream_demux.sv:32:17
					valid_in_sel = 1'sb0;
					// Trace: ../../rtl/libs/VX_stream_demux.sv:33:17
					valid_in_sel[sel_in[j * LOG_NUM_REQS+:LOG_NUM_REQS]] = valid_in[j];
				end
				// Trace: ../../rtl/libs/VX_stream_demux.sv:36:13
				assign ready_in[j] = ready_in_sel[sel_in[j * LOG_NUM_REQS+:LOG_NUM_REQS]];
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/libs/VX_stream_demux.sv:39:17
					VX_skid_buffer #(
						.DATAW(DATAW),
						.PASSTHRU(0 == BUFFERED),
						.OUT_REG(2 == BUFFERED)
					) out_buffer(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_in_sel[i]),
						.data_in(data_in[j * DATAW+:DATAW]),
						.ready_in(ready_in_sel[i]),
						.valid_out(valid_out[(i * LANES) + j]),
						.data_out(data_out[((i * LANES) + j) * DATAW+:DATAW]),
						.ready_out(ready_out[(i * LANES) + j])
					);
				end
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/libs/VX_stream_demux.sv:62:9
			assign valid_out = valid_in;
			// Trace: ../../rtl/libs/VX_stream_demux.sv:63:9
			assign data_out = data_in;
			// Trace: ../../rtl/libs/VX_stream_demux.sv:64:9
			assign ready_in = ready_out;
		end
	endgenerate
endmodule
// removed interface: VX_alu_req_if
// removed interface: VX_branch_ctl_if
// removed interface: VX_cmt_to_csr_if
// removed interface: VX_commit_if
// removed interface: VX_csr_req_if
// removed interface: VX_dcache_req_if
// removed interface: VX_dcache_rsp_if
// removed interface: VX_decode_if
// removed interface: VX_fetch_to_csr_if
// removed interface: VX_fpu_req_if
// removed interface: VX_fpu_to_csr_if
// removed interface: VX_gpr_req_if
// removed interface: VX_gpr_rsp_if
// removed interface: VX_gpu_req_if
// removed interface: VX_ibuffer_if
// removed interface: VX_icache_req_if
// removed interface: VX_icache_rsp_if
// removed interface: VX_ifetch_req_if
// removed interface: VX_ifetch_rsp_if
// removed interface: VX_join_if
// removed interface: VX_lsu_req_if
// removed interface: VX_mem_req_if
// removed interface: VX_mem_rsp_if
// removed interface: VX_perf_cache_if
// removed interface: VX_perf_memsys_if
// removed interface: VX_perf_pipeline_if
// removed interface: VX_perf_tex_if
// removed interface: VX_tex_csr_if
// removed interface: VX_tex_req_if
// removed interface: VX_tex_rsp_if
// removed interface: VX_warp_ctl_if
// removed interface: VX_writeback_if
// removed interface: VX_wstall_if
module VX_bank (
	clk,
	reset,
	core_req_valid,
	core_req_pmask,
	core_req_wsel,
	core_req_byteen,
	core_req_data,
	core_req_tid,
	core_req_tag,
	core_req_rw,
	core_req_addr,
	core_req_ready,
	core_rsp_valid,
	core_rsp_pmask,
	core_rsp_tid,
	core_rsp_data,
	core_rsp_tag,
	core_rsp_ready,
	mem_req_valid,
	mem_req_rw,
	mem_req_pmask,
	mem_req_byteen,
	mem_req_wsel,
	mem_req_addr,
	mem_req_id,
	mem_req_data,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_id,
	mem_rsp_data,
	mem_rsp_ready,
	flush_enable,
	flush_addr
);
	// Trace: ../../rtl/cache/VX_bank.sv:4:15
	parameter CACHE_ID = 0;
	// Trace: ../../rtl/cache/VX_bank.sv:5:15
	parameter BANK_ID = 0;
	// Trace: ../../rtl/cache/VX_bank.sv:8:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:11:15
	parameter CACHE_SIZE = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:13:15
	parameter CACHE_LINE_SIZE = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:15:15
	parameter NUM_BANKS = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:17:15
	parameter NUM_PORTS = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:19:15
	parameter WORD_SIZE = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:22:15
	parameter CREQ_SIZE = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:24:15
	parameter CRSQ_SIZE = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:26:15
	parameter MSHR_SIZE = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:28:15
	parameter MREQ_SIZE = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:31:15
	parameter WRITE_ENABLE = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:34:15
	parameter CORE_TAG_WIDTH = 1;
	// Trace: ../../rtl/cache/VX_bank.sv:37:15
	parameter BANK_ADDR_OFFSET = 0;
	// Trace: ../../rtl/cache/VX_bank.sv:39:15
	parameter MSHR_ADDR_WIDTH = $clog2(MSHR_SIZE);
	// Trace: ../../rtl/cache/VX_bank.sv:40:15
	parameter WORD_SELECT_BITS = ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1);
	// Trace: ../../rtl/cache/VX_bank.sv:44:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_bank.sv:45:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_bank.sv:54:5
	input wire core_req_valid;
	// Trace: ../../rtl/cache/VX_bank.sv:55:5
	input wire [NUM_PORTS - 1:0] core_req_pmask;
	// Trace: ../../rtl/cache/VX_bank.sv:56:5
	input wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] core_req_wsel;
	// Trace: ../../rtl/cache/VX_bank.sv:57:5
	input wire [(NUM_PORTS * WORD_SIZE) - 1:0] core_req_byteen;
	// Trace: ../../rtl/cache/VX_bank.sv:58:5
	input wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] core_req_data;
	// Trace: ../../rtl/cache/VX_bank.sv:59:5
	input wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] core_req_tid;
	// Trace: ../../rtl/cache/VX_bank.sv:60:5
	input wire [(NUM_PORTS * CORE_TAG_WIDTH) - 1:0] core_req_tag;
	// Trace: ../../rtl/cache/VX_bank.sv:61:5
	input wire core_req_rw;
	// Trace: ../../rtl/cache/VX_bank.sv:62:5
	input wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] core_req_addr;
	// Trace: ../../rtl/cache/VX_bank.sv:63:5
	output wire core_req_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:66:5
	output wire core_rsp_valid;
	// Trace: ../../rtl/cache/VX_bank.sv:67:5
	output wire [NUM_PORTS - 1:0] core_rsp_pmask;
	// Trace: ../../rtl/cache/VX_bank.sv:68:5
	output wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] core_rsp_tid;
	// Trace: ../../rtl/cache/VX_bank.sv:69:5
	output wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] core_rsp_data;
	// Trace: ../../rtl/cache/VX_bank.sv:70:5
	output wire [(NUM_PORTS * CORE_TAG_WIDTH) - 1:0] core_rsp_tag;
	// Trace: ../../rtl/cache/VX_bank.sv:71:5
	input wire core_rsp_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:74:5
	output wire mem_req_valid;
	// Trace: ../../rtl/cache/VX_bank.sv:75:5
	output wire mem_req_rw;
	// Trace: ../../rtl/cache/VX_bank.sv:76:5
	output wire [NUM_PORTS - 1:0] mem_req_pmask;
	// Trace: ../../rtl/cache/VX_bank.sv:77:5
	output wire [(NUM_PORTS * WORD_SIZE) - 1:0] mem_req_byteen;
	// Trace: ../../rtl/cache/VX_bank.sv:78:5
	output wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] mem_req_wsel;
	// Trace: ../../rtl/cache/VX_bank.sv:79:5
	output wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mem_req_addr;
	// Trace: ../../rtl/cache/VX_bank.sv:80:5
	output wire [MSHR_ADDR_WIDTH - 1:0] mem_req_id;
	// Trace: ../../rtl/cache/VX_bank.sv:81:5
	output wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] mem_req_data;
	// Trace: ../../rtl/cache/VX_bank.sv:82:5
	input wire mem_req_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:85:5
	input wire mem_rsp_valid;
	// Trace: ../../rtl/cache/VX_bank.sv:86:5
	input wire [MSHR_ADDR_WIDTH - 1:0] mem_rsp_id;
	// Trace: ../../rtl/cache/VX_bank.sv:87:5
	input wire [(8 * CACHE_LINE_SIZE) - 1:0] mem_rsp_data;
	// Trace: ../../rtl/cache/VX_bank.sv:88:5
	output wire mem_rsp_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:91:5
	input wire flush_enable;
	// Trace: ../../rtl/cache/VX_bank.sv:92:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0] flush_addr;
	// Trace: ../../rtl/cache/VX_bank.sv:96:5
	wire [43:0] req_id_sel;
	wire [43:0] req_id_st0;
	wire [43:0] req_id_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:99:5
	wire [NUM_PORTS - 1:0] creq_pmask;
	// Trace: ../../rtl/cache/VX_bank.sv:100:5
	wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] creq_wsel;
	// Trace: ../../rtl/cache/VX_bank.sv:101:5
	wire [(NUM_PORTS * WORD_SIZE) - 1:0] creq_byteen;
	// Trace: ../../rtl/cache/VX_bank.sv:102:5
	wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] creq_data;
	// Trace: ../../rtl/cache/VX_bank.sv:103:5
	wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] creq_tid;
	// Trace: ../../rtl/cache/VX_bank.sv:104:5
	wire [(NUM_PORTS * CORE_TAG_WIDTH) - 1:0] creq_tag;
	// Trace: ../../rtl/cache/VX_bank.sv:105:5
	wire creq_rw;
	// Trace: ../../rtl/cache/VX_bank.sv:106:5
	wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] creq_addr;
	// Trace: ../../rtl/cache/VX_bank.sv:108:5
	wire creq_valid;
	wire creq_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:110:5
	VX_elastic_buffer #(
		.DATAW((1 + ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) + (NUM_PORTS * (((((1 + WORD_SELECT_BITS) + WORD_SIZE) + (8 * WORD_SIZE)) + (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) + CORE_TAG_WIDTH))),
		.SIZE(CREQ_SIZE)
	) core_req_queue(
		.clk(clk),
		.reset(reset),
		.ready_in(core_req_ready),
		.valid_in(core_req_valid),
		.data_in({core_req_rw, core_req_addr, core_req_pmask, core_req_wsel, core_req_byteen, core_req_data, core_req_tid, core_req_tag}),
		.data_out({creq_rw, creq_addr, creq_pmask, creq_wsel, creq_byteen, creq_data, creq_tid, creq_tag}),
		.ready_out(creq_ready),
		.valid_out(creq_valid)
	);
	// Trace: ../../rtl/cache/VX_bank.sv:124:5
	wire mreq_alm_full;
	// Trace: ../../rtl/cache/VX_bank.sv:125:5
	wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mem_rsp_addr;
	// Trace: ../../rtl/cache/VX_bank.sv:126:5
	wire crsq_valid;
	wire crsq_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:127:5
	wire crsq_stall;
	// Trace: ../../rtl/cache/VX_bank.sv:129:5
	wire mshr_valid;
	// Trace: ../../rtl/cache/VX_bank.sv:130:5
	wire mshr_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:131:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_alloc_id;
	// Trace: ../../rtl/cache/VX_bank.sv:132:5
	wire mshr_alm_full;
	// Trace: ../../rtl/cache/VX_bank.sv:133:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_dequeue_id;
	// Trace: ../../rtl/cache/VX_bank.sv:134:5
	wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mshr_addr;
	// Trace: ../../rtl/cache/VX_bank.sv:135:5
	wire [(NUM_PORTS * CORE_TAG_WIDTH) - 1:0] mshr_tag;
	// Trace: ../../rtl/cache/VX_bank.sv:136:5
	wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] mshr_wsel;
	// Trace: ../../rtl/cache/VX_bank.sv:137:5
	wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] mshr_tid;
	// Trace: ../../rtl/cache/VX_bank.sv:138:5
	wire [NUM_PORTS - 1:0] mshr_pmask;
	// Trace: ../../rtl/cache/VX_bank.sv:140:5
	wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_st0;
	wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:141:5
	wire is_read_st0;
	wire is_read_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:142:5
	wire is_write_st0;
	wire is_write_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:143:5
	wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] wsel_st0;
	wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] wsel_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:144:5
	wire [(NUM_PORTS * WORD_SIZE) - 1:0] byteen_st0;
	wire [(NUM_PORTS * WORD_SIZE) - 1:0] byteen_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:145:5
	wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] req_tid_st0;
	wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] req_tid_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:146:5
	wire [NUM_PORTS - 1:0] pmask_st0;
	wire [NUM_PORTS - 1:0] pmask_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:147:5
	wire [(NUM_PORTS * CORE_TAG_WIDTH) - 1:0] tag_st0;
	wire [(NUM_PORTS * CORE_TAG_WIDTH) - 1:0] tag_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:148:5
	wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] rdata_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:149:5
	wire [(8 * CACHE_LINE_SIZE) - 1:0] wdata_st0;
	wire [(8 * CACHE_LINE_SIZE) - 1:0] wdata_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:150:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_id_st0;
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_id_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:151:5
	wire valid_st0;
	wire valid_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:152:5
	wire is_fill_st0;
	wire is_fill_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:153:5
	wire is_mshr_st0;
	wire is_mshr_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:154:5
	wire miss_st0;
	wire miss_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:155:5
	wire is_flush_st0;
	// Trace: ../../rtl/cache/VX_bank.sv:156:5
	wire mshr_pending_st0;
	wire mshr_pending_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:159:5
	wire rdw_fill_hazard = valid_st0 && is_fill_st0;
	// Trace: ../../rtl/cache/VX_bank.sv:160:5
	wire rdw_write_hazard = (valid_st0 && is_write_st0) && ~creq_rw;
	// Trace: ../../rtl/cache/VX_bank.sv:163:5
	wire mshr_grant = !flush_enable;
	// Trace: ../../rtl/cache/VX_bank.sv:164:5
	wire mshr_enable = mshr_grant && mshr_valid;
	// Trace: ../../rtl/cache/VX_bank.sv:166:5
	wire mrsq_grant = !flush_enable && !mshr_enable;
	// Trace: ../../rtl/cache/VX_bank.sv:167:5
	wire mrsq_enable = mrsq_grant && mem_rsp_valid;
	// Trace: ../../rtl/cache/VX_bank.sv:168:5
	wire creq_grant = (!flush_enable && !mshr_enable) && !mrsq_enable;
	// Trace: ../../rtl/cache/VX_bank.sv:170:5
	wire creq_enable = creq_grant && creq_valid;
	// Trace: ../../rtl/cache/VX_bank.sv:172:5
	assign mshr_ready = (mshr_grant && !rdw_fill_hazard) && !crsq_stall;
	// Trace: ../../rtl/cache/VX_bank.sv:177:5
	assign mem_rsp_ready = mrsq_grant && !crsq_stall;
	// Trace: ../../rtl/cache/VX_bank.sv:180:5
	assign creq_ready = (((creq_grant && !rdw_write_hazard) && !mreq_alm_full) && !mshr_alm_full) && !crsq_stall;
	// Trace: ../../rtl/cache/VX_bank.sv:186:5
	wire flush_fire = flush_enable;
	// Trace: ../../rtl/cache/VX_bank.sv:187:5
	wire mshr_fire = mshr_valid && mshr_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:188:5
	wire mem_rsp_fire = mem_rsp_valid && mem_rsp_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:189:5
	wire creq_fire = creq_valid && creq_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:191:5
	assign req_id_sel = (mshr_enable ? mshr_tag[0 + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? CORE_TAG_WIDTH - 1 : ((CORE_TAG_WIDTH - 1) + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)) - 1)-:((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)] : creq_tag[0 + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? CORE_TAG_WIDTH - 1 : ((CORE_TAG_WIDTH - 1) + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)) - 1)-:((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)]);
	// Trace: ../../rtl/cache/VX_bank.sv:193:5
	wire [(8 * CACHE_LINE_SIZE) - 1:0] wdata_sel;
	// Trace: ../../rtl/cache/VX_bank.sv:194:5
	assign wdata_sel[(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] = (mem_rsp_valid || !WRITE_ENABLE ? mem_rsp_data[(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] : creq_data);
	// Trace: ../../rtl/cache/VX_bank.sv:195:5
	genvar i;
	generate
		for (i = NUM_PORTS * (8 * WORD_SIZE); i < (8 * CACHE_LINE_SIZE); i = i + 1) begin : genblk1
			// Trace: ../../rtl/cache/VX_bank.sv:196:9
			assign wdata_sel[i] = mem_rsp_data[i];
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_bank.sv:199:5
	function automatic [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] sv2v_cast_FD4D3;
		input reg [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] inp;
		sv2v_cast_FD4D3 = inp;
	endfunction
	VX_pipe_register #(
		.DATAW((((6 + ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) + (8 * CACHE_LINE_SIZE)) + (NUM_PORTS * ((((WORD_SELECT_BITS + WORD_SIZE) + (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) + 1) + CORE_TAG_WIDTH))) + MSHR_ADDR_WIDTH),
		.RESETW(1)
	) pipe_reg0(
		.clk(clk),
		.reset(reset),
		.enable(!crsq_stall),
		.data_in({((flush_fire || mshr_fire) || mem_rsp_fire) || creq_fire, flush_enable, mshr_enable, mrsq_enable, creq_enable && ~creq_rw, creq_enable && creq_rw, (flush_enable ? sv2v_cast_FD4D3(flush_addr) : (mshr_valid ? mshr_addr : (mem_rsp_valid ? mem_rsp_addr : creq_addr))), wdata_sel, (mshr_valid ? mshr_wsel : creq_wsel), creq_byteen, (mshr_valid ? mshr_tid : creq_tid), (mshr_valid ? mshr_pmask : creq_pmask), (mshr_valid ? mshr_tag : creq_tag), (mshr_valid ? mshr_dequeue_id : mem_rsp_id)}),
		.data_out({valid_st0, is_flush_st0, is_mshr_st0, is_fill_st0, is_read_st0, is_write_st0, addr_st0, wdata_st0, wsel_st0, byteen_st0, req_tid_st0, pmask_st0, tag_st0, mshr_id_st0})
	);
	// Trace: ../../rtl/cache/VX_bank.sv:225:5
	assign req_id_st0 = tag_st0[0 + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? CORE_TAG_WIDTH - 1 : ((CORE_TAG_WIDTH - 1) + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)) - 1)-:((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)];
	// Trace: ../../rtl/cache/VX_bank.sv:227:5
	wire do_fill_st0 = valid_st0 && is_fill_st0;
	// Trace: ../../rtl/cache/VX_bank.sv:228:5
	wire do_flush_st0 = valid_st0 && is_flush_st0;
	// Trace: ../../rtl/cache/VX_bank.sv:229:5
	wire do_lookup_st0 = valid_st0 && ~(is_fill_st0 || is_flush_st0);
	// Trace: ../../rtl/cache/VX_bank.sv:231:5
	wire tag_match_st0;
	// Trace: ../../rtl/cache/VX_bank.sv:233:5
	VX_tag_access #(
		.BANK_ID(BANK_ID),
		.CACHE_ID(CACHE_ID),
		.CACHE_SIZE(CACHE_SIZE),
		.CACHE_LINE_SIZE(CACHE_LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.WORD_SIZE(WORD_SIZE),
		.BANK_ADDR_OFFSET(BANK_ADDR_OFFSET)
	) tag_access(
		.clk(clk),
		.reset(reset),
		.req_id(req_id_st0),
		.stall(crsq_stall),
		.lookup(do_lookup_st0),
		.addr(addr_st0),
		.fill(do_fill_st0),
		.flush(do_flush_st0),
		.tag_match(tag_match_st0)
	);
	// Trace: ../../rtl/cache/VX_bank.sv:258:5
	assign miss_st0 = (is_read_st0 || is_write_st0) && ~tag_match_st0;
	// Trace: ../../rtl/cache/VX_bank.sv:260:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_id_a_st0 = (is_read_st0 || is_write_st0 ? mshr_alloc_id : mshr_id_st0);
	// Trace: ../../rtl/cache/VX_bank.sv:262:5
	VX_pipe_register #(
		.DATAW(((((6 + ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) + (8 * CACHE_LINE_SIZE)) + (NUM_PORTS * ((((WORD_SELECT_BITS + WORD_SIZE) + (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) + 1) + CORE_TAG_WIDTH))) + MSHR_ADDR_WIDTH) + 1),
		.RESETW(1)
	) pipe_reg1(
		.clk(clk),
		.reset(reset),
		.enable(!crsq_stall),
		.data_in({valid_st0, is_mshr_st0, is_fill_st0, is_read_st0, is_write_st0, miss_st0, addr_st0, wdata_st0, wsel_st0, byteen_st0, req_tid_st0, pmask_st0, tag_st0, mshr_id_a_st0, mshr_pending_st0}),
		.data_out({valid_st1, is_mshr_st1, is_fill_st1, is_read_st1, is_write_st1, miss_st1, addr_st1, wdata_st1, wsel_st1, byteen_st1, req_tid_st1, pmask_st1, tag_st1, mshr_id_st1, mshr_pending_st1})
	);
	// Trace: ../../rtl/cache/VX_bank.sv:273:5
	assign req_id_st1 = tag_st1[0 + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? CORE_TAG_WIDTH - 1 : ((CORE_TAG_WIDTH - 1) + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)) - 1)-:((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)];
	// Trace: ../../rtl/cache/VX_bank.sv:275:5
	wire do_read_st0 = valid_st0 && is_read_st0;
	// Trace: ../../rtl/cache/VX_bank.sv:276:5
	wire do_read_st1 = valid_st1 && is_read_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:277:5
	wire do_fill_st1 = valid_st1 && is_fill_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:278:5
	wire do_write_st1 = valid_st1 && is_write_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:279:5
	wire do_mshr_st1 = valid_st1 && is_mshr_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:281:5
	wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] creq_data_st1 = wdata_st1[0+:NUM_PORTS * (8 * WORD_SIZE)];
	// Trace: ../../rtl/cache/VX_bank.sv:284:5
	VX_data_access #(
		.BANK_ID(BANK_ID),
		.CACHE_ID(CACHE_ID),
		.CACHE_SIZE(CACHE_SIZE),
		.CACHE_LINE_SIZE(CACHE_LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_PORTS(NUM_PORTS),
		.WORD_SIZE(WORD_SIZE),
		.WRITE_ENABLE(WRITE_ENABLE)
	) data_access(
		.clk(clk),
		.reset(reset),
		.req_id(req_id_st1),
		.stall(crsq_stall),
		.read(do_read_st1 || do_mshr_st1),
		.fill(do_fill_st1),
		.write(do_write_st1 && !miss_st1),
		.addr(addr_st1),
		.wsel(wsel_st1),
		.pmask(pmask_st1),
		.byteen(byteen_st1),
		.fill_data(wdata_st1),
		.write_data(creq_data_st1),
		.read_data(rdata_st1)
	);
	// Trace: ../../rtl/cache/VX_bank.sv:313:5
	wire mshr_allocate = do_read_st0 && !crsq_stall;
	// Trace: ../../rtl/cache/VX_bank.sv:314:5
	wire mshr_replay = do_fill_st0 && !crsq_stall;
	// Trace: ../../rtl/cache/VX_bank.sv:315:5
	wire mshr_lookup = mshr_allocate;
	// Trace: ../../rtl/cache/VX_bank.sv:316:5
	wire mshr_release = (do_read_st1 && !miss_st1) && !crsq_stall;
	// Trace: ../../rtl/cache/VX_bank.sv:318:5
	VX_pending_size #(.SIZE(MSHR_SIZE)) mshr_pending_size(
		.clk(clk),
		.reset(reset),
		.incr(creq_fire && ~creq_rw),
		.decr(mshr_fire || mshr_release),
		.full(mshr_alm_full)
	);
	// Trace: ../../rtl/cache/VX_bank.sv:330:5
	VX_miss_resrv #(
		.BANK_ID(BANK_ID),
		.CACHE_ID(CACHE_ID),
		.CACHE_LINE_SIZE(CACHE_LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_PORTS(NUM_PORTS),
		.WORD_SIZE(WORD_SIZE),
		.NUM_REQS(NUM_REQS),
		.MSHR_SIZE(MSHR_SIZE),
		.CORE_TAG_WIDTH(CORE_TAG_WIDTH)
	) miss_resrv(
		.clk(clk),
		.reset(reset),
		.deq_req_id(req_id_sel),
		.lkp_req_id(req_id_st0),
		.rel_req_id(req_id_st1),
		.allocate_valid(mshr_allocate),
		.allocate_addr(addr_st0),
		.allocate_data({wsel_st0, tag_st0, req_tid_st0, pmask_st0}),
		.allocate_id(mshr_alloc_id),
		.lookup_valid(mshr_lookup),
		.lookup_replay(mshr_replay),
		.lookup_id(mshr_alloc_id),
		.lookup_addr(addr_st0),
		.lookup_match(mshr_pending_st0),
		.fill_valid(mem_rsp_fire),
		.fill_id(mem_rsp_id),
		.fill_addr(mem_rsp_addr),
		.dequeue_valid(mshr_valid),
		.dequeue_id(mshr_dequeue_id),
		.dequeue_addr(mshr_addr),
		.dequeue_data({mshr_wsel, mshr_tag, mshr_tid, mshr_pmask}),
		.dequeue_ready(mshr_ready),
		.release_valid(mshr_release),
		.release_id(mshr_id_st1)
	);
	// Trace: ../../rtl/cache/VX_bank.sv:381:5
	wire [NUM_PORTS - 1:0] crsq_pmask;
	// Trace: ../../rtl/cache/VX_bank.sv:382:5
	wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] crsq_data;
	// Trace: ../../rtl/cache/VX_bank.sv:383:5
	wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] crsq_tid;
	// Trace: ../../rtl/cache/VX_bank.sv:384:5
	wire [(NUM_PORTS * CORE_TAG_WIDTH) - 1:0] crsq_tag;
	// Trace: ../../rtl/cache/VX_bank.sv:386:5
	assign crsq_valid = (do_read_st1 && !miss_st1) || do_mshr_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:389:5
	assign crsq_stall = crsq_valid && !crsq_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:391:5
	assign crsq_pmask = pmask_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:392:5
	assign crsq_tid = req_tid_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:393:5
	assign crsq_data = rdata_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:394:5
	assign crsq_tag = tag_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:396:5
	VX_elastic_buffer #(
		.DATAW(NUM_PORTS * (((CORE_TAG_WIDTH + 1) + (8 * WORD_SIZE)) + (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1))),
		.SIZE(CRSQ_SIZE),
		.OUT_REG(1)
	) core_rsp_req(
		.clk(clk),
		.reset(reset),
		.valid_in(crsq_valid),
		.data_in({crsq_tag, crsq_pmask, crsq_data, crsq_tid}),
		.ready_in(crsq_ready),
		.valid_out(core_rsp_valid),
		.data_out({core_rsp_tag, core_rsp_pmask, core_rsp_data, core_rsp_tid}),
		.ready_out(core_rsp_ready)
	);
	// Trace: ../../rtl/cache/VX_bank.sv:413:5
	wire mreq_push;
	wire mreq_pop;
	wire mreq_empty;
	// Trace: ../../rtl/cache/VX_bank.sv:414:5
	wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] mreq_data;
	// Trace: ../../rtl/cache/VX_bank.sv:415:5
	wire [(NUM_PORTS * WORD_SIZE) - 1:0] mreq_byteen;
	// Trace: ../../rtl/cache/VX_bank.sv:416:5
	wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] mreq_wsel;
	// Trace: ../../rtl/cache/VX_bank.sv:417:5
	wire [NUM_PORTS - 1:0] mreq_pmask;
	// Trace: ../../rtl/cache/VX_bank.sv:418:5
	wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mreq_addr;
	// Trace: ../../rtl/cache/VX_bank.sv:419:5
	wire [MSHR_ADDR_WIDTH - 1:0] mreq_id;
	// Trace: ../../rtl/cache/VX_bank.sv:420:5
	wire mreq_rw;
	// Trace: ../../rtl/cache/VX_bank.sv:422:5
	assign mreq_push = ((do_read_st1 && miss_st1) && !mshr_pending_st1) || do_write_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:425:5
	assign mreq_pop = mem_req_valid && mem_req_ready;
	// Trace: ../../rtl/cache/VX_bank.sv:427:5
	assign mreq_rw = WRITE_ENABLE && is_write_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:428:5
	assign mreq_addr = addr_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:429:5
	assign mreq_id = mshr_id_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:430:5
	assign mreq_pmask = pmask_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:431:5
	assign mreq_wsel = wsel_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:432:5
	assign mreq_byteen = byteen_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:433:5
	assign mreq_data = creq_data_st1;
	// Trace: ../../rtl/cache/VX_bank.sv:435:5
	VX_fifo_queue #(
		.DATAW(((1 + ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) + MSHR_ADDR_WIDTH) + (NUM_PORTS * (((1 + WORD_SIZE) + WORD_SELECT_BITS) + (8 * WORD_SIZE)))),
		.SIZE(MREQ_SIZE),
		.ALM_FULL(MREQ_SIZE - 2),
		.OUT_REG(1 == NUM_BANKS)
	) mem_req_queue(
		.clk(clk),
		.reset(reset),
		.push(mreq_push),
		.pop(mreq_pop),
		.data_in({mreq_rw, mreq_addr, mreq_id, mreq_pmask, mreq_byteen, mreq_wsel, mreq_data}),
		.data_out({mem_req_rw, mem_req_addr, mem_req_id, mem_req_pmask, mem_req_byteen, mem_req_wsel, mem_req_data}),
		.empty(mreq_empty),
		.alm_full(mreq_alm_full)
	);
	// Trace: ../../rtl/cache/VX_bank.sv:454:5
	assign mem_req_valid = !mreq_empty;
endmodule
module VX_cache (
	clk,
	reset,
	core_req_valid,
	core_req_rw,
	core_req_addr,
	core_req_byteen,
	core_req_data,
	core_req_tag,
	core_req_ready,
	core_rsp_valid,
	core_rsp_tmask,
	core_rsp_data,
	core_rsp_tag,
	core_rsp_ready,
	mem_req_valid,
	mem_req_rw,
	mem_req_byteen,
	mem_req_addr,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready
);
	// Trace: ../../rtl/cache/VX_cache.sv:4:15
	parameter CACHE_ID = 0;
	// Trace: ../../rtl/cache/VX_cache.sv:7:15
	parameter NUM_REQS = 4;
	// Trace: ../../rtl/cache/VX_cache.sv:10:15
	parameter CACHE_SIZE = 16384;
	// Trace: ../../rtl/cache/VX_cache.sv:12:15
	parameter CACHE_LINE_SIZE = 64;
	// Trace: ../../rtl/cache/VX_cache.sv:14:15
	parameter NUM_BANKS = NUM_REQS;
	// Trace: ../../rtl/cache/VX_cache.sv:16:15
	parameter NUM_PORTS = 1;
	// Trace: ../../rtl/cache/VX_cache.sv:18:15
	parameter WORD_SIZE = 4;
	// Trace: ../../rtl/cache/VX_cache.sv:21:15
	parameter CREQ_SIZE = 0;
	// Trace: ../../rtl/cache/VX_cache.sv:23:15
	parameter CRSQ_SIZE = 2;
	// Trace: ../../rtl/cache/VX_cache.sv:25:15
	parameter MSHR_SIZE = 8;
	// Trace: ../../rtl/cache/VX_cache.sv:27:15
	parameter MRSQ_SIZE = 0;
	// Trace: ../../rtl/cache/VX_cache.sv:29:15
	parameter MREQ_SIZE = 4;
	// Trace: ../../rtl/cache/VX_cache.sv:32:15
	parameter WRITE_ENABLE = 1;
	// Trace: ../../rtl/cache/VX_cache.sv:35:15
	parameter CORE_TAG_WIDTH = $clog2(MSHR_SIZE);
	// Trace: ../../rtl/cache/VX_cache.sv:38:15
	parameter CORE_TAG_ID_BITS = CORE_TAG_WIDTH;
	// Trace: ../../rtl/cache/VX_cache.sv:41:15
	parameter MEM_TAG_WIDTH = 32 - $clog2(CACHE_LINE_SIZE);
	// Trace: ../../rtl/cache/VX_cache.sv:44:15
	parameter BANK_ADDR_OFFSET = 0;
	// Trace: ../../rtl/cache/VX_cache.sv:47:15
	parameter NC_ENABLE = 0;
	// Trace: ../../rtl/cache/VX_cache.sv:49:15
	parameter WORD_SELECT_BITS = ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1);
	// Trace: ../../rtl/cache/VX_cache.sv:58:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_cache.sv:59:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_cache.sv:62:5
	input wire [NUM_REQS - 1:0] core_req_valid;
	// Trace: ../../rtl/cache/VX_cache.sv:63:5
	input wire [NUM_REQS - 1:0] core_req_rw;
	// Trace: ../../rtl/cache/VX_cache.sv:64:5
	input wire [(NUM_REQS * (32 - $clog2(WORD_SIZE))) - 1:0] core_req_addr;
	// Trace: ../../rtl/cache/VX_cache.sv:65:5
	input wire [(NUM_REQS * WORD_SIZE) - 1:0] core_req_byteen;
	// Trace: ../../rtl/cache/VX_cache.sv:66:5
	input wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_req_data;
	// Trace: ../../rtl/cache/VX_cache.sv:67:5
	input wire [(NUM_REQS * CORE_TAG_WIDTH) - 1:0] core_req_tag;
	// Trace: ../../rtl/cache/VX_cache.sv:68:5
	output wire [NUM_REQS - 1:0] core_req_ready;
	// Trace: ../../rtl/cache/VX_cache.sv:71:5
	output wire [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_valid;
	// Trace: ../../rtl/cache/VX_cache.sv:72:5
	output wire [NUM_REQS - 1:0] core_rsp_tmask;
	// Trace: ../../rtl/cache/VX_cache.sv:73:5
	output wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_rsp_data;
	// Trace: ../../rtl/cache/VX_cache.sv:74:5
	output wire [((CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) * CORE_TAG_WIDTH) - 1:0] core_rsp_tag;
	// Trace: ../../rtl/cache/VX_cache.sv:75:5
	input wire [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_ready;
	// Trace: ../../rtl/cache/VX_cache.sv:78:5
	output wire mem_req_valid;
	// Trace: ../../rtl/cache/VX_cache.sv:79:5
	output wire mem_req_rw;
	// Trace: ../../rtl/cache/VX_cache.sv:80:5
	output wire [CACHE_LINE_SIZE - 1:0] mem_req_byteen;
	// Trace: ../../rtl/cache/VX_cache.sv:81:5
	output wire [(32 - $clog2(CACHE_LINE_SIZE)) - 1:0] mem_req_addr;
	// Trace: ../../rtl/cache/VX_cache.sv:82:5
	output wire [(8 * CACHE_LINE_SIZE) - 1:0] mem_req_data;
	// Trace: ../../rtl/cache/VX_cache.sv:83:5
	output wire [MEM_TAG_WIDTH - 1:0] mem_req_tag;
	// Trace: ../../rtl/cache/VX_cache.sv:84:5
	input wire mem_req_ready;
	// Trace: ../../rtl/cache/VX_cache.sv:87:5
	input wire mem_rsp_valid;
	// Trace: ../../rtl/cache/VX_cache.sv:88:5
	input wire [(8 * CACHE_LINE_SIZE) - 1:0] mem_rsp_data;
	// Trace: ../../rtl/cache/VX_cache.sv:89:5
	input wire [MEM_TAG_WIDTH - 1:0] mem_rsp_tag;
	// Trace: ../../rtl/cache/VX_cache.sv:90:5
	output wire mem_rsp_ready;
	// Trace: ../../rtl/cache/VX_cache.sv:96:5
	localparam MSHR_ADDR_WIDTH = $clog2(MSHR_SIZE);
	// Trace: ../../rtl/cache/VX_cache.sv:97:5
	localparam MEM_TAG_IN_WIDTH = $clog2(NUM_BANKS) + MSHR_ADDR_WIDTH;
	// Trace: ../../rtl/cache/VX_cache.sv:98:5
	localparam CORE_TAG_X_WIDTH = CORE_TAG_WIDTH - NC_ENABLE;
	// Trace: ../../rtl/cache/VX_cache.sv:99:5
	localparam CORE_TAG_ID_X_BITS = (CORE_TAG_ID_BITS != 0 ? CORE_TAG_ID_BITS - NC_ENABLE : CORE_TAG_ID_BITS);
	// Trace: ../../rtl/cache/VX_cache.sv:109:5
	wire mem_req_valid_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:110:5
	wire mem_req_rw_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:111:5
	wire [CACHE_LINE_SIZE - 1:0] mem_req_byteen_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:112:5
	wire [(32 - $clog2(CACHE_LINE_SIZE)) - 1:0] mem_req_addr_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:113:5
	wire [(8 * CACHE_LINE_SIZE) - 1:0] mem_req_data_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:114:5
	wire [MEM_TAG_WIDTH - 1:0] mem_req_tag_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:115:5
	wire mem_req_ready_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:117:5
	VX_skid_buffer #(
		.DATAW((((1 + CACHE_LINE_SIZE) + (32 - $clog2(CACHE_LINE_SIZE))) + (8 * CACHE_LINE_SIZE)) + MEM_TAG_WIDTH),
		.PASSTHRU(1 == NUM_BANKS)
	) mem_req_sbuf(
		.clk(clk),
		.reset(reset),
		.valid_in(mem_req_valid_sb),
		.ready_in(mem_req_ready_sb),
		.data_in({mem_req_rw_sb, mem_req_byteen_sb, mem_req_addr_sb, mem_req_data_sb, mem_req_tag_sb}),
		.data_out({mem_req_rw, mem_req_byteen, mem_req_addr, mem_req_data, mem_req_tag}),
		.valid_out(mem_req_valid),
		.ready_out(mem_req_ready)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:133:5
	wire [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_valid_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:134:5
	wire [NUM_REQS - 1:0] core_rsp_tmask_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:135:5
	wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_rsp_data_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:136:5
	wire [((CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) * CORE_TAG_WIDTH) - 1:0] core_rsp_tag_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:137:5
	wire [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_ready_sb;
	// Trace: ../../rtl/cache/VX_cache.sv:139:5
	generate
		if (CORE_TAG_ID_BITS != 0) begin : genblk1
			// Trace: ../../rtl/cache/VX_cache.sv:140:9
			VX_skid_buffer #(
				.DATAW((NUM_REQS + (NUM_REQS * (8 * WORD_SIZE))) + CORE_TAG_WIDTH),
				.PASSTHRU(1 == NUM_BANKS)
			) core_rsp_sbuf(
				.clk(clk),
				.reset(reset),
				.valid_in(core_rsp_valid_sb),
				.ready_in(core_rsp_ready_sb),
				.data_in({core_rsp_tmask_sb, core_rsp_data_sb, core_rsp_tag_sb}),
				.data_out({core_rsp_tmask, core_rsp_data, core_rsp_tag}),
				.valid_out(core_rsp_valid),
				.ready_out(core_rsp_ready)
			);
		end
		else begin : genblk1
			genvar i;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_cache.sv:155:13
				VX_skid_buffer #(
					.DATAW((1 + (8 * WORD_SIZE)) + CORE_TAG_WIDTH),
					.PASSTHRU(1 == NUM_BANKS)
				) core_rsp_sbuf(
					.clk(clk),
					.reset(reset),
					.valid_in(core_rsp_valid_sb[i]),
					.ready_in(core_rsp_ready_sb[i]),
					.data_in({core_rsp_tmask_sb[i], core_rsp_data_sb[i * (8 * WORD_SIZE)+:8 * WORD_SIZE], core_rsp_tag_sb[i * CORE_TAG_WIDTH+:CORE_TAG_WIDTH]}),
					.data_out({core_rsp_tmask[i], core_rsp_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE], core_rsp_tag[i * CORE_TAG_WIDTH+:CORE_TAG_WIDTH]}),
					.valid_out(core_rsp_valid[i]),
					.ready_out(core_rsp_ready[i])
				);
			end
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_cache.sv:174:5
	wire [(NUM_PORTS * WORD_SIZE) - 1:0] mem_req_byteen_p;
	// Trace: ../../rtl/cache/VX_cache.sv:175:5
	wire [NUM_PORTS - 1:0] mem_req_pmask_p;
	// Trace: ../../rtl/cache/VX_cache.sv:176:5
	wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] mem_req_wsel_p;
	// Trace: ../../rtl/cache/VX_cache.sv:177:5
	wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] mem_req_data_p;
	// Trace: ../../rtl/cache/VX_cache.sv:178:5
	wire mem_req_rw_p;
	// Trace: ../../rtl/cache/VX_cache.sv:180:5
	generate
		if (WRITE_ENABLE) begin : genblk2
			if ((CACHE_LINE_SIZE / WORD_SIZE) > 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_cache.sv:182:13
				reg [CACHE_LINE_SIZE - 1:0] mem_req_byteen_r;
				// Trace: ../../rtl/cache/VX_cache.sv:183:13
				reg [(8 * CACHE_LINE_SIZE) - 1:0] mem_req_data_r;
				// Trace: ../../rtl/cache/VX_cache.sv:185:13
				always @(*) begin
					// Trace: ../../rtl/cache/VX_cache.sv:186:17
					mem_req_byteen_r = 0;
					// Trace: ../../rtl/cache/VX_cache.sv:187:17
					mem_req_data_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_cache.sv:188:17
					begin : sv2v_autoblock_1
						// Trace: ../../rtl/cache/VX_cache.sv:188:22
						integer i;
						// Trace: ../../rtl/cache/VX_cache.sv:188:22
						for (i = 0; i < NUM_PORTS; i = i + 1)
							begin
								// Trace: ../../rtl/cache/VX_cache.sv:189:21
								if ((1 == NUM_PORTS) || mem_req_pmask_p[i]) begin
									// Trace: ../../rtl/cache/VX_cache.sv:190:25
									mem_req_byteen_r[mem_req_wsel_p[i * WORD_SELECT_BITS+:WORD_SELECT_BITS] * WORD_SIZE+:WORD_SIZE] = mem_req_byteen_p[i * WORD_SIZE+:WORD_SIZE];
									// Trace: ../../rtl/cache/VX_cache.sv:191:25
									mem_req_data_r[mem_req_wsel_p[i * WORD_SELECT_BITS+:WORD_SELECT_BITS] * (8 * WORD_SIZE)+:8 * WORD_SIZE] = mem_req_data_p[i * (8 * WORD_SIZE)+:8 * WORD_SIZE];
								end
							end
					end
				end
				// Trace: ../../rtl/cache/VX_cache.sv:196:13
				assign mem_req_rw_sb = mem_req_rw_p;
				// Trace: ../../rtl/cache/VX_cache.sv:197:13
				assign mem_req_byteen_sb = mem_req_byteen_r;
				// Trace: ../../rtl/cache/VX_cache.sv:198:13
				assign mem_req_data_sb = mem_req_data_r;
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_cache.sv:202:13
				assign mem_req_rw_sb = mem_req_rw_p;
				// Trace: ../../rtl/cache/VX_cache.sv:203:13
				assign mem_req_byteen_sb = mem_req_byteen_p;
				// Trace: ../../rtl/cache/VX_cache.sv:204:13
				assign mem_req_data_sb = mem_req_data_p;
			end
		end
		else begin : genblk2
			// Trace: ../../rtl/cache/VX_cache.sv:213:9
			assign mem_req_rw_sb = 0;
			// Trace: ../../rtl/cache/VX_cache.sv:214:9
			assign mem_req_byteen_sb = 1'sbx;
			// Trace: ../../rtl/cache/VX_cache.sv:215:9
			assign mem_req_data_sb = 1'sbx;
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_cache.sv:221:5
	wire [NUM_REQS - 1:0] core_req_valid_c;
	// Trace: ../../rtl/cache/VX_cache.sv:222:5
	wire [NUM_REQS - 1:0] core_req_rw_c;
	// Trace: ../../rtl/cache/VX_cache.sv:223:5
	wire [(NUM_REQS * (32 - $clog2(WORD_SIZE))) - 1:0] core_req_addr_c;
	// Trace: ../../rtl/cache/VX_cache.sv:224:5
	wire [(NUM_REQS * WORD_SIZE) - 1:0] core_req_byteen_c;
	// Trace: ../../rtl/cache/VX_cache.sv:225:5
	wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_req_data_c;
	// Trace: ../../rtl/cache/VX_cache.sv:226:5
	wire [(NUM_REQS * CORE_TAG_X_WIDTH) - 1:0] core_req_tag_c;
	// Trace: ../../rtl/cache/VX_cache.sv:227:5
	wire [NUM_REQS - 1:0] core_req_ready_c;
	// Trace: ../../rtl/cache/VX_cache.sv:230:5
	wire [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_valid_c;
	// Trace: ../../rtl/cache/VX_cache.sv:231:5
	wire [NUM_REQS - 1:0] core_rsp_tmask_c;
	// Trace: ../../rtl/cache/VX_cache.sv:232:5
	wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_rsp_data_c;
	// Trace: ../../rtl/cache/VX_cache.sv:233:5
	wire [((CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) * CORE_TAG_X_WIDTH) - 1:0] core_rsp_tag_c;
	// Trace: ../../rtl/cache/VX_cache.sv:234:5
	wire [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_ready_c;
	// Trace: ../../rtl/cache/VX_cache.sv:237:5
	wire mem_req_valid_c;
	// Trace: ../../rtl/cache/VX_cache.sv:238:5
	wire mem_req_rw_c;
	// Trace: ../../rtl/cache/VX_cache.sv:239:5
	wire [(32 - $clog2(CACHE_LINE_SIZE)) - 1:0] mem_req_addr_c;
	// Trace: ../../rtl/cache/VX_cache.sv:240:5
	wire [NUM_PORTS - 1:0] mem_req_pmask_c;
	// Trace: ../../rtl/cache/VX_cache.sv:241:5
	wire [(NUM_PORTS * WORD_SIZE) - 1:0] mem_req_byteen_c;
	// Trace: ../../rtl/cache/VX_cache.sv:242:5
	wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] mem_req_wsel_c;
	// Trace: ../../rtl/cache/VX_cache.sv:243:5
	wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] mem_req_data_c;
	// Trace: ../../rtl/cache/VX_cache.sv:244:5
	wire [MEM_TAG_IN_WIDTH - 1:0] mem_req_tag_c;
	// Trace: ../../rtl/cache/VX_cache.sv:245:5
	wire mem_req_ready_c;
	// Trace: ../../rtl/cache/VX_cache.sv:248:5
	wire mem_rsp_valid_c;
	// Trace: ../../rtl/cache/VX_cache.sv:249:5
	wire [(8 * CACHE_LINE_SIZE) - 1:0] mem_rsp_data_c;
	// Trace: ../../rtl/cache/VX_cache.sv:250:5
	wire [MEM_TAG_IN_WIDTH - 1:0] mem_rsp_tag_c;
	// Trace: ../../rtl/cache/VX_cache.sv:251:5
	wire mem_rsp_ready_c;
	// Trace: ../../rtl/cache/VX_cache.sv:253:5
	generate
		if (NC_ENABLE) begin : genblk3
			// Trace: ../../rtl/cache/VX_cache.sv:254:9
			VX_nc_bypass #(
				.NUM_PORTS(NUM_PORTS),
				.NUM_REQS(NUM_REQS),
				.NUM_RSP_TAGS((CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS)),
				.NC_TAG_BIT(0),
				.CORE_ADDR_WIDTH(32 - $clog2(WORD_SIZE)),
				.CORE_DATA_SIZE(WORD_SIZE),
				.CORE_TAG_IN_WIDTH(CORE_TAG_WIDTH),
				.MEM_ADDR_WIDTH(32 - $clog2(CACHE_LINE_SIZE)),
				.MEM_DATA_SIZE(CACHE_LINE_SIZE),
				.MEM_TAG_IN_WIDTH(MEM_TAG_IN_WIDTH),
				.MEM_TAG_OUT_WIDTH(MEM_TAG_WIDTH)
			) nc_bypass(
				.clk(clk),
				.reset(reset),
				.core_req_valid_in(core_req_valid),
				.core_req_rw_in(core_req_rw),
				.core_req_byteen_in(core_req_byteen),
				.core_req_addr_in(core_req_addr),
				.core_req_data_in(core_req_data),
				.core_req_tag_in(core_req_tag),
				.core_req_ready_in(core_req_ready),
				.core_req_valid_out(core_req_valid_c),
				.core_req_rw_out(core_req_rw_c),
				.core_req_byteen_out(core_req_byteen_c),
				.core_req_addr_out(core_req_addr_c),
				.core_req_data_out(core_req_data_c),
				.core_req_tag_out(core_req_tag_c),
				.core_req_ready_out(core_req_ready_c),
				.core_rsp_valid_in(core_rsp_valid_c),
				.core_rsp_tmask_in(core_rsp_tmask_c),
				.core_rsp_data_in(core_rsp_data_c),
				.core_rsp_tag_in(core_rsp_tag_c),
				.core_rsp_ready_in(core_rsp_ready_c),
				.core_rsp_valid_out(core_rsp_valid_sb),
				.core_rsp_tmask_out(core_rsp_tmask_sb),
				.core_rsp_data_out(core_rsp_data_sb),
				.core_rsp_tag_out(core_rsp_tag_sb),
				.core_rsp_ready_out(core_rsp_ready_sb),
				.mem_req_valid_in(mem_req_valid_c),
				.mem_req_rw_in(mem_req_rw_c),
				.mem_req_addr_in(mem_req_addr_c),
				.mem_req_pmask_in(mem_req_pmask_c),
				.mem_req_byteen_in(mem_req_byteen_c),
				.mem_req_wsel_in(mem_req_wsel_c),
				.mem_req_data_in(mem_req_data_c),
				.mem_req_tag_in(mem_req_tag_c),
				.mem_req_ready_in(mem_req_ready_c),
				.mem_req_valid_out(mem_req_valid_sb),
				.mem_req_addr_out(mem_req_addr_sb),
				.mem_req_rw_out(mem_req_rw_p),
				.mem_req_pmask_out(mem_req_pmask_p),
				.mem_req_byteen_out(mem_req_byteen_p),
				.mem_req_wsel_out(mem_req_wsel_p),
				.mem_req_data_out(mem_req_data_p),
				.mem_req_tag_out(mem_req_tag_sb),
				.mem_req_ready_out(mem_req_ready_sb),
				.mem_rsp_valid_in(mem_rsp_valid),
				.mem_rsp_data_in(mem_rsp_data),
				.mem_rsp_tag_in(mem_rsp_tag),
				.mem_rsp_ready_in(mem_rsp_ready),
				.mem_rsp_valid_out(mem_rsp_valid_c),
				.mem_rsp_data_out(mem_rsp_data_c),
				.mem_rsp_tag_out(mem_rsp_tag_c),
				.mem_rsp_ready_out(mem_rsp_ready_c)
			);
		end
		else begin : genblk3
			// Trace: ../../rtl/cache/VX_cache.sv:339:9
			assign core_req_valid_c = core_req_valid;
			// Trace: ../../rtl/cache/VX_cache.sv:340:9
			assign core_req_rw_c = core_req_rw;
			// Trace: ../../rtl/cache/VX_cache.sv:341:9
			assign core_req_addr_c = core_req_addr;
			// Trace: ../../rtl/cache/VX_cache.sv:342:9
			assign core_req_byteen_c = core_req_byteen;
			// Trace: ../../rtl/cache/VX_cache.sv:343:9
			assign core_req_data_c = core_req_data;
			// Trace: ../../rtl/cache/VX_cache.sv:344:9
			assign core_req_tag_c = core_req_tag;
			// Trace: ../../rtl/cache/VX_cache.sv:345:9
			assign core_req_ready = core_req_ready_c;
			// Trace: ../../rtl/cache/VX_cache.sv:347:9
			assign core_rsp_valid_sb = core_rsp_valid_c;
			// Trace: ../../rtl/cache/VX_cache.sv:348:9
			assign core_rsp_tmask_sb = core_rsp_tmask_c;
			// Trace: ../../rtl/cache/VX_cache.sv:349:9
			assign core_rsp_data_sb = core_rsp_data_c;
			// Trace: ../../rtl/cache/VX_cache.sv:350:9
			assign core_rsp_tag_sb = core_rsp_tag_c;
			// Trace: ../../rtl/cache/VX_cache.sv:351:9
			assign core_rsp_ready_c = core_rsp_ready_sb;
			// Trace: ../../rtl/cache/VX_cache.sv:353:9
			assign mem_req_valid_sb = mem_req_valid_c;
			// Trace: ../../rtl/cache/VX_cache.sv:354:9
			assign mem_req_addr_sb = mem_req_addr_c;
			// Trace: ../../rtl/cache/VX_cache.sv:355:9
			assign mem_req_rw_p = mem_req_rw_c;
			// Trace: ../../rtl/cache/VX_cache.sv:356:9
			assign mem_req_pmask_p = mem_req_pmask_c;
			// Trace: ../../rtl/cache/VX_cache.sv:357:9
			assign mem_req_byteen_p = mem_req_byteen_c;
			// Trace: ../../rtl/cache/VX_cache.sv:358:9
			assign mem_req_wsel_p = mem_req_wsel_c;
			// Trace: ../../rtl/cache/VX_cache.sv:359:9
			assign mem_req_data_p = mem_req_data_c;
			// Trace: ../../rtl/cache/VX_cache.sv:360:9
			assign mem_req_tag_sb = mem_req_tag_c;
			// Trace: ../../rtl/cache/VX_cache.sv:361:9
			assign mem_req_ready_c = mem_req_ready_sb;
			// Trace: ../../rtl/cache/VX_cache.sv:363:9
			assign mem_rsp_valid_c = mem_rsp_valid;
			// Trace: ../../rtl/cache/VX_cache.sv:364:9
			assign mem_rsp_data_c = mem_rsp_data;
			// Trace: ../../rtl/cache/VX_cache.sv:365:9
			assign mem_rsp_tag_c = mem_rsp_tag;
			// Trace: ../../rtl/cache/VX_cache.sv:366:9
			assign mem_rsp_ready = mem_rsp_ready_c;
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_cache.sv:371:5
	wire [(8 * CACHE_LINE_SIZE) - 1:0] mem_rsp_data_qual;
	// Trace: ../../rtl/cache/VX_cache.sv:372:5
	wire [MEM_TAG_IN_WIDTH - 1:0] mem_rsp_tag_qual;
	// Trace: ../../rtl/cache/VX_cache.sv:374:5
	wire mrsq_out_valid;
	wire mrsq_out_ready;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/cache/VX_cache.sv:376:23
	wire mrsq_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/cache/VX_cache.sv:376:56
	VX_reset_relay __mrsq_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(mrsq_reset)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:378:5
	VX_elastic_buffer #(
		.DATAW(MEM_TAG_IN_WIDTH + (8 * CACHE_LINE_SIZE)),
		.SIZE(MRSQ_SIZE),
		.OUT_REG(MRSQ_SIZE > 2)
	) mem_rsp_queue(
		.clk(clk),
		.reset(mrsq_reset),
		.ready_in(mem_rsp_ready_c),
		.valid_in(mem_rsp_valid_c),
		.data_in({mem_rsp_tag_c, mem_rsp_data_c}),
		.data_out({mem_rsp_tag_qual, mem_rsp_data_qual}),
		.ready_out(mrsq_out_ready),
		.valid_out(mrsq_out_valid)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:397:5
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0] flush_addr;
	// Trace: ../../rtl/cache/VX_cache.sv:398:5
	wire flush_enable;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/cache/VX_cache.sv:400:24
	wire flush_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/cache/VX_cache.sv:400:57
	VX_reset_relay __flush_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(flush_reset)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:402:5
	VX_flush_ctrl #(
		.CACHE_SIZE(CACHE_SIZE),
		.CACHE_LINE_SIZE(CACHE_LINE_SIZE),
		.NUM_BANKS(NUM_BANKS)
	) flush_ctrl(
		.clk(clk),
		.reset(flush_reset),
		.addr_out(flush_addr),
		.valid_out(flush_enable)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:415:5
	wire [NUM_BANKS - 1:0] per_bank_core_req_valid;
	// Trace: ../../rtl/cache/VX_cache.sv:416:5
	wire [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_req_pmask;
	// Trace: ../../rtl/cache/VX_cache.sv:417:5
	wire [((NUM_BANKS * NUM_PORTS) * WORD_SELECT_BITS) - 1:0] per_bank_core_req_wsel;
	// Trace: ../../rtl/cache/VX_cache.sv:418:5
	wire [((NUM_BANKS * NUM_PORTS) * WORD_SIZE) - 1:0] per_bank_core_req_byteen;
	// Trace: ../../rtl/cache/VX_cache.sv:419:5
	wire [((NUM_BANKS * NUM_PORTS) * (8 * WORD_SIZE)) - 1:0] per_bank_core_req_data;
	// Trace: ../../rtl/cache/VX_cache.sv:420:5
	wire [((NUM_BANKS * NUM_PORTS) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] per_bank_core_req_tid;
	// Trace: ../../rtl/cache/VX_cache.sv:421:5
	wire [((NUM_BANKS * NUM_PORTS) * CORE_TAG_X_WIDTH) - 1:0] per_bank_core_req_tag;
	// Trace: ../../rtl/cache/VX_cache.sv:422:5
	wire [NUM_BANKS - 1:0] per_bank_core_req_rw;
	// Trace: ../../rtl/cache/VX_cache.sv:423:5
	wire [(NUM_BANKS * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] per_bank_core_req_addr;
	// Trace: ../../rtl/cache/VX_cache.sv:424:5
	wire [NUM_BANKS - 1:0] per_bank_core_req_ready;
	// Trace: ../../rtl/cache/VX_cache.sv:426:5
	wire [NUM_BANKS - 1:0] per_bank_core_rsp_valid;
	// Trace: ../../rtl/cache/VX_cache.sv:427:5
	wire [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_pmask;
	// Trace: ../../rtl/cache/VX_cache.sv:428:5
	wire [((NUM_BANKS * NUM_PORTS) * (8 * WORD_SIZE)) - 1:0] per_bank_core_rsp_data;
	// Trace: ../../rtl/cache/VX_cache.sv:429:5
	wire [((NUM_BANKS * NUM_PORTS) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] per_bank_core_rsp_tid;
	// Trace: ../../rtl/cache/VX_cache.sv:430:5
	wire [((NUM_BANKS * NUM_PORTS) * CORE_TAG_X_WIDTH) - 1:0] per_bank_core_rsp_tag;
	// Trace: ../../rtl/cache/VX_cache.sv:431:5
	wire [NUM_BANKS - 1:0] per_bank_core_rsp_ready;
	// Trace: ../../rtl/cache/VX_cache.sv:433:5
	wire [NUM_BANKS - 1:0] per_bank_mem_req_valid;
	// Trace: ../../rtl/cache/VX_cache.sv:434:5
	wire [NUM_BANKS - 1:0] per_bank_mem_req_rw;
	// Trace: ../../rtl/cache/VX_cache.sv:435:5
	wire [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_mem_req_pmask;
	// Trace: ../../rtl/cache/VX_cache.sv:436:5
	wire [((NUM_BANKS * NUM_PORTS) * WORD_SIZE) - 1:0] per_bank_mem_req_byteen;
	// Trace: ../../rtl/cache/VX_cache.sv:437:5
	wire [((NUM_BANKS * NUM_PORTS) * WORD_SELECT_BITS) - 1:0] per_bank_mem_req_wsel;
	// Trace: ../../rtl/cache/VX_cache.sv:438:5
	wire [(NUM_BANKS * (32 - $clog2(CACHE_LINE_SIZE))) - 1:0] per_bank_mem_req_addr;
	// Trace: ../../rtl/cache/VX_cache.sv:439:5
	wire [(NUM_BANKS * MSHR_ADDR_WIDTH) - 1:0] per_bank_mem_req_id;
	// Trace: ../../rtl/cache/VX_cache.sv:440:5
	wire [((NUM_BANKS * NUM_PORTS) * (8 * WORD_SIZE)) - 1:0] per_bank_mem_req_data;
	// Trace: ../../rtl/cache/VX_cache.sv:441:5
	wire [NUM_BANKS - 1:0] per_bank_mem_req_ready;
	// Trace: ../../rtl/cache/VX_cache.sv:443:5
	wire [NUM_BANKS - 1:0] per_bank_mem_rsp_ready;
	// Trace: ../../rtl/cache/VX_cache.sv:445:5
	generate
		if (NUM_BANKS == 1) begin : genblk4
			// Trace: ../../rtl/cache/VX_cache.sv:446:9
			assign mrsq_out_ready = per_bank_mem_rsp_ready;
		end
		else begin : genblk4
			// Trace: ../../rtl/cache/VX_cache.sv:448:9
			assign mrsq_out_ready = per_bank_mem_rsp_ready[mem_rsp_tag_qual[MSHR_ADDR_WIDTH+:$clog2(NUM_BANKS)]];
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_cache.sv:451:5
	VX_core_req_bank_sel #(
		.CACHE_ID(CACHE_ID),
		.CACHE_LINE_SIZE(CACHE_LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_PORTS(NUM_PORTS),
		.WORD_SIZE(WORD_SIZE),
		.NUM_REQS(NUM_REQS),
		.CORE_TAG_WIDTH(CORE_TAG_X_WIDTH),
		.BANK_ADDR_OFFSET(BANK_ADDR_OFFSET)
	) core_req_bank_sel(
		.clk(clk),
		.reset(reset),
		.core_req_valid(core_req_valid_c),
		.core_req_rw(core_req_rw_c),
		.core_req_addr(core_req_addr_c),
		.core_req_byteen(core_req_byteen_c),
		.core_req_data(core_req_data_c),
		.core_req_tag(core_req_tag_c),
		.core_req_ready(core_req_ready_c),
		.per_bank_core_req_valid(per_bank_core_req_valid),
		.per_bank_core_req_pmask(per_bank_core_req_pmask),
		.per_bank_core_req_rw(per_bank_core_req_rw),
		.per_bank_core_req_addr(per_bank_core_req_addr),
		.per_bank_core_req_wsel(per_bank_core_req_wsel),
		.per_bank_core_req_byteen(per_bank_core_req_byteen),
		.per_bank_core_req_data(per_bank_core_req_data),
		.per_bank_core_req_tag(per_bank_core_req_tag),
		.per_bank_core_req_tid(per_bank_core_req_tid),
		.per_bank_core_req_ready(per_bank_core_req_ready)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:487:5
	genvar i;
	function automatic signed [$clog2(NUM_BANKS) - 1:0] sv2v_cast_748B1_signed;
		input reg signed [$clog2(NUM_BANKS) - 1:0] inp;
		sv2v_cast_748B1_signed = inp;
	endfunction
	generate
		for (i = 0; i < NUM_BANKS; i = i + 1) begin : genblk5
			// Trace: ../../rtl/cache/VX_cache.sv:488:9
			wire curr_bank_core_req_valid;
			// Trace: ../../rtl/cache/VX_cache.sv:489:9
			wire [NUM_PORTS - 1:0] curr_bank_core_req_pmask;
			// Trace: ../../rtl/cache/VX_cache.sv:490:9
			wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] curr_bank_core_req_wsel;
			// Trace: ../../rtl/cache/VX_cache.sv:491:9
			wire [(NUM_PORTS * WORD_SIZE) - 1:0] curr_bank_core_req_byteen;
			// Trace: ../../rtl/cache/VX_cache.sv:492:9
			wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] curr_bank_core_req_data;
			// Trace: ../../rtl/cache/VX_cache.sv:493:9
			wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] curr_bank_core_req_tid;
			// Trace: ../../rtl/cache/VX_cache.sv:494:9
			wire [(NUM_PORTS * CORE_TAG_X_WIDTH) - 1:0] curr_bank_core_req_tag;
			// Trace: ../../rtl/cache/VX_cache.sv:495:9
			wire curr_bank_core_req_rw;
			// Trace: ../../rtl/cache/VX_cache.sv:496:9
			wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] curr_bank_core_req_addr;
			// Trace: ../../rtl/cache/VX_cache.sv:497:9
			wire curr_bank_core_req_ready;
			// Trace: ../../rtl/cache/VX_cache.sv:499:9
			wire curr_bank_core_rsp_valid;
			// Trace: ../../rtl/cache/VX_cache.sv:500:9
			wire [NUM_PORTS - 1:0] curr_bank_core_rsp_pmask;
			// Trace: ../../rtl/cache/VX_cache.sv:501:9
			wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] curr_bank_core_rsp_data;
			// Trace: ../../rtl/cache/VX_cache.sv:502:9
			wire [(NUM_PORTS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] curr_bank_core_rsp_tid;
			// Trace: ../../rtl/cache/VX_cache.sv:503:9
			wire [(NUM_PORTS * CORE_TAG_X_WIDTH) - 1:0] curr_bank_core_rsp_tag;
			// Trace: ../../rtl/cache/VX_cache.sv:504:9
			wire curr_bank_core_rsp_ready;
			// Trace: ../../rtl/cache/VX_cache.sv:506:9
			wire curr_bank_mem_req_valid;
			// Trace: ../../rtl/cache/VX_cache.sv:507:9
			wire curr_bank_mem_req_rw;
			// Trace: ../../rtl/cache/VX_cache.sv:508:9
			wire [NUM_PORTS - 1:0] curr_bank_mem_req_pmask;
			// Trace: ../../rtl/cache/VX_cache.sv:509:9
			wire [(NUM_PORTS * WORD_SIZE) - 1:0] curr_bank_mem_req_byteen;
			// Trace: ../../rtl/cache/VX_cache.sv:510:9
			wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] curr_bank_mem_req_wsel;
			// Trace: ../../rtl/cache/VX_cache.sv:511:9
			wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] curr_bank_mem_req_addr;
			// Trace: ../../rtl/cache/VX_cache.sv:512:9
			wire [MSHR_ADDR_WIDTH - 1:0] curr_bank_mem_req_id;
			// Trace: ../../rtl/cache/VX_cache.sv:513:9
			wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] curr_bank_mem_req_data;
			// Trace: ../../rtl/cache/VX_cache.sv:514:9
			wire curr_bank_mem_req_ready;
			// Trace: ../../rtl/cache/VX_cache.sv:516:9
			wire curr_bank_mem_rsp_valid;
			// Trace: ../../rtl/cache/VX_cache.sv:517:9
			wire [MSHR_ADDR_WIDTH - 1:0] curr_bank_mem_rsp_id;
			// Trace: ../../rtl/cache/VX_cache.sv:518:9
			wire [(8 * CACHE_LINE_SIZE) - 1:0] curr_bank_mem_rsp_data;
			// Trace: ../../rtl/cache/VX_cache.sv:519:9
			wire curr_bank_mem_rsp_ready;
			// Trace: ../../rtl/cache/VX_cache.sv:522:9
			assign curr_bank_core_req_valid = per_bank_core_req_valid[i];
			// Trace: ../../rtl/cache/VX_cache.sv:523:9
			assign curr_bank_core_req_pmask = per_bank_core_req_pmask[i * NUM_PORTS+:NUM_PORTS];
			// Trace: ../../rtl/cache/VX_cache.sv:524:9
			assign curr_bank_core_req_addr = per_bank_core_req_addr[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)];
			// Trace: ../../rtl/cache/VX_cache.sv:525:9
			assign curr_bank_core_req_rw = per_bank_core_req_rw[i];
			// Trace: ../../rtl/cache/VX_cache.sv:526:9
			assign curr_bank_core_req_wsel = per_bank_core_req_wsel[WORD_SELECT_BITS * (i * NUM_PORTS)+:WORD_SELECT_BITS * NUM_PORTS];
			// Trace: ../../rtl/cache/VX_cache.sv:527:9
			assign curr_bank_core_req_byteen = per_bank_core_req_byteen[WORD_SIZE * (i * NUM_PORTS)+:WORD_SIZE * NUM_PORTS];
			// Trace: ../../rtl/cache/VX_cache.sv:528:9
			assign curr_bank_core_req_data = per_bank_core_req_data[(8 * WORD_SIZE) * (i * NUM_PORTS)+:(8 * WORD_SIZE) * NUM_PORTS];
			// Trace: ../../rtl/cache/VX_cache.sv:529:9
			assign curr_bank_core_req_tag = per_bank_core_req_tag[CORE_TAG_X_WIDTH * (i * NUM_PORTS)+:CORE_TAG_X_WIDTH * NUM_PORTS];
			// Trace: ../../rtl/cache/VX_cache.sv:530:9
			assign curr_bank_core_req_tid = per_bank_core_req_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS];
			// Trace: ../../rtl/cache/VX_cache.sv:531:9
			assign per_bank_core_req_ready[i] = curr_bank_core_req_ready;
			// Trace: ../../rtl/cache/VX_cache.sv:534:9
			assign curr_bank_core_rsp_ready = per_bank_core_rsp_ready[i];
			// Trace: ../../rtl/cache/VX_cache.sv:535:9
			assign per_bank_core_rsp_valid[i] = curr_bank_core_rsp_valid;
			// Trace: ../../rtl/cache/VX_cache.sv:536:9
			assign per_bank_core_rsp_pmask[i * NUM_PORTS+:NUM_PORTS] = curr_bank_core_rsp_pmask;
			// Trace: ../../rtl/cache/VX_cache.sv:537:9
			assign per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS] = curr_bank_core_rsp_tid;
			// Trace: ../../rtl/cache/VX_cache.sv:538:9
			assign per_bank_core_rsp_tag[CORE_TAG_X_WIDTH * (i * NUM_PORTS)+:CORE_TAG_X_WIDTH * NUM_PORTS] = curr_bank_core_rsp_tag;
			// Trace: ../../rtl/cache/VX_cache.sv:539:9
			assign per_bank_core_rsp_data[(8 * WORD_SIZE) * (i * NUM_PORTS)+:(8 * WORD_SIZE) * NUM_PORTS] = curr_bank_core_rsp_data;
			// Trace: ../../rtl/cache/VX_cache.sv:542:9
			assign per_bank_mem_req_valid[i] = curr_bank_mem_req_valid;
			// Trace: ../../rtl/cache/VX_cache.sv:543:9
			assign per_bank_mem_req_rw[i] = curr_bank_mem_req_rw;
			// Trace: ../../rtl/cache/VX_cache.sv:544:9
			assign per_bank_mem_req_pmask[i * NUM_PORTS+:NUM_PORTS] = curr_bank_mem_req_pmask;
			// Trace: ../../rtl/cache/VX_cache.sv:545:9
			assign per_bank_mem_req_byteen[WORD_SIZE * (i * NUM_PORTS)+:WORD_SIZE * NUM_PORTS] = curr_bank_mem_req_byteen;
			// Trace: ../../rtl/cache/VX_cache.sv:546:9
			assign per_bank_mem_req_wsel[WORD_SELECT_BITS * (i * NUM_PORTS)+:WORD_SELECT_BITS * NUM_PORTS] = curr_bank_mem_req_wsel;
			if (NUM_BANKS == 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_cache.sv:548:13
				assign per_bank_mem_req_addr[i * (32 - $clog2(CACHE_LINE_SIZE))+:32 - $clog2(CACHE_LINE_SIZE)] = curr_bank_mem_req_addr;
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_cache.sv:550:13
				assign per_bank_mem_req_addr[i * (32 - $clog2(CACHE_LINE_SIZE))+:32 - $clog2(CACHE_LINE_SIZE)] = {curr_bank_mem_req_addr, sv2v_cast_748B1_signed(i)};
			end
			// Trace: ../../rtl/cache/VX_cache.sv:552:9
			assign per_bank_mem_req_id[i * MSHR_ADDR_WIDTH+:MSHR_ADDR_WIDTH] = curr_bank_mem_req_id;
			// Trace: ../../rtl/cache/VX_cache.sv:553:9
			assign per_bank_mem_req_data[(8 * WORD_SIZE) * (i * NUM_PORTS)+:(8 * WORD_SIZE) * NUM_PORTS] = curr_bank_mem_req_data;
			// Trace: ../../rtl/cache/VX_cache.sv:554:9
			assign curr_bank_mem_req_ready = per_bank_mem_req_ready[i];
			if (NUM_BANKS == 1) begin : genblk2
				// Trace: ../../rtl/cache/VX_cache.sv:558:13
				assign curr_bank_mem_rsp_valid = mrsq_out_valid;
			end
			else begin : genblk2
				// Trace: ../../rtl/cache/VX_cache.sv:560:13
				assign curr_bank_mem_rsp_valid = mrsq_out_valid && (mem_rsp_tag_qual[MSHR_ADDR_WIDTH+:$clog2(NUM_BANKS)] == i);
			end
			// Trace: ../../rtl/cache/VX_cache.sv:562:9
			assign curr_bank_mem_rsp_id = mem_rsp_tag_qual[MSHR_ADDR_WIDTH - 1:0];
			// Trace: ../../rtl/cache/VX_cache.sv:563:9
			assign curr_bank_mem_rsp_data = mem_rsp_data_qual;
			// Trace: ../../rtl/cache/VX_cache.sv:564:9
			assign per_bank_mem_rsp_ready[i] = curr_bank_mem_rsp_ready;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/cache/VX_cache.sv:566:27
			wire bank_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/cache/VX_cache.sv:566:60
			VX_reset_relay __bank_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(bank_reset)
			);
			// Trace: ../../rtl/cache/VX_cache.sv:568:9
			VX_bank #(
				.BANK_ID(i),
				.CACHE_ID(CACHE_ID),
				.CACHE_SIZE(CACHE_SIZE),
				.CACHE_LINE_SIZE(CACHE_LINE_SIZE),
				.NUM_BANKS(NUM_BANKS),
				.NUM_PORTS(NUM_PORTS),
				.WORD_SIZE(WORD_SIZE),
				.NUM_REQS(NUM_REQS),
				.CREQ_SIZE(CREQ_SIZE),
				.CRSQ_SIZE(CRSQ_SIZE),
				.MSHR_SIZE(MSHR_SIZE),
				.MREQ_SIZE(MREQ_SIZE),
				.WRITE_ENABLE(WRITE_ENABLE),
				.CORE_TAG_WIDTH(CORE_TAG_X_WIDTH),
				.BANK_ADDR_OFFSET(BANK_ADDR_OFFSET)
			) bank(
				.clk(clk),
				.reset(bank_reset),
				.core_req_valid(curr_bank_core_req_valid),
				.core_req_pmask(curr_bank_core_req_pmask),
				.core_req_rw(curr_bank_core_req_rw),
				.core_req_byteen(curr_bank_core_req_byteen),
				.core_req_addr(curr_bank_core_req_addr),
				.core_req_wsel(curr_bank_core_req_wsel),
				.core_req_data(curr_bank_core_req_data),
				.core_req_tag(curr_bank_core_req_tag),
				.core_req_tid(curr_bank_core_req_tid),
				.core_req_ready(curr_bank_core_req_ready),
				.core_rsp_valid(curr_bank_core_rsp_valid),
				.core_rsp_pmask(curr_bank_core_rsp_pmask),
				.core_rsp_tid(curr_bank_core_rsp_tid),
				.core_rsp_data(curr_bank_core_rsp_data),
				.core_rsp_tag(curr_bank_core_rsp_tag),
				.core_rsp_ready(curr_bank_core_rsp_ready),
				.mem_req_valid(curr_bank_mem_req_valid),
				.mem_req_rw(curr_bank_mem_req_rw),
				.mem_req_pmask(curr_bank_mem_req_pmask),
				.mem_req_byteen(curr_bank_mem_req_byteen),
				.mem_req_wsel(curr_bank_mem_req_wsel),
				.mem_req_addr(curr_bank_mem_req_addr),
				.mem_req_id(curr_bank_mem_req_id),
				.mem_req_data(curr_bank_mem_req_data),
				.mem_req_ready(curr_bank_mem_req_ready),
				.mem_rsp_valid(curr_bank_mem_rsp_valid),
				.mem_rsp_id(curr_bank_mem_rsp_id),
				.mem_rsp_data(curr_bank_mem_rsp_data),
				.mem_rsp_ready(curr_bank_mem_rsp_ready),
				.flush_enable(flush_enable),
				.flush_addr(flush_addr)
			);
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_cache.sv:639:5
	VX_core_rsp_merge #(
		.CACHE_ID(CACHE_ID),
		.NUM_BANKS(NUM_BANKS),
		.NUM_PORTS(NUM_PORTS),
		.WORD_SIZE(WORD_SIZE),
		.NUM_REQS(NUM_REQS),
		.CORE_TAG_WIDTH(CORE_TAG_X_WIDTH),
		.CORE_TAG_ID_BITS(CORE_TAG_ID_X_BITS)
	) core_rsp_merge(
		.clk(clk),
		.reset(reset),
		.per_bank_core_rsp_valid(per_bank_core_rsp_valid),
		.per_bank_core_rsp_pmask(per_bank_core_rsp_pmask),
		.per_bank_core_rsp_data(per_bank_core_rsp_data),
		.per_bank_core_rsp_tag(per_bank_core_rsp_tag),
		.per_bank_core_rsp_tid(per_bank_core_rsp_tid),
		.per_bank_core_rsp_ready(per_bank_core_rsp_ready),
		.core_rsp_valid(core_rsp_valid_c),
		.core_rsp_tmask(core_rsp_tmask_c),
		.core_rsp_tag(core_rsp_tag_c),
		.core_rsp_data(core_rsp_data_c),
		.core_rsp_ready(core_rsp_ready_c)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:663:5
	wire [(NUM_BANKS * ((((32 - $clog2(CACHE_LINE_SIZE)) + MSHR_ADDR_WIDTH) + 1) + (NUM_PORTS * (((1 + WORD_SIZE) + WORD_SELECT_BITS) + (8 * WORD_SIZE))))) - 1:0] data_in;
	// Trace: ../../rtl/cache/VX_cache.sv:664:5
	generate
		for (i = 0; i < NUM_BANKS; i = i + 1) begin : genblk6
			// Trace: ../../rtl/cache/VX_cache.sv:665:9
			assign data_in[i * ((((32 - $clog2(CACHE_LINE_SIZE)) + MSHR_ADDR_WIDTH) + 1) + (NUM_PORTS * (((1 + WORD_SIZE) + WORD_SELECT_BITS) + (8 * WORD_SIZE))))+:(((32 - $clog2(CACHE_LINE_SIZE)) + MSHR_ADDR_WIDTH) + 1) + (NUM_PORTS * (((1 + WORD_SIZE) + WORD_SELECT_BITS) + (8 * WORD_SIZE)))] = {per_bank_mem_req_addr[i * (32 - $clog2(CACHE_LINE_SIZE))+:32 - $clog2(CACHE_LINE_SIZE)], per_bank_mem_req_id[i * MSHR_ADDR_WIDTH+:MSHR_ADDR_WIDTH], per_bank_mem_req_rw[i], per_bank_mem_req_pmask[i * NUM_PORTS+:NUM_PORTS], per_bank_mem_req_byteen[WORD_SIZE * (i * NUM_PORTS)+:WORD_SIZE * NUM_PORTS], per_bank_mem_req_wsel[WORD_SELECT_BITS * (i * NUM_PORTS)+:WORD_SELECT_BITS * NUM_PORTS], per_bank_mem_req_data[(8 * WORD_SIZE) * (i * NUM_PORTS)+:(8 * WORD_SIZE) * NUM_PORTS]};
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_cache.sv:668:5
	wire [MSHR_ADDR_WIDTH - 1:0] mem_req_id;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/cache/VX_cache.sv:670:23
	wire mreq_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/cache/VX_cache.sv:670:56
	VX_reset_relay __mreq_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(mreq_reset)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:672:5
	VX_stream_arbiter #(
		.NUM_REQS(NUM_BANKS),
		.DATAW((((32 - $clog2(CACHE_LINE_SIZE)) + MSHR_ADDR_WIDTH) + 1) + (NUM_PORTS * (((1 + WORD_SIZE) + WORD_SELECT_BITS) + (8 * WORD_SIZE)))),
		.TYPE("R")
	) mem_req_arb(
		.clk(clk),
		.reset(mreq_reset),
		.valid_in(per_bank_mem_req_valid),
		.data_in(data_in),
		.ready_in(per_bank_mem_req_ready),
		.valid_out(mem_req_valid_c),
		.data_out({mem_req_addr_c, mem_req_id, mem_req_rw_c, mem_req_pmask_c, mem_req_byteen_c, mem_req_wsel_c, mem_req_data_c}),
		.ready_out(mem_req_ready_c)
	);
	// Trace: ../../rtl/cache/VX_cache.sv:687:5
	function automatic [MEM_TAG_IN_WIDTH - 1:0] sv2v_cast_4ECAF;
		input reg [MEM_TAG_IN_WIDTH - 1:0] inp;
		sv2v_cast_4ECAF = inp;
	endfunction
	generate
		if (NUM_BANKS == 1) begin : genblk7
			// Trace: ../../rtl/cache/VX_cache.sv:688:9
			assign mem_req_tag_c = sv2v_cast_4ECAF(mem_req_id);
		end
		else begin : genblk7
			// Trace: ../../rtl/cache/VX_cache.sv:690:9
			assign mem_req_tag_c = sv2v_cast_4ECAF({mem_req_addr_c[0+:$clog2(NUM_BANKS)], mem_req_id});
		end
	endgenerate
endmodule
module VX_core_req_bank_sel (
	clk,
	reset,
	core_req_valid,
	core_req_rw,
	core_req_addr,
	core_req_byteen,
	core_req_data,
	core_req_tag,
	core_req_ready,
	per_bank_core_req_valid,
	per_bank_core_req_pmask,
	per_bank_core_req_rw,
	per_bank_core_req_addr,
	per_bank_core_req_wsel,
	per_bank_core_req_byteen,
	per_bank_core_req_data,
	per_bank_core_req_tid,
	per_bank_core_req_tag,
	per_bank_core_req_ready
);
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:4:15
	parameter CACHE_ID = 0;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:7:15
	parameter CACHE_LINE_SIZE = 64;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:9:15
	parameter WORD_SIZE = 4;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:11:15
	parameter NUM_BANKS = 4;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:13:15
	parameter NUM_PORTS = 1;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:15:15
	parameter NUM_REQS = 4;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:17:15
	parameter CORE_TAG_WIDTH = 3;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:19:15
	parameter BANK_ADDR_OFFSET = 0;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:21:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:22:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:28:5
	input wire [NUM_REQS - 1:0] core_req_valid;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:29:5
	input wire [NUM_REQS - 1:0] core_req_rw;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:30:5
	input wire [(NUM_REQS * (32 - $clog2(WORD_SIZE))) - 1:0] core_req_addr;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:31:5
	input wire [(NUM_REQS * WORD_SIZE) - 1:0] core_req_byteen;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:32:5
	input wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_req_data;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:33:5
	input wire [(NUM_REQS * CORE_TAG_WIDTH) - 1:0] core_req_tag;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:34:5
	output wire [NUM_REQS - 1:0] core_req_ready;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:36:5
	output wire [NUM_BANKS - 1:0] per_bank_core_req_valid;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:37:5
	output wire [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_req_pmask;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:38:5
	output wire [NUM_BANKS - 1:0] per_bank_core_req_rw;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:39:5
	output wire [(NUM_BANKS * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] per_bank_core_req_addr;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:40:5
	output wire [((NUM_BANKS * NUM_PORTS) * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)) - 1:0] per_bank_core_req_wsel;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:41:5
	output wire [((NUM_BANKS * NUM_PORTS) * WORD_SIZE) - 1:0] per_bank_core_req_byteen;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:42:5
	output wire [((NUM_BANKS * NUM_PORTS) * (8 * WORD_SIZE)) - 1:0] per_bank_core_req_data;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:43:5
	output wire [((NUM_BANKS * NUM_PORTS) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] per_bank_core_req_tid;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:44:5
	output wire [((NUM_BANKS * NUM_PORTS) * CORE_TAG_WIDTH) - 1:0] per_bank_core_req_tag;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:45:5
	input wire [NUM_BANKS - 1:0] per_bank_core_req_ready;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:54:5
	wire [(NUM_REQS * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] core_req_line_addr;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:55:5
	wire [(NUM_REQS * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)) - 1:0] core_req_wsel;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:56:5
	wire [(NUM_REQS * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)) - 1:0] core_req_bid;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:58:5
	genvar i;
	generate
		for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
			if (BANK_ADDR_OFFSET == 0) begin : genblk1
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:60:13
				assign core_req_line_addr[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] = core_req_addr[(i * (32 - $clog2(WORD_SIZE))) + (((32 - $clog2(WORD_SIZE)) - 1) >= (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) ? (32 - $clog2(WORD_SIZE)) - 1 : (((32 - $clog2(WORD_SIZE)) - 1) + (((32 - $clog2(WORD_SIZE)) - 1) >= (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) ? (((32 - $clog2(WORD_SIZE)) - 1) - (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0)) + 1 : ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) - ((32 - $clog2(WORD_SIZE)) - 1)) + 1)) - 1)-:(((32 - $clog2(WORD_SIZE)) - 1) >= (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) ? (((32 - $clog2(WORD_SIZE)) - 1) - (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0)) + 1 : ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) - ((32 - $clog2(WORD_SIZE)) - 1)) + 1)];
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:62:13
				assign core_req_line_addr[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] = {core_req_addr[(i * (32 - $clog2(WORD_SIZE))) + (((32 - $clog2(WORD_SIZE)) - 1) >= (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) ? (32 - $clog2(WORD_SIZE)) - 1 : (((32 - $clog2(WORD_SIZE)) - 1) + (((32 - $clog2(WORD_SIZE)) - 1) >= (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) ? (((32 - $clog2(WORD_SIZE)) - 1) - (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0)) + 1 : ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) - ((32 - $clog2(WORD_SIZE)) - 1)) + 1)) - 1)-:(((32 - $clog2(WORD_SIZE)) - 1) >= (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) ? (((32 - $clog2(WORD_SIZE)) - 1) - (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0)) + 1 : ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) - ((32 - $clog2(WORD_SIZE)) - 1)) + 1)], core_req_addr[(i * (32 - $clog2(WORD_SIZE))) + (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1) >= ((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) ? (((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1 : (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1) + (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1) >= ((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) ? (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1) - ((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0)) + 1 : (((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) - ((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1)) + 1)) - 1)-:(((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1) >= ((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) ? (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1) - ((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0)) + 1 : (((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) - ((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - 1)) + 1)]};
			end
			// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:64:9
			assign core_req_wsel[i * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)+:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)] = core_req_addr[(i * (32 - $clog2(WORD_SIZE))) + (($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1) - 1)-:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)];
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:67:5
	generate
		for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk2
			if (NUM_BANKS > 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:69:13
				assign core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] = core_req_addr[(i * (32 - $clog2(WORD_SIZE))) + ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1) >= (((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) ? ((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1 : ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1) + ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1) >= (((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) ? ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1) - (((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET)) + 1 : ((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1)) + 1)) - 1)-:((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1) >= (((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) ? ((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1) - (((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET)) + 1 : ((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) - (((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) - 1)) + 1)];
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:71:13
				assign core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] = 0;
			end
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:75:5
	reg [NUM_BANKS - 1:0] per_bank_core_req_valid_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:76:5
	reg [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_req_pmask_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:77:5
	reg [((NUM_BANKS * NUM_PORTS) * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)) - 1:0] per_bank_core_req_wsel_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:78:5
	reg [((NUM_BANKS * NUM_PORTS) * WORD_SIZE) - 1:0] per_bank_core_req_byteen_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:79:5
	reg [((NUM_BANKS * NUM_PORTS) * (8 * WORD_SIZE)) - 1:0] per_bank_core_req_data_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:80:5
	reg [((NUM_BANKS * NUM_PORTS) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] per_bank_core_req_tid_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:81:5
	reg [((NUM_BANKS * NUM_PORTS) * CORE_TAG_WIDTH) - 1:0] per_bank_core_req_tag_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:82:5
	reg [NUM_BANKS - 1:0] per_bank_core_req_rw_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:83:5
	reg [(NUM_BANKS * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] per_bank_core_req_addr_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:84:5
	reg [NUM_REQS - 1:0] core_req_ready_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:86:5
	function automatic signed [(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) - 1:0] sv2v_cast_CC627_signed;
		input reg signed [(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) - 1:0] inp;
		sv2v_cast_CC627_signed = inp;
	endfunction
	generate
		if (NUM_REQS > 1) begin : genblk3
			if (NUM_PORTS > 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:90:13
				reg [(NUM_BANKS * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] per_bank_line_addr_r;
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:91:13
				reg [NUM_BANKS - 1:0] per_bank_rw_r;
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:92:13
				wire [NUM_REQS - 1:0] core_req_line_match;
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:94:13
				always @(*) begin
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:95:17
					per_bank_line_addr_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:96:17
					begin : sv2v_autoblock_1
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:96:22
						integer i;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:96:22
						for (i = NUM_REQS - 1; i >= 0; i = i - 1)
							begin
								// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:97:21
								if (core_req_valid[i]) begin
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:98:25
									per_bank_line_addr_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] = core_req_line_addr[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)];
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:99:25
									per_bank_rw_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = core_req_rw[i];
								end
							end
					end
				end
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:105:17
					assign core_req_line_match[i] = (core_req_line_addr[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] == per_bank_line_addr_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)]) && (core_req_rw[i] == per_bank_rw_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]]);
				end
				if (NUM_PORTS < NUM_REQS) begin : genblk2
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:111:17
					reg [((NUM_BANKS * NUM_PORTS) * NUM_REQS) - 1:0] req_select_table_r;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:113:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:114:21
						per_bank_core_req_valid_r = 0;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:115:21
						per_bank_core_req_pmask_r = 0;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:116:21
						per_bank_core_req_rw_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:117:21
						per_bank_core_req_addr_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:118:21
						per_bank_core_req_wsel_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:119:21
						per_bank_core_req_byteen_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:120:21
						per_bank_core_req_data_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:121:21
						per_bank_core_req_tag_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:122:21
						per_bank_core_req_tid_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:123:21
						req_select_table_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:125:21
						begin : sv2v_autoblock_2
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:125:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:125:26
							for (i = NUM_REQS - 1; i >= 0; i = i - 1)
								begin
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:126:25
									if (core_req_valid[i]) begin
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:127:29
										per_bank_core_req_valid_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = 1;
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:128:29
										per_bank_core_req_pmask_r[(core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)] = core_req_line_match[i];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:129:29
										per_bank_core_req_wsel_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)+:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)] = core_req_wsel[i * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)+:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:130:29
										per_bank_core_req_byteen_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * WORD_SIZE+:WORD_SIZE] = core_req_byteen[i * WORD_SIZE+:WORD_SIZE];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:131:29
										per_bank_core_req_data_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * (8 * WORD_SIZE)+:8 * WORD_SIZE] = core_req_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:132:29
										per_bank_core_req_tid_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)] = sv2v_cast_CC627_signed(i);
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:133:29
										per_bank_core_req_tag_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * CORE_TAG_WIDTH+:CORE_TAG_WIDTH] = core_req_tag[i * CORE_TAG_WIDTH+:CORE_TAG_WIDTH];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:134:29
										per_bank_core_req_rw_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = core_req_rw[i];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:135:29
										per_bank_core_req_addr_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] = core_req_line_addr[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:136:29
										req_select_table_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * NUM_REQS+:NUM_REQS] = 1 << i;
									end
								end
						end
					end
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:141:17
					always @(*)
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:142:21
						begin : sv2v_autoblock_3
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:142:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:142:26
							for (i = 0; i < NUM_REQS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:143:25
									core_req_ready_r[i] = (per_bank_core_req_ready[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] && core_req_line_match[i]) && req_select_table_r[(((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * NUM_REQS) + i];
								end
						end
				end
				else begin : genblk2
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:151:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:152:21
						per_bank_core_req_valid_r = 0;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:153:21
						per_bank_core_req_pmask_r = 0;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:154:21
						per_bank_core_req_rw_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:155:21
						per_bank_core_req_addr_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:156:21
						per_bank_core_req_wsel_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:157:21
						per_bank_core_req_byteen_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:158:21
						per_bank_core_req_data_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:159:21
						per_bank_core_req_tag_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:160:21
						per_bank_core_req_tid_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:162:21
						begin : sv2v_autoblock_4
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:162:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:162:26
							for (i = NUM_REQS - 1; i >= 0; i = i - 1)
								begin
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:163:25
									if (core_req_valid[i]) begin
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:164:29
										per_bank_core_req_valid_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = 1;
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:165:29
										per_bank_core_req_pmask_r[(core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)] = core_req_line_match[i];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:166:29
										per_bank_core_req_wsel_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)+:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)] = core_req_wsel[i * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)+:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:167:29
										per_bank_core_req_byteen_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * WORD_SIZE+:WORD_SIZE] = core_req_byteen[i * WORD_SIZE+:WORD_SIZE];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:168:29
										per_bank_core_req_data_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * (8 * WORD_SIZE)+:8 * WORD_SIZE] = core_req_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:169:29
										per_bank_core_req_tid_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)] = sv2v_cast_CC627_signed(i);
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:170:29
										per_bank_core_req_tag_r[((core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS) + (i % NUM_PORTS)) * CORE_TAG_WIDTH+:CORE_TAG_WIDTH] = core_req_tag[i * CORE_TAG_WIDTH+:CORE_TAG_WIDTH];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:171:29
										per_bank_core_req_rw_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = core_req_rw[i];
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:172:29
										per_bank_core_req_addr_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] = core_req_line_addr[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)];
									end
								end
						end
					end
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:177:17
					always @(*)
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:178:21
						begin : sv2v_autoblock_5
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:178:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:178:26
							for (i = 0; i < NUM_REQS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:179:25
									core_req_ready_r[i] = per_bank_core_req_ready[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] && core_req_line_match[i];
								end
						end
				end
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:187:13
				always @(*) begin
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:188:17
					per_bank_core_req_valid_r = 0;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:189:17
					per_bank_core_req_rw_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:190:17
					per_bank_core_req_addr_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:191:17
					per_bank_core_req_wsel_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:192:17
					per_bank_core_req_byteen_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:193:17
					per_bank_core_req_data_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:194:17
					per_bank_core_req_tag_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:195:17
					per_bank_core_req_tid_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:197:17
					begin : sv2v_autoblock_6
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:197:22
						integer i;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:197:22
						for (i = NUM_REQS - 1; i >= 0; i = i - 1)
							begin
								// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:198:21
								if (core_req_valid[i]) begin
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:199:25
									per_bank_core_req_valid_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = 1;
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:200:25
									per_bank_core_req_rw_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = core_req_rw[i];
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:201:25
									per_bank_core_req_addr_r[core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] = core_req_line_addr[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)];
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:202:25
									per_bank_core_req_wsel_r[($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1) * (core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1) * NUM_PORTS] = core_req_wsel[i * ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)+:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)];
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:203:25
									per_bank_core_req_byteen_r[WORD_SIZE * (core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:WORD_SIZE * NUM_PORTS] = core_req_byteen[i * WORD_SIZE+:WORD_SIZE];
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:204:25
									per_bank_core_req_data_r[(8 * WORD_SIZE) * (core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:(8 * WORD_SIZE) * NUM_PORTS] = core_req_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE];
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:205:25
									per_bank_core_req_tag_r[CORE_TAG_WIDTH * (core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:CORE_TAG_WIDTH * NUM_PORTS] = core_req_tag[i * CORE_TAG_WIDTH+:CORE_TAG_WIDTH];
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:206:25
									per_bank_core_req_tid_r[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (core_req_bid[i * ($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS] = sv2v_cast_CC627_signed(i);
								end
							end
					end
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:210:17
					per_bank_core_req_pmask_r = per_bank_core_req_valid_r;
				end
				if (NUM_BANKS > 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:214:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:215:21
						core_req_ready_r = 0;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:216:21
						begin : sv2v_autoblock_7
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:216:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:216:26
							for (i = 0; i < NUM_BANKS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:217:25
									if (per_bank_core_req_valid_r[i])
										// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:218:29
										core_req_ready_r[per_bank_core_req_tid_r[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS]] = per_bank_core_req_ready[i];
								end
						end
					end
				end
				else begin : genblk1
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:223:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:224:21
						core_req_ready_r = 0;
						// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:225:21
						core_req_ready_r[per_bank_core_req_tid_r[0+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS]] = per_bank_core_req_ready;
					end
				end
			end
		end
		else begin : genblk3
			if (NUM_BANKS > 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:233:13
				always @(*) begin
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:234:17
					per_bank_core_req_valid_r = 0;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:235:17
					per_bank_core_req_rw_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:236:17
					per_bank_core_req_addr_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:237:17
					per_bank_core_req_wsel_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:238:17
					per_bank_core_req_byteen_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:239:17
					per_bank_core_req_data_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:240:17
					per_bank_core_req_tag_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:241:17
					per_bank_core_req_tid_r = 1'sbx;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:242:17
					per_bank_core_req_valid_r[core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = core_req_valid;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:243:17
					per_bank_core_req_rw_r[core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]] = core_req_rw;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:244:17
					per_bank_core_req_addr_r[core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] = core_req_line_addr;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:245:17
					per_bank_core_req_wsel_r[($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1) * (core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1) * NUM_PORTS] = core_req_wsel;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:246:17
					per_bank_core_req_byteen_r[WORD_SIZE * (core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:WORD_SIZE * NUM_PORTS] = core_req_byteen;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:247:17
					per_bank_core_req_data_r[(8 * WORD_SIZE) * (core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:(8 * WORD_SIZE) * NUM_PORTS] = core_req_data;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:248:17
					per_bank_core_req_tag_r[CORE_TAG_WIDTH * (core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:CORE_TAG_WIDTH * NUM_PORTS] = core_req_tag;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:249:17
					per_bank_core_req_tid_r[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)] * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS] = 0;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:250:17
					core_req_ready_r = per_bank_core_req_ready[core_req_bid[0+:($clog2(NUM_BANKS) > 0 ? $clog2(NUM_BANKS) : 1)]];
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:252:17
					per_bank_core_req_pmask_r = per_bank_core_req_valid_r;
				end
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:256:13
				always @(*) begin
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:257:17
					per_bank_core_req_valid_r = core_req_valid;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:258:17
					per_bank_core_req_rw_r = core_req_rw;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:259:17
					per_bank_core_req_addr_r = core_req_line_addr;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:260:17
					per_bank_core_req_wsel_r = core_req_wsel;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:261:17
					per_bank_core_req_byteen_r = core_req_byteen;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:262:17
					per_bank_core_req_data_r = core_req_data;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:263:17
					per_bank_core_req_tag_r = core_req_tag;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:264:17
					per_bank_core_req_tid_r = 0;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:265:17
					core_req_ready_r = per_bank_core_req_ready;
					// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:267:17
					per_bank_core_req_pmask_r = per_bank_core_req_valid_r;
				end
			end
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:273:5
	assign per_bank_core_req_valid = per_bank_core_req_valid_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:274:5
	assign per_bank_core_req_pmask = per_bank_core_req_pmask_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:275:5
	assign per_bank_core_req_rw = per_bank_core_req_rw_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:276:5
	assign per_bank_core_req_addr = per_bank_core_req_addr_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:277:5
	assign per_bank_core_req_wsel = per_bank_core_req_wsel_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:278:5
	assign per_bank_core_req_byteen = per_bank_core_req_byteen_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:279:5
	assign per_bank_core_req_data = per_bank_core_req_data_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:280:5
	assign per_bank_core_req_tag = per_bank_core_req_tag_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:281:5
	assign per_bank_core_req_tid = per_bank_core_req_tid_r;
	// Trace: ../../rtl/cache/VX_core_req_bank_sel.sv:282:5
	assign core_req_ready = core_req_ready_r;
endmodule
module VX_core_rsp_merge (
	clk,
	reset,
	per_bank_core_rsp_valid,
	per_bank_core_rsp_pmask,
	per_bank_core_rsp_data,
	per_bank_core_rsp_tid,
	per_bank_core_rsp_tag,
	per_bank_core_rsp_ready,
	core_rsp_valid,
	core_rsp_tmask,
	core_rsp_tag,
	core_rsp_data,
	core_rsp_ready
);
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:4:15
	parameter CACHE_ID = 0;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:7:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:9:15
	parameter NUM_BANKS = 1;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:11:15
	parameter NUM_PORTS = 1;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:13:15
	parameter WORD_SIZE = 1;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:15:15
	parameter CORE_TAG_WIDTH = 1;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:17:15
	parameter CORE_TAG_ID_BITS = 0;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:19:15
	parameter OUT_REG = 0;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:21:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:22:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:25:5
	input wire [NUM_BANKS - 1:0] per_bank_core_rsp_valid;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:26:5
	input wire [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_pmask;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:27:5
	input wire [((NUM_BANKS * NUM_PORTS) * (8 * WORD_SIZE)) - 1:0] per_bank_core_rsp_data;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:28:5
	input wire [((NUM_BANKS * NUM_PORTS) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] per_bank_core_rsp_tid;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:29:5
	input wire [((NUM_BANKS * NUM_PORTS) * CORE_TAG_WIDTH) - 1:0] per_bank_core_rsp_tag;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:30:5
	output wire [NUM_BANKS - 1:0] per_bank_core_rsp_ready;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:33:5
	output wire [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_valid;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:34:5
	output wire [NUM_REQS - 1:0] core_rsp_tmask;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:35:5
	output wire [((CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) * CORE_TAG_WIDTH) - 1:0] core_rsp_tag;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:36:5
	output wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_rsp_data;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:37:5
	input wire [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_ready;
	// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:41:5
	function automatic signed [(NUM_PORTS > 1 ? $clog2(NUM_PORTS) : 1) - 1:0] sv2v_cast_B86A1_signed;
		input reg signed [(NUM_PORTS > 1 ? $clog2(NUM_PORTS) : 1) - 1:0] inp;
		sv2v_cast_B86A1_signed = inp;
	endfunction
	function automatic signed [$clog2(NUM_BANKS) - 1:0] sv2v_cast_748B1_signed;
		input reg signed [$clog2(NUM_BANKS) - 1:0] inp;
		sv2v_cast_748B1_signed = inp;
	endfunction
	generate
		if (NUM_BANKS > 1) begin : genblk1
			// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:43:9
			reg [NUM_REQS - 1:0] core_rsp_valid_unqual;
			// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:44:9
			reg [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_rsp_data_unqual;
			// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:45:9
			reg [NUM_BANKS - 1:0] per_bank_core_rsp_ready_r;
			if (CORE_TAG_ID_BITS != 0) begin : genblk1
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:53:13
				wire [CORE_TAG_WIDTH - 1:0] core_rsp_tag_unqual;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:54:13
				wire core_rsp_ready_unqual;
				if (NUM_PORTS > 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:58:17
					reg [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_sent_r;
					reg [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_sent;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:59:17
					wire [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_sent_n;
					genvar i;
					for (i = 0; i < NUM_BANKS; i = i + 1) begin : genblk1
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:62:21
						assign per_bank_core_rsp_sent_n[i * NUM_PORTS+:NUM_PORTS] = per_bank_core_rsp_sent_r[i * NUM_PORTS+:NUM_PORTS] | per_bank_core_rsp_sent[i * NUM_PORTS+:NUM_PORTS];
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:65:17
					always @(posedge clk)
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:66:21
						if (reset)
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:67:25
							per_bank_core_rsp_sent_r <= 1'sb0;
						else
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:69:25
							begin : sv2v_autoblock_1
								// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:69:30
								integer i;
								// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:69:30
								for (i = 0; i < NUM_BANKS; i = i + 1)
									begin
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:70:29
										if (per_bank_core_rsp_sent_n[i * NUM_PORTS+:NUM_PORTS] == per_bank_core_rsp_pmask[i * NUM_PORTS+:NUM_PORTS])
											// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:71:33
											per_bank_core_rsp_sent_r[i * NUM_PORTS+:NUM_PORTS] <= 1'sb0;
										else
											// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:73:33
											per_bank_core_rsp_sent_r[i * NUM_PORTS+:NUM_PORTS] <= per_bank_core_rsp_sent_n[i * NUM_PORTS+:NUM_PORTS];
									end
							end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:79:17
					wire [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_valid_p;
					for (i = 0; i < NUM_BANKS; i = i + 1) begin : genblk2
						genvar p;
						for (p = 0; p < NUM_PORTS; p = p + 1) begin : genblk1
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:82:25
							assign per_bank_core_rsp_valid_p[(i * NUM_PORTS) + p] = (per_bank_core_rsp_valid[i] && per_bank_core_rsp_pmask[(i * NUM_PORTS) + p]) && !per_bank_core_rsp_sent_r[(i * NUM_PORTS) + p];
						end
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:88:17
					VX_find_first #(
						.N(NUM_BANKS * NUM_PORTS),
						.DATAW(CORE_TAG_WIDTH)
					) find_first(
						.valid_i(per_bank_core_rsp_valid_p),
						.data_i(per_bank_core_rsp_tag),
						.data_o(core_rsp_tag_unqual)
					);
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:98:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:99:21
						core_rsp_valid_unqual = 0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:100:21
						core_rsp_data_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:101:21
						per_bank_core_rsp_sent = 0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:103:21
						begin : sv2v_autoblock_2
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:103:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:103:26
							for (i = 0; i < NUM_BANKS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:104:25
									begin : sv2v_autoblock_3
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:104:30
										integer p;
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:104:30
										for (p = 0; p < NUM_PORTS; p = p + 1)
											begin
												// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:105:29
												if (((per_bank_core_rsp_valid[i] && per_bank_core_rsp_pmask[(i * NUM_PORTS) + p]) && !per_bank_core_rsp_sent_r[(i * NUM_PORTS) + p]) && (per_bank_core_rsp_tag[(((i * NUM_PORTS) + p) * CORE_TAG_WIDTH) + (CORE_TAG_ID_BITS - 1)-:CORE_TAG_ID_BITS] == core_rsp_tag_unqual[CORE_TAG_ID_BITS - 1:0])) begin
													// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:109:33
													core_rsp_valid_unqual[per_bank_core_rsp_tid[((i * NUM_PORTS) + p) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)]] = 1;
													// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:110:33
													core_rsp_data_unqual[per_bank_core_rsp_tid[((i * NUM_PORTS) + p) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)] * (8 * WORD_SIZE)+:8 * WORD_SIZE] = per_bank_core_rsp_data[((i * NUM_PORTS) + p) * (8 * WORD_SIZE)+:8 * WORD_SIZE];
													// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:111:33
													per_bank_core_rsp_sent[(i * NUM_PORTS) + p] = core_rsp_ready_unqual;
												end
											end
									end
								end
						end
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:117:17
					always @(*)
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:118:21
						begin : sv2v_autoblock_4
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:118:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:118:26
							for (i = 0; i < NUM_BANKS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:119:25
									per_bank_core_rsp_ready_r[i] = per_bank_core_rsp_sent_n[i * NUM_PORTS+:NUM_PORTS] == per_bank_core_rsp_pmask[i * NUM_PORTS+:NUM_PORTS];
								end
						end
				end
				else begin : genblk1
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:127:17
					VX_find_first #(
						.N(NUM_BANKS),
						.DATAW(CORE_TAG_WIDTH)
					) find_first(
						.valid_i(per_bank_core_rsp_valid),
						.data_i(per_bank_core_rsp_tag),
						.data_o(core_rsp_tag_unqual)
					);
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:137:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:138:21
						core_rsp_valid_unqual = 0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:139:21
						core_rsp_data_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:140:21
						per_bank_core_rsp_ready_r = 0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:142:21
						begin : sv2v_autoblock_5
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:142:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:142:26
							for (i = 0; i < NUM_BANKS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:143:25
									if (per_bank_core_rsp_valid[i] && (per_bank_core_rsp_tag[((i * NUM_PORTS) * CORE_TAG_WIDTH) + (CORE_TAG_ID_BITS - 1)-:CORE_TAG_ID_BITS] == core_rsp_tag_unqual[CORE_TAG_ID_BITS - 1:0])) begin
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:145:29
										core_rsp_valid_unqual[per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS]] = 1;
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:146:29
										core_rsp_data_unqual[per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS] * (8 * WORD_SIZE)+:8 * WORD_SIZE] = per_bank_core_rsp_data[(8 * WORD_SIZE) * (i * NUM_PORTS)+:(8 * WORD_SIZE) * NUM_PORTS];
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:147:29
										per_bank_core_rsp_ready_r[i] = core_rsp_ready_unqual;
									end
								end
						end
					end
				end
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:153:13
				wire core_rsp_valid_any = |per_bank_core_rsp_valid;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:155:13
				VX_skid_buffer #(
					.DATAW((NUM_REQS + CORE_TAG_WIDTH) + (NUM_REQS * (8 * WORD_SIZE))),
					.PASSTHRU(0 == OUT_REG)
				) out_sbuf(
					.clk(clk),
					.reset(reset),
					.valid_in(core_rsp_valid_any),
					.data_in({core_rsp_valid_unqual, core_rsp_tag_unqual, core_rsp_data_unqual}),
					.ready_in(core_rsp_ready_unqual),
					.valid_out(core_rsp_valid),
					.data_out({core_rsp_tmask, core_rsp_tag, core_rsp_data}),
					.ready_out(core_rsp_ready)
				);
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:171:13
				reg [(NUM_REQS * CORE_TAG_WIDTH) - 1:0] core_rsp_tag_unqual;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:172:13
				wire [NUM_REQS - 1:0] core_rsp_ready_unqual;
				if (NUM_PORTS > 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:176:17
					reg [(NUM_REQS * ((NUM_PORTS > 1 ? $clog2(NUM_PORTS) : 1) + $clog2(NUM_BANKS))) - 1:0] bank_select_table;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:178:17
					reg [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_sent_r;
					reg [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_sent;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:179:17
					wire [(NUM_BANKS * NUM_PORTS) - 1:0] per_bank_core_rsp_sent_n;
					genvar i;
					for (i = 0; i < NUM_BANKS; i = i + 1) begin : genblk1
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:182:21
						assign per_bank_core_rsp_sent_n[i * NUM_PORTS+:NUM_PORTS] = per_bank_core_rsp_sent_r[i * NUM_PORTS+:NUM_PORTS] | per_bank_core_rsp_sent[i * NUM_PORTS+:NUM_PORTS];
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:185:17
					always @(posedge clk)
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:186:21
						if (reset)
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:187:25
							per_bank_core_rsp_sent_r <= 1'sb0;
						else
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:189:25
							begin : sv2v_autoblock_6
								// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:189:30
								integer i;
								// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:189:30
								for (i = 0; i < NUM_BANKS; i = i + 1)
									begin
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:190:29
										if (per_bank_core_rsp_sent_n[i * NUM_PORTS+:NUM_PORTS] == per_bank_core_rsp_pmask[i * NUM_PORTS+:NUM_PORTS])
											// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:191:33
											per_bank_core_rsp_sent_r[i * NUM_PORTS+:NUM_PORTS] <= 1'sb0;
										else
											// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:193:33
											per_bank_core_rsp_sent_r[i * NUM_PORTS+:NUM_PORTS] <= per_bank_core_rsp_sent_n[i * NUM_PORTS+:NUM_PORTS];
									end
							end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:199:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:200:21
						core_rsp_valid_unqual = 1'sb0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:201:21
						core_rsp_tag_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:202:21
						core_rsp_data_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:203:21
						bank_select_table = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:205:21
						begin : sv2v_autoblock_7
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:205:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:205:26
							for (i = NUM_BANKS - 1; i >= 0; i = i - 1)
								begin
									// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:206:25
									begin : sv2v_autoblock_8
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:206:30
										integer p;
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:206:30
										for (p = 0; p < NUM_PORTS; p = p + 1)
											begin
												// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:207:29
												if ((per_bank_core_rsp_valid[i] && per_bank_core_rsp_pmask[(i * NUM_PORTS) + p]) && !per_bank_core_rsp_sent_r[(i * NUM_PORTS) + p]) begin
													// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:210:33
													core_rsp_valid_unqual[per_bank_core_rsp_tid[((i * NUM_PORTS) + p) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)]] = 1;
													// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:211:33
													core_rsp_tag_unqual[per_bank_core_rsp_tid[((i * NUM_PORTS) + p) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)] * CORE_TAG_WIDTH+:CORE_TAG_WIDTH] = per_bank_core_rsp_tag[((i * NUM_PORTS) + p) * CORE_TAG_WIDTH+:CORE_TAG_WIDTH];
													// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:212:33
													core_rsp_data_unqual[per_bank_core_rsp_tid[((i * NUM_PORTS) + p) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)] * (8 * WORD_SIZE)+:8 * WORD_SIZE] = per_bank_core_rsp_data[((i * NUM_PORTS) + p) * (8 * WORD_SIZE)+:8 * WORD_SIZE];
													// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:213:33
													bank_select_table[per_bank_core_rsp_tid[((i * NUM_PORTS) + p) * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)] * ((NUM_PORTS > 1 ? $clog2(NUM_PORTS) : 1) + $clog2(NUM_BANKS))+:(NUM_PORTS > 1 ? $clog2(NUM_PORTS) : 1) + $clog2(NUM_BANKS)] = {sv2v_cast_B86A1_signed(p), sv2v_cast_748B1_signed(i)};
												end
											end
									end
								end
						end
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:219:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:220:21
						per_bank_core_rsp_sent = 1'sb0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:221:21
						begin : sv2v_autoblock_9
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:221:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:221:26
							for (i = 0; i < NUM_REQS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:222:25
									if (core_rsp_valid_unqual[i])
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:223:29
										per_bank_core_rsp_sent[(bank_select_table[i * ((NUM_PORTS > 1 ? $clog2(NUM_PORTS) : 1) + $clog2(NUM_BANKS))+:$clog2(NUM_BANKS)] * NUM_PORTS) + bank_select_table[(i * ((NUM_PORTS > 1 ? $clog2(NUM_PORTS) : 1) + $clog2(NUM_BANKS))) + $clog2(NUM_BANKS)+:(NUM_PORTS > 1 ? $clog2(NUM_PORTS) : 1)]] = core_rsp_ready_unqual[i];
								end
						end
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:228:17
					always @(*)
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:229:21
						begin : sv2v_autoblock_10
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:229:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:229:26
							for (i = 0; i < NUM_BANKS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:230:25
									per_bank_core_rsp_ready_r[i] = per_bank_core_rsp_sent_n[i * NUM_PORTS+:NUM_PORTS] == per_bank_core_rsp_pmask[i * NUM_PORTS+:NUM_PORTS];
								end
						end
				end
				else begin : genblk1
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:237:17
					reg [(NUM_REQS * NUM_BANKS) - 1:0] bank_select_table;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:239:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:240:21
						core_rsp_valid_unqual = 0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:241:21
						core_rsp_tag_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:242:21
						core_rsp_data_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:243:21
						bank_select_table = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:245:21
						begin : sv2v_autoblock_11
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:245:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:245:26
							for (i = NUM_BANKS - 1; i >= 0; i = i - 1)
								begin
									// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:246:25
									if (per_bank_core_rsp_valid[i]) begin
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:247:29
										core_rsp_valid_unqual[per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS]] = 1;
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:248:29
										core_rsp_tag_unqual[per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS] * CORE_TAG_WIDTH+:CORE_TAG_WIDTH] = per_bank_core_rsp_tag[CORE_TAG_WIDTH * (i * NUM_PORTS)+:CORE_TAG_WIDTH * NUM_PORTS];
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:249:29
										core_rsp_data_unqual[per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS] * (8 * WORD_SIZE)+:8 * WORD_SIZE] = per_bank_core_rsp_data[(8 * WORD_SIZE) * (i * NUM_PORTS)+:(8 * WORD_SIZE) * NUM_PORTS];
										// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:250:29
										bank_select_table[per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS] * NUM_BANKS+:NUM_BANKS] = 1 << i;
									end
								end
						end
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:255:17
					always @(*)
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:256:21
						begin : sv2v_autoblock_12
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:256:26
							integer i;
							// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:256:26
							for (i = 0; i < NUM_BANKS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:257:25
									per_bank_core_rsp_ready_r[i] = core_rsp_ready_unqual[per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS]] && bank_select_table[(per_bank_core_rsp_tid[(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * (i * NUM_PORTS)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1) * NUM_PORTS] * NUM_BANKS) + i];
								end
						end
				end
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk2
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:264:17
					VX_skid_buffer #(
						.DATAW(CORE_TAG_WIDTH + (8 * WORD_SIZE)),
						.PASSTHRU(0 == OUT_REG)
					) out_sbuf(
						.clk(clk),
						.reset(reset),
						.valid_in(core_rsp_valid_unqual[i]),
						.data_in({core_rsp_tag_unqual[i * CORE_TAG_WIDTH+:CORE_TAG_WIDTH], core_rsp_data_unqual[i * (8 * WORD_SIZE)+:8 * WORD_SIZE]}),
						.ready_in(core_rsp_ready_unqual[i]),
						.valid_out(core_rsp_valid[i]),
						.data_out({core_rsp_tag[i * CORE_TAG_WIDTH+:CORE_TAG_WIDTH], core_rsp_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE]}),
						.ready_out(core_rsp_ready[i])
					);
				end
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:279:13
				assign core_rsp_tmask = core_rsp_valid;
			end
			// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:283:9
			assign per_bank_core_rsp_ready = per_bank_core_rsp_ready_r;
		end
		else begin : genblk1
			if (NUM_REQS > 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:293:13
				reg [((CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) * CORE_TAG_WIDTH) - 1:0] core_rsp_tag_unqual;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:294:13
				reg [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_rsp_data_unqual;
				if (CORE_TAG_ID_BITS != 0) begin : genblk1
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:298:17
					reg [NUM_REQS - 1:0] core_rsp_tmask_unqual;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:300:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:301:21
						core_rsp_tmask_unqual = 0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:302:21
						core_rsp_tmask_unqual[per_bank_core_rsp_tid] = per_bank_core_rsp_valid;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:304:21
						core_rsp_tag_unqual = per_bank_core_rsp_tag;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:306:21
						core_rsp_data_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:307:21
						core_rsp_data_unqual[per_bank_core_rsp_tid * (8 * WORD_SIZE)+:8 * WORD_SIZE] = per_bank_core_rsp_data;
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:310:17
					assign core_rsp_valid = per_bank_core_rsp_valid;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:311:17
					assign core_rsp_tmask = core_rsp_tmask_unqual;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:312:17
					assign per_bank_core_rsp_ready = core_rsp_ready;
				end
				else begin : genblk1
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:316:17
					reg [(CORE_TAG_ID_BITS != 0 ? 1 : NUM_REQS) - 1:0] core_rsp_valid_unqual;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:318:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:319:21
						core_rsp_valid_unqual = 0;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:320:21
						core_rsp_valid_unqual[per_bank_core_rsp_tid] = per_bank_core_rsp_valid;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:322:21
						core_rsp_tag_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:323:21
						core_rsp_tag_unqual[per_bank_core_rsp_tid * CORE_TAG_WIDTH+:CORE_TAG_WIDTH] = per_bank_core_rsp_tag;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:325:21
						core_rsp_data_unqual = 1'sbx;
						// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:326:21
						core_rsp_data_unqual[per_bank_core_rsp_tid * (8 * WORD_SIZE)+:8 * WORD_SIZE] = per_bank_core_rsp_data;
					end
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:329:17
					assign core_rsp_valid = core_rsp_valid_unqual;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:330:17
					assign core_rsp_tmask = core_rsp_valid_unqual;
					// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:331:17
					assign per_bank_core_rsp_ready = core_rsp_ready[per_bank_core_rsp_tid];
				end
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:335:13
				assign core_rsp_tag = core_rsp_tag_unqual;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:336:13
				assign core_rsp_data = core_rsp_data_unqual;
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:341:13
				assign core_rsp_valid = per_bank_core_rsp_valid;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:342:13
				assign core_rsp_tmask = per_bank_core_rsp_valid;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:343:13
				assign core_rsp_tag = per_bank_core_rsp_tag;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:344:13
				assign core_rsp_data = per_bank_core_rsp_data;
				// Trace: ../../rtl/cache/VX_core_rsp_merge.sv:345:13
				assign per_bank_core_rsp_ready = core_rsp_ready;
			end
		end
	endgenerate
endmodule
module VX_data_access (
	clk,
	reset,
	req_id,
	stall,
	read,
	fill,
	write,
	addr,
	wsel,
	pmask,
	byteen,
	fill_data,
	write_data,
	read_data
);
	// Trace: ../../rtl/cache/VX_data_access.sv:4:15
	parameter CACHE_ID = 0;
	// Trace: ../../rtl/cache/VX_data_access.sv:5:15
	parameter BANK_ID = 0;
	// Trace: ../../rtl/cache/VX_data_access.sv:7:15
	parameter CACHE_SIZE = 1;
	// Trace: ../../rtl/cache/VX_data_access.sv:9:15
	parameter CACHE_LINE_SIZE = 1;
	// Trace: ../../rtl/cache/VX_data_access.sv:11:15
	parameter NUM_BANKS = 1;
	// Trace: ../../rtl/cache/VX_data_access.sv:13:15
	parameter NUM_PORTS = 1;
	// Trace: ../../rtl/cache/VX_data_access.sv:15:15
	parameter WORD_SIZE = 1;
	// Trace: ../../rtl/cache/VX_data_access.sv:17:15
	parameter WRITE_ENABLE = 1;
	// Trace: ../../rtl/cache/VX_data_access.sv:19:15
	parameter WORD_SELECT_BITS = ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1);
	// Trace: ../../rtl/cache/VX_data_access.sv:21:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_data_access.sv:22:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_data_access.sv:25:5
	input wire [43:0] req_id;
	// Trace: ../../rtl/cache/VX_data_access.sv:28:5
	input wire stall;
	// Trace: ../../rtl/cache/VX_data_access.sv:30:5
	input wire read;
	// Trace: ../../rtl/cache/VX_data_access.sv:31:5
	input wire fill;
	// Trace: ../../rtl/cache/VX_data_access.sv:32:5
	input wire write;
	// Trace: ../../rtl/cache/VX_data_access.sv:33:5
	input wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr;
	// Trace: ../../rtl/cache/VX_data_access.sv:34:5
	input wire [(NUM_PORTS * WORD_SELECT_BITS) - 1:0] wsel;
	// Trace: ../../rtl/cache/VX_data_access.sv:35:5
	input wire [NUM_PORTS - 1:0] pmask;
	// Trace: ../../rtl/cache/VX_data_access.sv:36:5
	input wire [(NUM_PORTS * WORD_SIZE) - 1:0] byteen;
	// Trace: ../../rtl/cache/VX_data_access.sv:37:5
	input wire [((CACHE_LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] fill_data;
	// Trace: ../../rtl/cache/VX_data_access.sv:38:5
	input wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] write_data;
	// Trace: ../../rtl/cache/VX_data_access.sv:39:5
	output wire [(NUM_PORTS * (8 * WORD_SIZE)) - 1:0] read_data;
	// Trace: ../../rtl/cache/VX_data_access.sv:48:5
	localparam BYTEENW = (WRITE_ENABLE ? CACHE_LINE_SIZE : 1);
	// Trace: ../../rtl/cache/VX_data_access.sv:50:5
	wire [((CACHE_LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] rdata;
	// Trace: ../../rtl/cache/VX_data_access.sv:51:5
	wire [((CACHE_LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] wdata;
	// Trace: ../../rtl/cache/VX_data_access.sv:52:5
	wire [BYTEENW - 1:0] wren;
	// Trace: ../../rtl/cache/VX_data_access.sv:54:5
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0] line_addr = addr[$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0];
	// Trace: ../../rtl/cache/VX_data_access.sv:56:5
	generate
		if (WRITE_ENABLE) begin : genblk1
			if ((CACHE_LINE_SIZE / WORD_SIZE) > 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_data_access.sv:58:13
				reg [((CACHE_LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] wdata_r;
				// Trace: ../../rtl/cache/VX_data_access.sv:59:13
				reg [((CACHE_LINE_SIZE / WORD_SIZE) * WORD_SIZE) - 1:0] wren_r;
				if (NUM_PORTS > 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_data_access.sv:61:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_data_access.sv:62:21
						wdata_r = 1'sbx;
						// Trace: ../../rtl/cache/VX_data_access.sv:63:21
						wren_r = 0;
						// Trace: ../../rtl/cache/VX_data_access.sv:64:21
						begin : sv2v_autoblock_1
							// Trace: ../../rtl/cache/VX_data_access.sv:64:26
							integer i;
							// Trace: ../../rtl/cache/VX_data_access.sv:64:26
							for (i = 0; i < NUM_PORTS; i = i + 1)
								begin
									// Trace: ../../rtl/cache/VX_data_access.sv:65:25
									if (pmask[i]) begin
										// Trace: ../../rtl/cache/VX_data_access.sv:66:29
										wdata_r[wsel[i * WORD_SELECT_BITS+:WORD_SELECT_BITS] * (8 * WORD_SIZE)+:8 * WORD_SIZE] = write_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE];
										// Trace: ../../rtl/cache/VX_data_access.sv:67:29
										wren_r[wsel[i * WORD_SELECT_BITS+:WORD_SELECT_BITS] * WORD_SIZE+:WORD_SIZE] = byteen[i * WORD_SIZE+:WORD_SIZE];
									end
								end
						end
					end
				end
				else begin : genblk1
					// Trace: ../../rtl/cache/VX_data_access.sv:73:17
					always @(*) begin
						// Trace: ../../rtl/cache/VX_data_access.sv:74:21
						wdata_r = {CACHE_LINE_SIZE / WORD_SIZE {write_data}};
						// Trace: ../../rtl/cache/VX_data_access.sv:75:21
						wren_r = 0;
						// Trace: ../../rtl/cache/VX_data_access.sv:76:21
						wren_r[wsel * WORD_SIZE+:WORD_SIZE] = byteen;
					end
				end
				// Trace: ../../rtl/cache/VX_data_access.sv:79:13
				assign wdata = (write ? wdata_r : fill_data);
				// Trace: ../../rtl/cache/VX_data_access.sv:80:13
				assign wren = (write ? wren_r : {BYTEENW {fill}});
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_data_access.sv:84:13
				assign wdata = (write ? write_data : fill_data);
				// Trace: ../../rtl/cache/VX_data_access.sv:85:13
				assign wren = (write ? byteen : {BYTEENW {fill}});
			end
		end
		else begin : genblk1
			// Trace: ../../rtl/cache/VX_data_access.sv:92:9
			assign wdata = fill_data;
			// Trace: ../../rtl/cache/VX_data_access.sv:93:9
			assign wren = fill;
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_data_access.sv:96:5
	VX_sp_ram #(
		.DATAW(8 * CACHE_LINE_SIZE),
		.SIZE((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE),
		.BYTEENW(BYTEENW),
		.NO_RWCHECK(1)
	) data_store(
		.clk(clk),
		.addr(line_addr),
		.wren(wren),
		.wdata(wdata),
		.rdata(rdata)
	);
	// Trace: ../../rtl/cache/VX_data_access.sv:109:5
	generate
		if ((CACHE_LINE_SIZE / WORD_SIZE) > 1) begin : genblk2
			genvar i;
			for (i = 0; i < NUM_PORTS; i = i + 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_data_access.sv:111:13
				assign read_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE] = rdata[wsel[i * WORD_SELECT_BITS+:WORD_SELECT_BITS] * (8 * WORD_SIZE)+:8 * WORD_SIZE];
			end
		end
		else begin : genblk2
			// Trace: ../../rtl/cache/VX_data_access.sv:114:9
			assign read_data = rdata;
		end
	endgenerate
endmodule
module VX_flush_ctrl (
	clk,
	reset,
	addr_out,
	valid_out
);
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:5:15
	parameter CACHE_SIZE = 16384;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:7:15
	parameter CACHE_LINE_SIZE = 1;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:9:15
	parameter NUM_BANKS = 1;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:11:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:12:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:13:5
	output wire [$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0] addr_out;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:14:5
	output wire valid_out;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:16:5
	reg flush_enable;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:17:5
	reg [$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0] flush_ctr;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:19:5
	always @(posedge clk)
		// Trace: ../../rtl/cache/VX_flush_ctrl.sv:20:9
		if (reset) begin
			// Trace: ../../rtl/cache/VX_flush_ctrl.sv:21:13
			flush_enable <= 1;
			// Trace: ../../rtl/cache/VX_flush_ctrl.sv:22:13
			flush_ctr <= 0;
		end
		else
			// Trace: ../../rtl/cache/VX_flush_ctrl.sv:24:13
			if (flush_enable) begin
				// Trace: ../../rtl/cache/VX_flush_ctrl.sv:25:17
				if (flush_ctr == ((2 ** $clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE)) - 1))
					// Trace: ../../rtl/cache/VX_flush_ctrl.sv:26:21
					flush_enable <= 0;
				// Trace: ../../rtl/cache/VX_flush_ctrl.sv:28:17
				flush_ctr <= flush_ctr + 1;
			end
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:33:5
	assign addr_out = flush_ctr;
	// Trace: ../../rtl/cache/VX_flush_ctrl.sv:34:5
	assign valid_out = flush_enable;
endmodule
module VX_miss_resrv (
	clk,
	reset,
	deq_req_id,
	lkp_req_id,
	rel_req_id,
	allocate_valid,
	allocate_addr,
	allocate_data,
	allocate_id,
	allocate_ready,
	fill_valid,
	fill_id,
	fill_addr,
	lookup_valid,
	lookup_replay,
	lookup_id,
	lookup_addr,
	lookup_match,
	dequeue_valid,
	dequeue_id,
	dequeue_addr,
	dequeue_data,
	dequeue_ready,
	release_valid,
	release_id
);
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:4:15
	parameter CACHE_ID = 0;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:5:15
	parameter BANK_ID = 0;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:8:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:11:15
	parameter CACHE_LINE_SIZE = 1;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:13:15
	parameter NUM_BANKS = 1;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:15:15
	parameter NUM_PORTS = 1;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:17:15
	parameter WORD_SIZE = 1;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:19:15
	parameter MSHR_SIZE = 1;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:21:15
	parameter CORE_TAG_WIDTH = 1;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:23:15
	parameter MSHR_ADDR_WIDTH = $clog2(MSHR_SIZE);
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:25:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:26:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:29:5
	input wire [43:0] deq_req_id;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:30:5
	input wire [43:0] lkp_req_id;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:31:5
	input wire [43:0] rel_req_id;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:35:5
	input wire allocate_valid;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:36:5
	input wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] allocate_addr;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:37:5
	input wire [((((CORE_TAG_WIDTH + 1) + (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) + ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)) * NUM_PORTS) - 1:0] allocate_data;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:38:5
	output wire [MSHR_ADDR_WIDTH - 1:0] allocate_id;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:39:5
	output wire allocate_ready;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:42:5
	input wire fill_valid;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:43:5
	input wire [MSHR_ADDR_WIDTH - 1:0] fill_id;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:44:5
	output wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] fill_addr;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:47:5
	input wire lookup_valid;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:48:5
	input wire lookup_replay;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:49:5
	input wire [MSHR_ADDR_WIDTH - 1:0] lookup_id;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:50:5
	input wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] lookup_addr;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:51:5
	output wire lookup_match;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:54:5
	output wire dequeue_valid;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:55:5
	output wire [MSHR_ADDR_WIDTH - 1:0] dequeue_id;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:56:5
	output wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] dequeue_addr;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:57:5
	output wire [((((CORE_TAG_WIDTH + 1) + (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) + ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)) * NUM_PORTS) - 1:0] dequeue_data;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:58:5
	input wire dequeue_ready;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:61:5
	input wire release_valid;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:62:5
	input wire [MSHR_ADDR_WIDTH - 1:0] release_id;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:67:5
	reg [(MSHR_SIZE * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] addr_table;
	reg [(MSHR_SIZE * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] addr_table_n;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:68:5
	reg [MSHR_SIZE - 1:0] valid_table;
	reg [MSHR_SIZE - 1:0] valid_table_n;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:69:5
	reg [MSHR_SIZE - 1:0] ready_table;
	reg [MSHR_SIZE - 1:0] ready_table_n;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:71:5
	reg allocate_rdy_r;
	reg allocate_rdy_n;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:72:5
	reg [MSHR_ADDR_WIDTH - 1:0] allocate_id_r;
	reg [MSHR_ADDR_WIDTH - 1:0] allocate_id_n;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:74:5
	reg dequeue_val_r;
	reg dequeue_val_n;
	reg dequeue_val_x;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:75:5
	reg [MSHR_ADDR_WIDTH - 1:0] dequeue_id_r;
	reg [MSHR_ADDR_WIDTH - 1:0] dequeue_id_n;
	reg [MSHR_ADDR_WIDTH - 1:0] dequeue_id_x;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:77:5
	reg [MSHR_SIZE - 1:0] valid_table_x;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:78:5
	reg [MSHR_SIZE - 1:0] ready_table_x;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:80:5
	wire [MSHR_SIZE - 1:0] addr_matches;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:82:5
	wire allocate_fire = allocate_valid && allocate_ready;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:84:5
	wire dequeue_fire = dequeue_valid && dequeue_ready;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:86:5
	genvar i;
	generate
		for (i = 0; i < MSHR_SIZE; i = i + 1) begin : genblk1
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:87:9
			assign addr_matches[i] = addr_table[i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] == lookup_addr;
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:90:5
	always @(*) begin
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:91:9
		valid_table_x = valid_table;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:92:9
		ready_table_x = ready_table;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:93:9
		if (dequeue_fire)
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:94:13
			valid_table_x[dequeue_id] = 0;
		if (lookup_replay)
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:97:13
			ready_table_x = ready_table_x | addr_matches;
	end
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:101:5
	// rewrote reg-to-output bindings
	wire [MSHR_ADDR_WIDTH:1] sv2v_tmp_dequeue_sel_cnt_o;
	always @(*) dequeue_id_x = sv2v_tmp_dequeue_sel_cnt_o;
	wire [1:1] sv2v_tmp_dequeue_sel_valid_o;
	always @(*) dequeue_val_x = sv2v_tmp_dequeue_sel_valid_o;
	VX_lzc #(.N(MSHR_SIZE)) dequeue_sel(
		.in_i(valid_table_x & ready_table_x),
		.cnt_o(sv2v_tmp_dequeue_sel_cnt_o),
		.valid_o(sv2v_tmp_dequeue_sel_valid_o)
	);
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:109:5
	// rewrote reg-to-output bindings
	wire [MSHR_ADDR_WIDTH:1] sv2v_tmp_allocate_sel_cnt_o;
	always @(*) allocate_id_n = sv2v_tmp_allocate_sel_cnt_o;
	wire [1:1] sv2v_tmp_allocate_sel_valid_o;
	always @(*) allocate_rdy_n = sv2v_tmp_allocate_sel_valid_o;
	VX_lzc #(.N(MSHR_SIZE)) allocate_sel(
		.in_i(~valid_table_n),
		.cnt_o(sv2v_tmp_allocate_sel_cnt_o),
		.valid_o(sv2v_tmp_allocate_sel_valid_o)
	);
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:117:5
	always @(*) begin
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:118:9
		valid_table_n = valid_table_x;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:119:9
		ready_table_n = ready_table_x;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:120:9
		addr_table_n = addr_table;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:121:9
		dequeue_val_n = dequeue_val_r;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:122:9
		dequeue_id_n = dequeue_id_r;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:124:9
		if (dequeue_fire) begin
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:125:13
			dequeue_val_n = dequeue_val_x;
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:126:13
			dequeue_id_n = dequeue_id_x;
		end
		if (allocate_fire) begin
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:130:13
			valid_table_n[allocate_id] = 1;
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:131:13
			ready_table_n[allocate_id] = 0;
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:132:13
			addr_table_n[allocate_id * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)] = allocate_addr;
		end
		if (fill_valid) begin
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:136:13
			dequeue_val_n = 1;
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:137:13
			dequeue_id_n = fill_id;
		end
		if (release_valid)
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:141:13
			valid_table_n[release_id] = 0;
	end
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:145:5
	always @(posedge clk) begin
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:146:9
		if (reset) begin
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:147:13
			valid_table <= 0;
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:148:13
			allocate_rdy_r <= 0;
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:149:13
			dequeue_val_r <= 0;
		end
		else begin
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:151:13
			valid_table <= valid_table_n;
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:152:13
			allocate_rdy_r <= allocate_rdy_n;
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:153:13
			dequeue_val_r <= dequeue_val_n;
		end
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:155:9
		ready_table <= ready_table_n;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:156:9
		addr_table <= addr_table_n;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:157:9
		dequeue_id_r <= dequeue_id_n;
		// Trace: ../../rtl/cache/VX_miss_resrv.sv:158:9
		allocate_id_r <= allocate_id_n;
		if (!allocate_fire || !valid_table[allocate_id_r])
			;
		if (!release_valid || valid_table[release_id])
			;
	end
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:170:5
	VX_dp_ram #(
		.DATAW((((CORE_TAG_WIDTH + 1) + (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) + ($clog2(CACHE_LINE_SIZE / WORD_SIZE) > 0 ? $clog2(CACHE_LINE_SIZE / WORD_SIZE) : 1)) * NUM_PORTS),
		.SIZE(MSHR_SIZE),
		.LUTRAM(1)
	) entries(
		.clk(clk),
		.waddr(allocate_id_r),
		.raddr(dequeue_id_r),
		.wren(allocate_valid),
		.wdata(allocate_data),
		.rdata(dequeue_data)
	);
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:183:5
	assign fill_addr = addr_table[fill_id * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)];
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:185:5
	assign allocate_ready = allocate_rdy_r;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:186:5
	assign allocate_id = allocate_id_r;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:188:5
	assign dequeue_valid = dequeue_val_r;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:189:5
	assign dequeue_id = dequeue_id_r;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:190:5
	assign dequeue_addr = addr_table[dequeue_id_r * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))+:(32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)];
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:192:5
	wire [MSHR_SIZE - 1:0] lookup_entries;
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:193:5
	generate
		for (i = 0; i < MSHR_SIZE; i = i + 1) begin : genblk2
			// Trace: ../../rtl/cache/VX_miss_resrv.sv:194:9
			assign lookup_entries[i] = i != lookup_id;
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_miss_resrv.sv:196:5
	assign lookup_match = |((lookup_entries & valid_table) & addr_matches);
endmodule
module VX_nc_bypass (
	clk,
	reset,
	core_req_valid_in,
	core_req_rw_in,
	core_req_addr_in,
	core_req_byteen_in,
	core_req_data_in,
	core_req_tag_in,
	core_req_ready_in,
	core_req_valid_out,
	core_req_rw_out,
	core_req_addr_out,
	core_req_byteen_out,
	core_req_data_out,
	core_req_tag_out,
	core_req_ready_out,
	core_rsp_valid_in,
	core_rsp_tmask_in,
	core_rsp_data_in,
	core_rsp_tag_in,
	core_rsp_ready_in,
	core_rsp_valid_out,
	core_rsp_tmask_out,
	core_rsp_data_out,
	core_rsp_tag_out,
	core_rsp_ready_out,
	mem_req_valid_in,
	mem_req_rw_in,
	mem_req_addr_in,
	mem_req_pmask_in,
	mem_req_byteen_in,
	mem_req_wsel_in,
	mem_req_data_in,
	mem_req_tag_in,
	mem_req_ready_in,
	mem_req_valid_out,
	mem_req_rw_out,
	mem_req_addr_out,
	mem_req_pmask_out,
	mem_req_byteen_out,
	mem_req_wsel_out,
	mem_req_data_out,
	mem_req_tag_out,
	mem_req_ready_out,
	mem_rsp_valid_in,
	mem_rsp_data_in,
	mem_rsp_tag_in,
	mem_rsp_ready_in,
	mem_rsp_valid_out,
	mem_rsp_data_out,
	mem_rsp_tag_out,
	mem_rsp_ready_out
);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:4:15
	parameter NUM_PORTS = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:5:15
	parameter NUM_REQS = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:6:15
	parameter NUM_RSP_TAGS = 0;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:7:15
	parameter NC_TAG_BIT = 0;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:9:15
	parameter CORE_ADDR_WIDTH = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:10:15
	parameter CORE_DATA_SIZE = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:11:15
	parameter CORE_TAG_IN_WIDTH = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:13:15
	parameter MEM_ADDR_WIDTH = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:14:15
	parameter MEM_DATA_SIZE = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:15:15
	parameter MEM_TAG_IN_WIDTH = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:16:15
	parameter MEM_TAG_OUT_WIDTH = 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:18:15
	parameter CORE_DATA_WIDTH = CORE_DATA_SIZE * 8;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:19:15
	parameter MEM_DATA_WIDTH = MEM_DATA_SIZE * 8;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:20:15
	parameter CORE_TAG_OUT_WIDTH = CORE_TAG_IN_WIDTH - 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:21:15
	parameter MEM_SELECT_BITS = ($clog2(MEM_DATA_SIZE / CORE_DATA_SIZE) > 0 ? $clog2(MEM_DATA_SIZE / CORE_DATA_SIZE) : 1);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:23:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:24:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:27:5
	input wire [NUM_REQS - 1:0] core_req_valid_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:28:5
	input wire [NUM_REQS - 1:0] core_req_rw_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:29:5
	input wire [(NUM_REQS * CORE_ADDR_WIDTH) - 1:0] core_req_addr_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:30:5
	input wire [(NUM_REQS * CORE_DATA_SIZE) - 1:0] core_req_byteen_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:31:5
	input wire [(NUM_REQS * CORE_DATA_WIDTH) - 1:0] core_req_data_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:32:5
	input wire [(NUM_REQS * CORE_TAG_IN_WIDTH) - 1:0] core_req_tag_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:33:5
	output wire [NUM_REQS - 1:0] core_req_ready_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:36:5
	output wire [NUM_REQS - 1:0] core_req_valid_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:37:5
	output wire [NUM_REQS - 1:0] core_req_rw_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:38:5
	output wire [(NUM_REQS * CORE_ADDR_WIDTH) - 1:0] core_req_addr_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:39:5
	output wire [(NUM_REQS * CORE_DATA_SIZE) - 1:0] core_req_byteen_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:40:5
	output wire [(NUM_REQS * CORE_DATA_WIDTH) - 1:0] core_req_data_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:41:5
	output wire [(NUM_REQS * CORE_TAG_OUT_WIDTH) - 1:0] core_req_tag_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:42:5
	input wire [NUM_REQS - 1:0] core_req_ready_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:45:5
	input wire [NUM_RSP_TAGS - 1:0] core_rsp_valid_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:46:5
	input wire [NUM_REQS - 1:0] core_rsp_tmask_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:47:5
	input wire [(NUM_REQS * CORE_DATA_WIDTH) - 1:0] core_rsp_data_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:48:5
	input wire [(NUM_RSP_TAGS * CORE_TAG_OUT_WIDTH) - 1:0] core_rsp_tag_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:49:5
	output wire [NUM_RSP_TAGS - 1:0] core_rsp_ready_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:52:5
	output wire [NUM_RSP_TAGS - 1:0] core_rsp_valid_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:53:5
	output wire [NUM_REQS - 1:0] core_rsp_tmask_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:54:5
	output wire [(NUM_REQS * CORE_DATA_WIDTH) - 1:0] core_rsp_data_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:55:5
	output wire [(NUM_RSP_TAGS * CORE_TAG_IN_WIDTH) - 1:0] core_rsp_tag_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:56:5
	input wire [NUM_RSP_TAGS - 1:0] core_rsp_ready_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:59:5
	input wire mem_req_valid_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:60:5
	input wire mem_req_rw_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:61:5
	input wire [MEM_ADDR_WIDTH - 1:0] mem_req_addr_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:62:5
	input wire [NUM_PORTS - 1:0] mem_req_pmask_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:63:5
	input wire [(NUM_PORTS * CORE_DATA_SIZE) - 1:0] mem_req_byteen_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:64:5
	input wire [(NUM_PORTS * MEM_SELECT_BITS) - 1:0] mem_req_wsel_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:65:5
	input wire [(NUM_PORTS * CORE_DATA_WIDTH) - 1:0] mem_req_data_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:66:5
	input wire [MEM_TAG_IN_WIDTH - 1:0] mem_req_tag_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:67:5
	output wire mem_req_ready_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:70:5
	output wire mem_req_valid_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:71:5
	output wire mem_req_rw_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:72:5
	output wire [MEM_ADDR_WIDTH - 1:0] mem_req_addr_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:73:5
	output wire [NUM_PORTS - 1:0] mem_req_pmask_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:74:5
	output wire [(NUM_PORTS * CORE_DATA_SIZE) - 1:0] mem_req_byteen_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:75:5
	output wire [(NUM_PORTS * MEM_SELECT_BITS) - 1:0] mem_req_wsel_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:76:5
	output wire [(NUM_PORTS * CORE_DATA_WIDTH) - 1:0] mem_req_data_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:77:5
	output wire [MEM_TAG_OUT_WIDTH - 1:0] mem_req_tag_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:78:5
	input wire mem_req_ready_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:81:5
	input wire mem_rsp_valid_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:82:5
	input wire [MEM_DATA_WIDTH - 1:0] mem_rsp_data_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:83:5
	input wire [MEM_TAG_OUT_WIDTH - 1:0] mem_rsp_tag_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:84:5
	output wire mem_rsp_ready_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:87:5
	output wire mem_rsp_valid_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:88:5
	output wire [MEM_DATA_WIDTH - 1:0] mem_rsp_data_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:89:5
	output wire [MEM_TAG_IN_WIDTH - 1:0] mem_rsp_tag_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:90:5
	input wire mem_rsp_ready_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:97:5
	localparam CORE_REQ_TIDW = $clog2(NUM_REQS);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:98:5
	localparam MUX_DATAW = (((CORE_TAG_IN_WIDTH + CORE_DATA_WIDTH) + CORE_DATA_SIZE) + CORE_ADDR_WIDTH) + 1;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:100:5
	localparam CORE_LDATAW = $clog2(CORE_DATA_WIDTH);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:101:5
	localparam MEM_LDATAW = $clog2(MEM_DATA_WIDTH);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:102:5
	localparam D = MEM_LDATAW - CORE_LDATAW;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:106:5
	wire [NUM_REQS - 1:0] core_req_valid_in_nc;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:107:5
	wire [NUM_REQS - 1:0] core_req_nc_tids;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:108:5
	wire [(CORE_REQ_TIDW > 0 ? CORE_REQ_TIDW : 1) - 1:0] core_req_nc_tid;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:109:5
	wire [NUM_REQS - 1:0] core_req_nc_sel;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:110:5
	wire core_req_nc_valid;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:112:5
	genvar i;
	generate
		for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:113:9
			assign core_req_nc_tids[i] = core_req_tag_in[(i * CORE_TAG_IN_WIDTH) + NC_TAG_BIT];
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:116:5
	assign core_req_valid_in_nc = core_req_valid_in & core_req_nc_tids;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:118:5
	VX_priority_encoder #(.N(NUM_REQS)) core_req_sel(
		.data_in(core_req_valid_in_nc),
		.index(core_req_nc_tid),
		.onehot(core_req_nc_sel),
		.valid_out(core_req_nc_valid)
	);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:127:5
	assign core_req_valid_out = core_req_valid_in & ~core_req_nc_tids;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:128:5
	assign core_req_rw_out = core_req_rw_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:129:5
	assign core_req_addr_out = core_req_addr_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:130:5
	assign core_req_byteen_out = core_req_byteen_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:131:5
	assign core_req_data_out = core_req_data_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:133:5
	generate
		for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk2
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:134:9
			VX_bits_remove #(
				.N(CORE_TAG_IN_WIDTH),
				.S(1),
				.POS(NC_TAG_BIT)
			) core_req_tag_remove(
				.data_in(core_req_tag_in[i * CORE_TAG_IN_WIDTH+:CORE_TAG_IN_WIDTH]),
				.data_out(core_req_tag_out[i * CORE_TAG_OUT_WIDTH+:CORE_TAG_OUT_WIDTH])
			);
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:144:5
	generate
		if (NUM_REQS > 1) begin : genblk3
			genvar i;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:146:13
				assign core_req_ready_in[i] = (core_req_valid_in_nc[i] ? (~mem_req_valid_in && mem_req_ready_out) && core_req_nc_sel[i] : core_req_ready_out[i]);
			end
		end
		else begin : genblk3
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:150:9
			assign core_req_ready_in = (core_req_valid_in_nc ? ~mem_req_valid_in && mem_req_ready_out : core_req_ready_out);
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:155:5
	assign mem_req_valid_out = mem_req_valid_in || core_req_nc_valid;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:156:5
	assign mem_req_ready_in = mem_req_ready_out;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:158:5
	wire [MEM_TAG_IN_WIDTH + 0:0] mem_req_tag_in_c;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:160:5
	localparam sv2v_uu_mem_req_tag_insert_S = 1;
	// removed localparam type sv2v_uu_mem_req_tag_insert_sel_in
	localparam [0:0] sv2v_uu_mem_req_tag_insert_ext_sel_in_0 = 1'sb0;
	VX_bits_insert #(
		.N(MEM_TAG_IN_WIDTH),
		.S(1),
		.POS(NC_TAG_BIT)
	) mem_req_tag_insert(
		.data_in(mem_req_tag_in),
		.sel_in(sv2v_uu_mem_req_tag_insert_ext_sel_in_0),
		.data_out(mem_req_tag_in_c)
	);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:170:5
	wire [CORE_TAG_IN_WIDTH - 1:0] core_req_tag_in_sel;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:171:5
	wire [CORE_DATA_WIDTH - 1:0] core_req_data_in_sel;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:172:5
	wire [CORE_DATA_SIZE - 1:0] core_req_byteen_in_sel;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:173:5
	wire [CORE_ADDR_WIDTH - 1:0] core_req_addr_in_sel;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:174:5
	wire core_req_rw_in_sel;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:176:5
	generate
		if (NUM_REQS > 1) begin : genblk4
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:177:9
			wire [(NUM_REQS * MUX_DATAW) - 1:0] core_req_nc_mux_in;
			genvar i;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:179:13
				assign core_req_nc_mux_in[i * MUX_DATAW+:MUX_DATAW] = {core_req_tag_in[i * CORE_TAG_IN_WIDTH+:CORE_TAG_IN_WIDTH], core_req_data_in[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH], core_req_byteen_in[i * CORE_DATA_SIZE+:CORE_DATA_SIZE], core_req_addr_in[i * CORE_ADDR_WIDTH+:CORE_ADDR_WIDTH], core_req_rw_in[i]};
			end
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:182:9
			assign {core_req_tag_in_sel, core_req_data_in_sel, core_req_byteen_in_sel, core_req_addr_in_sel, core_req_rw_in_sel} = core_req_nc_mux_in[core_req_nc_tid * MUX_DATAW+:MUX_DATAW];
		end
		else begin : genblk4
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:184:9
			assign core_req_tag_in_sel = core_req_tag_in;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:185:9
			assign core_req_data_in_sel = core_req_data_in;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:186:9
			assign core_req_byteen_in_sel = core_req_byteen_in;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:187:9
			assign core_req_addr_in_sel = core_req_addr_in;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:188:9
			assign core_req_rw_in_sel = core_req_rw_in;
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:191:5
	assign mem_req_rw_out = (mem_req_valid_in ? mem_req_rw_in : core_req_rw_in_sel);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:192:5
	assign mem_req_addr_out = (mem_req_valid_in ? mem_req_addr_in : core_req_addr_in_sel[D+:MEM_ADDR_WIDTH]);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:194:5
	function automatic [MEM_TAG_OUT_WIDTH - 1:0] sv2v_cast_CEA83;
		input reg [MEM_TAG_OUT_WIDTH - 1:0] inp;
		sv2v_cast_CEA83 = inp;
	endfunction
	function automatic [NUM_PORTS - 1:0] sv2v_cast_1AD22;
		input reg [NUM_PORTS - 1:0] inp;
		sv2v_cast_1AD22 = inp;
	endfunction
	generate
		if (D != 0) begin : genblk5
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:195:9
			reg [(NUM_PORTS * CORE_DATA_SIZE) - 1:0] mem_req_byteen_in_r;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:196:9
			reg [(NUM_PORTS * MEM_SELECT_BITS) - 1:0] mem_req_wsel_in_r;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:197:9
			reg [(NUM_PORTS * CORE_DATA_WIDTH) - 1:0] mem_req_data_in_r;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:199:9
			wire [D - 1:0] req_addr_idx = core_req_addr_in_sel[D - 1:0];
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:201:9
			always @(*) begin
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:202:13
				mem_req_byteen_in_r = 0;
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:203:13
				mem_req_byteen_in_r[0+:CORE_DATA_SIZE] = core_req_byteen_in_sel;
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:205:13
				mem_req_wsel_in_r = 1'sbx;
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:206:13
				mem_req_wsel_in_r[0+:MEM_SELECT_BITS] = req_addr_idx;
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:208:13
				mem_req_data_in_r = 1'sbx;
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:209:13
				mem_req_data_in_r[0+:CORE_DATA_WIDTH] = core_req_data_in_sel;
			end
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:212:9
			assign mem_req_pmask_out = (mem_req_valid_in ? mem_req_pmask_in : sv2v_cast_1AD22(1'b1));
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:213:9
			assign mem_req_byteen_out = (mem_req_valid_in ? mem_req_byteen_in : mem_req_byteen_in_r);
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:214:9
			assign mem_req_wsel_out = (mem_req_valid_in ? mem_req_wsel_in : mem_req_wsel_in_r);
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:215:9
			assign mem_req_data_out = (mem_req_valid_in ? mem_req_data_in : mem_req_data_in_r);
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:216:9
			assign mem_req_tag_out = (mem_req_valid_in ? sv2v_cast_CEA83(mem_req_tag_in_c) : sv2v_cast_CEA83({core_req_nc_tid, req_addr_idx, core_req_tag_in_sel}));
		end
		else begin : genblk5
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:220:9
			assign mem_req_pmask_out = 0;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:221:9
			assign mem_req_byteen_out = (mem_req_valid_in ? mem_req_byteen_in : core_req_byteen_in_sel);
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:222:9
			assign mem_req_data_out = (mem_req_valid_in ? mem_req_data_in : core_req_data_in_sel);
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:223:9
			assign mem_req_wsel_out = 0;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:224:9
			assign mem_req_tag_out = (mem_req_valid_in ? sv2v_cast_CEA83(mem_req_tag_in_c) : sv2v_cast_CEA83({core_req_nc_tid, core_req_tag_in_sel}));
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:229:5
	wire [(NUM_RSP_TAGS * CORE_TAG_IN_WIDTH) - 1:0] core_rsp_tag_out_c;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:231:5
	wire is_mem_rsp_nc = mem_rsp_valid_in && mem_rsp_tag_in[NC_TAG_BIT];
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:233:5
	generate
		for (i = 0; i < NUM_RSP_TAGS; i = i + 1) begin : genblk6
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:234:9
			localparam sv2v_uu_core_rsp_tag_insert_S = 1;
			// removed localparam type sv2v_uu_core_rsp_tag_insert_sel_in
			localparam [0:0] sv2v_uu_core_rsp_tag_insert_ext_sel_in_0 = 1'sb0;
			VX_bits_insert #(
				.N(CORE_TAG_OUT_WIDTH),
				.S(1),
				.POS(NC_TAG_BIT)
			) core_rsp_tag_insert(
				.data_in(core_rsp_tag_in[i * CORE_TAG_OUT_WIDTH+:CORE_TAG_OUT_WIDTH]),
				.sel_in(sv2v_uu_core_rsp_tag_insert_ext_sel_in_0),
				.data_out(core_rsp_tag_out_c[i * CORE_TAG_IN_WIDTH+:CORE_TAG_IN_WIDTH])
			);
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:245:5
	generate
		if (NUM_RSP_TAGS > 1) begin : genblk7
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:246:9
			wire [CORE_REQ_TIDW - 1:0] rsp_tid = mem_rsp_tag_in[CORE_TAG_IN_WIDTH + D+:CORE_REQ_TIDW];
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:247:9
			reg [NUM_REQS - 1:0] rsp_nc_valid_r;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:248:9
			always @(*) begin
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:249:13
				rsp_nc_valid_r = 0;
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:250:13
				rsp_nc_valid_r[rsp_tid] = is_mem_rsp_nc;
			end
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:253:9
			assign core_rsp_valid_out = core_rsp_valid_in | rsp_nc_valid_r;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:254:9
			assign core_rsp_tmask_out = core_rsp_tmask_in;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:255:9
			assign core_rsp_ready_in = core_rsp_ready_out;
			if (D != 0) begin : genblk1
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:258:13
				wire [D - 1:0] rsp_addr_idx = mem_rsp_tag_in[CORE_TAG_IN_WIDTH+:D];
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_nc_bypass.sv:260:17
					assign core_rsp_data_out[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH] = (core_rsp_valid_in[i] ? core_rsp_data_in[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH] : mem_rsp_data_in[rsp_addr_idx * CORE_DATA_WIDTH+:CORE_DATA_WIDTH]);
				end
			end
			else begin : genblk1
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_nc_bypass.sv:265:17
					assign core_rsp_data_out[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH] = (core_rsp_valid_in[i] ? core_rsp_data_in[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH] : mem_rsp_data_in);
				end
			end
			genvar i;
			for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk2
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:270:13
				assign core_rsp_tag_out[i * CORE_TAG_IN_WIDTH+:CORE_TAG_IN_WIDTH] = (core_rsp_valid_in[i] ? core_rsp_tag_out_c[i * CORE_TAG_IN_WIDTH+:CORE_TAG_IN_WIDTH] : mem_rsp_tag_in[CORE_TAG_IN_WIDTH - 1:0]);
			end
		end
		else begin : genblk7
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:273:9
			assign core_rsp_valid_out = core_rsp_valid_in || is_mem_rsp_nc;
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:274:9
			assign core_rsp_tag_out = (core_rsp_valid_in ? core_rsp_tag_out_c : mem_rsp_tag_in[CORE_TAG_IN_WIDTH - 1:0]);
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:275:9
			assign core_rsp_ready_in = core_rsp_ready_out;
			if (NUM_REQS > 1) begin : genblk1
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:278:13
				wire [CORE_REQ_TIDW - 1:0] rsp_tid = mem_rsp_tag_in[CORE_TAG_IN_WIDTH + D+:CORE_REQ_TIDW];
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:279:13
				reg [NUM_REQS - 1:0] core_rsp_tmask_in_r;
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:280:13
				always @(*) begin
					// Trace: ../../rtl/cache/VX_nc_bypass.sv:281:17
					core_rsp_tmask_in_r = 0;
					// Trace: ../../rtl/cache/VX_nc_bypass.sv:282:17
					core_rsp_tmask_in_r[rsp_tid] = 1;
				end
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:284:13
				assign core_rsp_tmask_out = (core_rsp_valid_in ? core_rsp_tmask_in : core_rsp_tmask_in_r);
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:286:13
				assign core_rsp_tmask_out = core_rsp_tmask_in || is_mem_rsp_nc;
			end
			if (D != 0) begin : genblk2
				// Trace: ../../rtl/cache/VX_nc_bypass.sv:290:13
				wire [D - 1:0] rsp_addr_idx = mem_rsp_tag_in[CORE_TAG_IN_WIDTH+:D];
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_nc_bypass.sv:292:17
					assign core_rsp_data_out[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH] = (core_rsp_valid_in ? core_rsp_data_in[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH] : mem_rsp_data_in[rsp_addr_idx * CORE_DATA_WIDTH+:CORE_DATA_WIDTH]);
				end
			end
			else begin : genblk2
				genvar i;
				for (i = 0; i < NUM_REQS; i = i + 1) begin : genblk1
					// Trace: ../../rtl/cache/VX_nc_bypass.sv:297:17
					assign core_rsp_data_out[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH] = (core_rsp_valid_in ? core_rsp_data_in[i * CORE_DATA_WIDTH+:CORE_DATA_WIDTH] : mem_rsp_data_in);
				end
			end
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:304:5
	assign mem_rsp_valid_out = mem_rsp_valid_in && ~mem_rsp_tag_in[NC_TAG_BIT];
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:305:5
	assign mem_rsp_data_out = mem_rsp_data_in;
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:307:5
	VX_bits_remove #(
		.N(MEM_TAG_IN_WIDTH + 1),
		.S(1),
		.POS(NC_TAG_BIT)
	) mem_rsp_tag_remove(
		.data_in(mem_rsp_tag_in[MEM_TAG_IN_WIDTH + 0:0]),
		.data_out(mem_rsp_tag_out)
	);
	// Trace: ../../rtl/cache/VX_nc_bypass.sv:316:5
	generate
		if (NUM_RSP_TAGS > 1) begin : genblk8
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:317:9
			wire [CORE_REQ_TIDW - 1:0] rsp_tid = mem_rsp_tag_in[CORE_TAG_IN_WIDTH + D+:CORE_REQ_TIDW];
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:318:9
			assign mem_rsp_ready_in = (is_mem_rsp_nc ? ~core_rsp_valid_in[rsp_tid] && core_rsp_ready_out[rsp_tid] : mem_rsp_ready_out);
		end
		else begin : genblk8
			// Trace: ../../rtl/cache/VX_nc_bypass.sv:320:9
			assign mem_rsp_ready_in = (is_mem_rsp_nc ? ~core_rsp_valid_in && core_rsp_ready_out : mem_rsp_ready_out);
		end
	endgenerate
endmodule
module VX_shared_mem (
	clk,
	reset,
	core_req_valid,
	core_req_rw,
	core_req_addr,
	core_req_byteen,
	core_req_data,
	core_req_tag,
	core_req_ready,
	core_rsp_valid,
	core_rsp_tmask,
	core_rsp_data,
	core_rsp_tag,
	core_rsp_ready
);
	// Trace: ../../rtl/cache/VX_shared_mem.sv:4:15
	parameter CACHE_ID = 0;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:7:15
	parameter CACHE_SIZE = 16384;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:9:15
	parameter NUM_BANKS = 2;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:11:15
	parameter WORD_SIZE = 4;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:13:15
	parameter NUM_REQS = 4;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:16:15
	parameter CREQ_SIZE = 2;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:18:15
	parameter CRSQ_SIZE = 2;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:21:15
	parameter CORE_TAG_ID_BITS = 8;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:24:15
	parameter CORE_TAG_WIDTH = 2 + CORE_TAG_ID_BITS;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:27:15
	parameter BANK_ADDR_OFFSET = 8;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:29:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:30:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:38:5
	input wire [NUM_REQS - 1:0] core_req_valid;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:39:5
	input wire [NUM_REQS - 1:0] core_req_rw;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:40:5
	input wire [(NUM_REQS * (32 - $clog2(WORD_SIZE))) - 1:0] core_req_addr;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:41:5
	input wire [(NUM_REQS * WORD_SIZE) - 1:0] core_req_byteen;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:42:5
	input wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_req_data;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:43:5
	input wire [(NUM_REQS * CORE_TAG_WIDTH) - 1:0] core_req_tag;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:44:5
	output wire [NUM_REQS - 1:0] core_req_ready;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:47:5
	output wire core_rsp_valid;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:48:5
	output wire [NUM_REQS - 1:0] core_rsp_tmask;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:49:5
	output wire [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_rsp_data;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:50:5
	output wire [CORE_TAG_WIDTH - 1:0] core_rsp_tag;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:51:5
	input wire core_rsp_ready;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:58:5
	localparam CACHE_LINE_SIZE = WORD_SIZE;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:60:5
	wire [NUM_BANKS - 1:0] per_bank_core_req_valid_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:61:5
	wire [NUM_BANKS - 1:0] per_bank_core_req_rw_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:62:5
	wire [(NUM_BANKS * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] per_bank_core_req_addr_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:63:5
	wire [(NUM_BANKS * WORD_SIZE) - 1:0] per_bank_core_req_byteen_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:64:5
	wire [(NUM_BANKS * (8 * WORD_SIZE)) - 1:0] per_bank_core_req_data_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:65:5
	wire [(NUM_BANKS * CORE_TAG_WIDTH) - 1:0] per_bank_core_req_tag_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:66:5
	wire [(NUM_BANKS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] per_bank_core_req_tid_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:67:5
	wire [NUM_BANKS - 1:0] per_bank_core_req_ready_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:69:5
	VX_core_req_bank_sel #(
		.CACHE_ID(CACHE_ID),
		.CACHE_LINE_SIZE(WORD_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_PORTS(1),
		.WORD_SIZE(WORD_SIZE),
		.NUM_REQS(NUM_REQS),
		.CORE_TAG_WIDTH(CORE_TAG_WIDTH),
		.BANK_ADDR_OFFSET(BANK_ADDR_OFFSET)
	) core_req_bank_sel(
		.clk(clk),
		.reset(reset),
		.core_req_valid(core_req_valid),
		.core_req_rw(core_req_rw),
		.core_req_addr(core_req_addr),
		.core_req_byteen(core_req_byteen),
		.core_req_data(core_req_data),
		.core_req_tag(core_req_tag),
		.core_req_ready(core_req_ready),
		.per_bank_core_req_valid(per_bank_core_req_valid_unqual),
		.per_bank_core_req_tid(per_bank_core_req_tid_unqual),
		.per_bank_core_req_rw(per_bank_core_req_rw_unqual),
		.per_bank_core_req_addr(per_bank_core_req_addr_unqual),
		.per_bank_core_req_byteen(per_bank_core_req_byteen_unqual),
		.per_bank_core_req_tag(per_bank_core_req_tag_unqual),
		.per_bank_core_req_data(per_bank_core_req_data_unqual),
		.per_bank_core_req_ready(per_bank_core_req_ready_unqual)
	);
	// Trace: ../../rtl/cache/VX_shared_mem.sv:103:5
	wire [NUM_BANKS - 1:0] per_bank_core_req_valid;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:104:5
	wire [NUM_BANKS - 1:0] per_bank_core_req_rw;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:105:5
	wire [(NUM_BANKS * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) - 1:0] per_bank_core_req_addr;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:106:5
	wire [(NUM_BANKS * WORD_SIZE) - 1:0] per_bank_core_req_byteen;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:107:5
	wire [(NUM_BANKS * (8 * WORD_SIZE)) - 1:0] per_bank_core_req_data;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:108:5
	wire [(NUM_BANKS * CORE_TAG_WIDTH) - 1:0] per_bank_core_req_tag;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:109:5
	wire [(NUM_BANKS * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)) - 1:0] per_bank_core_req_tid;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:111:5
	wire creq_out_valid;
	wire creq_out_ready;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:112:5
	wire creq_in_valid;
	wire creq_in_ready;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:114:5
	wire creq_in_fire = creq_in_valid && creq_in_ready;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:117:5
	wire creq_out_fire = creq_out_valid && creq_out_ready;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:120:5
	assign creq_in_valid = |core_req_valid;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:121:5
	assign per_bank_core_req_ready_unqual = {NUM_BANKS {creq_in_ready}};
	// Trace: ../../rtl/cache/VX_shared_mem.sv:123:5
	wire [NUM_BANKS - 1:0] core_req_read_mask;
	wire [NUM_BANKS - 1:0] core_req_read_mask_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:124:5
	wire core_req_writeonly;
	wire core_req_writeonly_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:126:5
	assign core_req_read_mask_unqual = per_bank_core_req_valid_unqual & ~per_bank_core_req_rw_unqual;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:127:5
	assign core_req_writeonly_unqual = ~(|core_req_read_mask_unqual);
	// Trace: ../../rtl/cache/VX_shared_mem.sv:129:5
	VX_elastic_buffer #(
		.DATAW(((NUM_BANKS * (((((2 + ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) + WORD_SIZE) + (8 * WORD_SIZE)) + CORE_TAG_WIDTH) + (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1))) + NUM_BANKS) + 1),
		.SIZE(CREQ_SIZE),
		.OUT_REG(1)
	) core_req_queue(
		.clk(clk),
		.reset(reset),
		.ready_in(creq_in_ready),
		.valid_in(creq_in_valid),
		.data_in({per_bank_core_req_valid_unqual, per_bank_core_req_rw_unqual, per_bank_core_req_addr_unqual, per_bank_core_req_byteen_unqual, per_bank_core_req_data_unqual, per_bank_core_req_tag_unqual, per_bank_core_req_tid_unqual, core_req_read_mask_unqual, core_req_writeonly_unqual}),
		.data_out({per_bank_core_req_valid, per_bank_core_req_rw, per_bank_core_req_addr, per_bank_core_req_byteen, per_bank_core_req_data, per_bank_core_req_tag, per_bank_core_req_tid, core_req_read_mask, core_req_writeonly}),
		.ready_out(creq_out_ready),
		.valid_out(creq_out_valid)
	);
	// Trace: ../../rtl/cache/VX_shared_mem.sv:160:5
	wire crsq_in_valid;
	wire crsq_in_ready;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:161:5
	wire crsq_last_read;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:163:5
	assign creq_out_ready = core_req_writeonly || (crsq_in_ready && crsq_last_read);
	// Trace: ../../rtl/cache/VX_shared_mem.sv:166:5
	wire [(NUM_BANKS * (8 * WORD_SIZE)) - 1:0] per_bank_core_rsp_data;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:168:5
	genvar i;
	generate
		for (i = 0; i < NUM_BANKS; i = i + 1) begin : genblk1
			// Trace: ../../rtl/cache/VX_shared_mem.sv:170:9
			wire [WORD_SIZE - 1:0] wren = per_bank_core_req_byteen[i * WORD_SIZE+:WORD_SIZE] & {WORD_SIZE {per_bank_core_req_valid[i] && per_bank_core_req_rw[i]}};
			// Trace: ../../rtl/cache/VX_shared_mem.sv:174:9
			wire [$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0] addr = per_bank_core_req_addr[(i * ((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS))) + ($clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1)-:$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE)];
			// Trace: ../../rtl/cache/VX_shared_mem.sv:176:9
			VX_sp_ram #(
				.DATAW(8 * WORD_SIZE),
				.SIZE((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE),
				.BYTEENW(WORD_SIZE),
				.NO_RWCHECK(1)
			) data_store(
				.clk(clk),
				.addr(addr),
				.wren(wren),
				.wdata(per_bank_core_req_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE]),
				.rdata(per_bank_core_rsp_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE])
			);
		end
	endgenerate
	// Trace: ../../rtl/cache/VX_shared_mem.sv:194:5
	reg [NUM_REQS - 1:0] core_rsp_valids_in;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:195:5
	reg [(NUM_REQS * (8 * WORD_SIZE)) - 1:0] core_rsp_data_in;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:196:5
	wire [CORE_TAG_WIDTH - 1:0] core_rsp_tag_in;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:197:5
	reg [NUM_BANKS - 1:0] bank_rsp_sel_r;
	reg [NUM_BANKS - 1:0] bank_rsp_sel_n;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:199:5
	wire crsq_in_fire = crsq_in_valid && crsq_in_ready;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:201:5
	assign crsq_last_read = bank_rsp_sel_n == core_req_read_mask;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:203:5
	always @(posedge clk)
		// Trace: ../../rtl/cache/VX_shared_mem.sv:204:9
		if (reset)
			// Trace: ../../rtl/cache/VX_shared_mem.sv:205:13
			bank_rsp_sel_r <= 0;
		else
			// Trace: ../../rtl/cache/VX_shared_mem.sv:207:13
			if (crsq_in_fire)
				// Trace: ../../rtl/cache/VX_shared_mem.sv:208:17
				if (crsq_last_read)
					// Trace: ../../rtl/cache/VX_shared_mem.sv:209:21
					bank_rsp_sel_r <= 0;
				else
					// Trace: ../../rtl/cache/VX_shared_mem.sv:211:21
					bank_rsp_sel_r <= bank_rsp_sel_n;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:217:5
	VX_find_first #(
		.N(NUM_BANKS),
		.DATAW(CORE_TAG_WIDTH)
	) find_first(
		.valid_i(core_req_read_mask & ~bank_rsp_sel_r),
		.data_i(per_bank_core_req_tag),
		.data_o(core_rsp_tag_in)
	);
	// Trace: ../../rtl/cache/VX_shared_mem.sv:227:5
	always @(*) begin
		// Trace: ../../rtl/cache/VX_shared_mem.sv:228:9
		core_rsp_valids_in = 0;
		// Trace: ../../rtl/cache/VX_shared_mem.sv:229:9
		core_rsp_data_in = 1'sbx;
		// Trace: ../../rtl/cache/VX_shared_mem.sv:230:9
		bank_rsp_sel_n = bank_rsp_sel_r;
		// Trace: ../../rtl/cache/VX_shared_mem.sv:231:9
		begin : sv2v_autoblock_1
			// Trace: ../../rtl/cache/VX_shared_mem.sv:231:14
			integer i;
			// Trace: ../../rtl/cache/VX_shared_mem.sv:231:14
			for (i = 0; i < NUM_BANKS; i = i + 1)
				begin
					// Trace: ../../rtl/cache/VX_shared_mem.sv:232:13
					if (core_req_read_mask[i] && (core_rsp_tag_in[CORE_TAG_ID_BITS - 1:0] == per_bank_core_req_tag[(i * CORE_TAG_WIDTH) + (CORE_TAG_ID_BITS - 1)-:CORE_TAG_ID_BITS])) begin
						// Trace: ../../rtl/cache/VX_shared_mem.sv:234:17
						core_rsp_valids_in[per_bank_core_req_tid[i * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)]] = 1;
						// Trace: ../../rtl/cache/VX_shared_mem.sv:235:17
						core_rsp_data_in[per_bank_core_req_tid[i * (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)+:(NUM_REQS > 1 ? $clog2(NUM_REQS) : 1)] * (8 * WORD_SIZE)+:8 * WORD_SIZE] = per_bank_core_rsp_data[i * (8 * WORD_SIZE)+:8 * WORD_SIZE];
						// Trace: ../../rtl/cache/VX_shared_mem.sv:236:17
						bank_rsp_sel_n[i] = 1;
					end
				end
		end
	end
	// Trace: ../../rtl/cache/VX_shared_mem.sv:241:5
	assign crsq_in_valid = creq_out_valid && ~core_req_writeonly;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:243:5
	VX_elastic_buffer #(
		.DATAW((NUM_BANKS * (1 + (8 * WORD_SIZE))) + CORE_TAG_WIDTH),
		.SIZE(CRSQ_SIZE)
	) core_rsp_req(
		.clk(clk),
		.reset(reset),
		.valid_in(crsq_in_valid),
		.data_in({core_rsp_valids_in, core_rsp_data_in, core_rsp_tag_in}),
		.ready_in(crsq_in_ready),
		.valid_out(core_rsp_valid),
		.data_out({core_rsp_tmask, core_rsp_data, core_rsp_tag}),
		.ready_out(core_rsp_ready)
	);
	// Trace: ../../rtl/cache/VX_shared_mem.sv:258:5
	wire [(NUM_BANKS * 44) - 1:0] req_id_st0;
	wire [(NUM_BANKS * 44) - 1:0] req_id_st1;
	// Trace: ../../rtl/cache/VX_shared_mem.sv:261:5
	generate
		for (i = 0; i < NUM_BANKS; i = i + 1) begin : genblk2
			if ((CORE_TAG_WIDTH != CORE_TAG_ID_BITS) && (CORE_TAG_ID_BITS != 0)) begin : genblk1
				// Trace: ../../rtl/cache/VX_shared_mem.sv:263:13
				assign req_id_st0[i * 44+:44] = per_bank_core_req_tag_unqual[(i * CORE_TAG_WIDTH) + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? CORE_TAG_WIDTH - 1 : ((CORE_TAG_WIDTH - 1) + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)) - 1)-:((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)];
				// Trace: ../../rtl/cache/VX_shared_mem.sv:264:13
				assign req_id_st1[i * 44+:44] = per_bank_core_req_tag[(i * CORE_TAG_WIDTH) + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? CORE_TAG_WIDTH - 1 : ((CORE_TAG_WIDTH - 1) + ((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)) - 1)-:((CORE_TAG_WIDTH - 1) >= (CORE_TAG_WIDTH - 44) ? ((CORE_TAG_WIDTH - 1) - (CORE_TAG_WIDTH - 44)) + 1 : ((CORE_TAG_WIDTH - 44) - (CORE_TAG_WIDTH - 1)) + 1)];
			end
			else begin : genblk1
				// Trace: ../../rtl/cache/VX_shared_mem.sv:266:13
				assign req_id_st0[i * 44+:44] = 0;
				// Trace: ../../rtl/cache/VX_shared_mem.sv:267:13
				assign req_id_st1[i * 44+:44] = 0;
			end
		end
	endgenerate
endmodule
module VX_tag_access (
	clk,
	reset,
	req_id,
	stall,
	lookup,
	addr,
	fill,
	flush,
	tag_match
);
	// Trace: ../../rtl/cache/VX_tag_access.sv:4:15
	parameter CACHE_ID = 0;
	// Trace: ../../rtl/cache/VX_tag_access.sv:5:15
	parameter BANK_ID = 0;
	// Trace: ../../rtl/cache/VX_tag_access.sv:7:15
	parameter CACHE_SIZE = 1;
	// Trace: ../../rtl/cache/VX_tag_access.sv:9:15
	parameter CACHE_LINE_SIZE = 1;
	// Trace: ../../rtl/cache/VX_tag_access.sv:11:15
	parameter NUM_BANKS = 1;
	// Trace: ../../rtl/cache/VX_tag_access.sv:13:15
	parameter WORD_SIZE = 1;
	// Trace: ../../rtl/cache/VX_tag_access.sv:15:15
	parameter BANK_ADDR_OFFSET = 0;
	// Trace: ../../rtl/cache/VX_tag_access.sv:17:5
	input wire clk;
	// Trace: ../../rtl/cache/VX_tag_access.sv:18:5
	input wire reset;
	// Trace: ../../rtl/cache/VX_tag_access.sv:21:5
	input wire [43:0] req_id;
	// Trace: ../../rtl/cache/VX_tag_access.sv:24:5
	input wire stall;
	// Trace: ../../rtl/cache/VX_tag_access.sv:27:5
	input wire lookup;
	// Trace: ../../rtl/cache/VX_tag_access.sv:28:5
	input wire [((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr;
	// Trace: ../../rtl/cache/VX_tag_access.sv:29:5
	input wire fill;
	// Trace: ../../rtl/cache/VX_tag_access.sv:30:5
	input wire flush;
	// Trace: ../../rtl/cache/VX_tag_access.sv:31:5
	output wire tag_match;
	// Trace: ../../rtl/cache/VX_tag_access.sv:39:5
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) - BANK_ADDR_OFFSET) + $clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE)) - 1)) - 1:0] read_tag;
	// Trace: ../../rtl/cache/VX_tag_access.sv:40:5
	wire read_valid;
	// Trace: ../../rtl/cache/VX_tag_access.sv:42:5
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0] line_addr = addr[$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE) - 1:0];
	// Trace: ../../rtl/cache/VX_tag_access.sv:43:5
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) - BANK_ADDR_OFFSET) + $clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE)) - 1)) - 1:0] line_tag = addr[((32 - $clog2(CACHE_LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:$clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE)];
	// Trace: ../../rtl/cache/VX_tag_access.sv:45:5
	VX_sp_ram #(
		.DATAW((((32 - $clog2(WORD_SIZE)) - 1) - ((((((((0 + $clog2(CACHE_LINE_SIZE / WORD_SIZE)) + 0) + BANK_ADDR_OFFSET) + $clog2(NUM_BANKS)) + 0) - BANK_ADDR_OFFSET) + $clog2((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE)) - 1)) + 1),
		.SIZE((CACHE_SIZE / NUM_BANKS) / CACHE_LINE_SIZE),
		.NO_RWCHECK(1)
	) tag_store(
		.clk(clk),
		.addr(line_addr),
		.wren(fill || flush),
		.wdata({!flush, line_tag}),
		.rdata({read_valid, read_tag})
	);
	// Trace: ../../rtl/cache/VX_tag_access.sv:57:5
	assign tag_match = read_valid && (line_tag == read_tag);
endmodule
// Trace: ../../rtl/fp_cores/VX_fpu_define.vh:11:1
// removed ["import fpu_types::*;"]
module VX_fp_class (
	exp_i,
	man_i,
	clss_o
);
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:5:15
	parameter MAN_BITS = 23;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:6:15
	parameter EXP_BITS = 8;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:8:5
	input [EXP_BITS - 1:0] exp_i;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:9:5
	input [MAN_BITS - 1:0] man_i;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:10:5
	// removed localparam type fpu_types_fp_class_t
	output wire [6:0] clss_o;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:12:5
	wire is_normal = (exp_i != {EXP_BITS {1'sb0}}) && (exp_i != {EXP_BITS {1'sb1}});
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:13:5
	wire is_zero = (exp_i == {EXP_BITS {1'sb0}}) && (man_i == {MAN_BITS {1'sb0}});
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:14:5
	wire is_subnormal = (exp_i == {EXP_BITS {1'sb0}}) && (man_i != {MAN_BITS {1'sb0}});
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:15:5
	wire is_inf = (exp_i == {EXP_BITS {1'sb1}}) && (man_i == {MAN_BITS {1'sb0}});
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:16:5
	wire is_nan = (exp_i == {EXP_BITS {1'sb1}}) && (man_i != {MAN_BITS {1'sb0}});
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:17:5
	wire is_signaling = is_nan && ~man_i[MAN_BITS - 1];
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:18:5
	wire is_quiet = is_nan && ~is_signaling;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:20:5
	assign clss_o[6] = is_normal;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:21:5
	assign clss_o[5] = is_zero;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:22:5
	assign clss_o[4] = is_subnormal;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:23:5
	assign clss_o[3] = is_inf;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:24:5
	assign clss_o[2] = is_nan;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:25:5
	assign clss_o[1] = is_quiet;
	// Trace: ../../rtl/fp_cores/VX_fp_class.sv:26:5
	assign clss_o[0] = is_signaling;
endmodule
module VX_fp_cvt (
	clk,
	reset,
	ready_in,
	valid_in,
	tag_in,
	frm,
	is_itof,
	is_signed,
	dataa,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:7:15
	parameter TAGW = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:8:15
	parameter LANES = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:10:5
	input wire clk;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:11:5
	input wire reset;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:13:5
	output wire ready_in;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:14:5
	input wire valid_in;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:16:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:18:5
	input wire [2:0] frm;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:20:5
	input wire is_itof;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:21:5
	input wire is_signed;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:23:5
	input wire [(LANES * 32) - 1:0] dataa;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:24:5
	output wire [(LANES * 32) - 1:0] result;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:26:5
	output wire has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:27:5
	// removed localparam type fpu_types_fflags_t
	output wire [(LANES * 5) - 1:0] fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:29:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:31:5
	input wire ready_out;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:32:5
	output wire valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:36:5
	localparam MAN_BITS = 23;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:37:5
	localparam EXP_BITS = 8;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:38:5
	localparam EXP_BIAS = 127;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:41:5
	localparam MAX_INT_WIDTH = 32;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:44:5
	localparam INT_MAN_WIDTH = MAX_INT_WIDTH;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:47:5
	localparam LZC_RESULT_WIDTH = 5;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:51:5
	localparam INT_EXP_WIDTH = 9;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:54:5
	localparam SHAMT_BITS = 6;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:56:5
	localparam FMT_SHIFT_COMPENSATION = 8;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:57:5
	localparam NUM_FP_STICKY = 40;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:58:5
	localparam NUM_INT_STICKY = 32;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:62:5
	// removed localparam type fpu_types_fp_class_t
	wire [(LANES * 7) - 1:0] fp_clss;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:64:5
	genvar i;
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk1
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:65:9
			VX_fp_class #(
				.EXP_BITS(EXP_BITS),
				.MAN_BITS(MAN_BITS)
			) fp_class(
				.exp_i(dataa[(i * 32) + 30-:8]),
				.man_i(dataa[(i * 32) + 22-:23]),
				.clss_o(fp_clss[i * 7+:7])
			);
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:75:5
	wire [(LANES * 32) - 1:0] encoded_mant;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:76:5
	wire [(LANES * 9) - 1:0] fmt_exponent;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:77:5
	wire [LANES - 1:0] input_sign;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:79:5
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk2
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:81:9
			wire [31:0] int_mantissa;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:82:9
			wire [31:0] fmt_mantissa;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:83:9
			wire fmt_sign = dataa[(i * 32) + 31];
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:84:9
			wire int_sign = dataa[(i * 32) + 31] & is_signed;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:85:9
			assign int_mantissa = (int_sign ? -dataa[i * 32+:32] : dataa[i * 32+:32]);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:86:9
			assign fmt_mantissa = sv2v_cast_32({fp_clss[(i * 7) + 6], dataa[(i * 32) + 22-:23]});
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:87:9
			assign fmt_exponent[i * 9+:9] = {1'b0, dataa[(i * 32) + MAN_BITS+:EXP_BITS]} + {1'b0, fp_clss[(i * 7) + 4]};
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:89:9
			assign encoded_mant[i * 32+:32] = (is_itof ? int_mantissa : fmt_mantissa);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:90:9
			assign input_sign[i] = (is_itof ? int_sign : fmt_sign);
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:96:5
	wire valid_in_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:97:5
	wire [TAGW - 1:0] tag_in_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:98:5
	wire is_itof_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:99:5
	wire unsigned_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:100:5
	wire [2:0] rnd_mode_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:101:5
	wire [(LANES * 7) - 1:0] fp_clss_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:102:5
	wire [LANES - 1:0] input_sign_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:103:5
	wire [(LANES * 9) - 1:0] fmt_exponent_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:104:5
	wire [(LANES * 32) - 1:0] encoded_mant_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:106:5
	wire stall;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:108:5
	VX_pipe_register #(
		.DATAW(((1 + TAGW) + 5) + (LANES * 49)),
		.RESETW(1)
	) pipe_reg0(
		.clk(clk),
		.reset(reset),
		.enable(~stall),
		.data_in({valid_in, tag_in, is_itof, !is_signed, frm, fp_clss, input_sign, fmt_exponent, encoded_mant}),
		.data_out({valid_in_s0, tag_in_s0, is_itof_s0, unsigned_s0, rnd_mode_s0, fp_clss_s0, input_sign_s0, fmt_exponent_s0, encoded_mant_s0})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:121:5
	wire [(LANES * 5) - 1:0] renorm_shamt_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:122:5
	wire [LANES - 1:0] mant_is_zero_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:124:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk3
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:125:9
			wire mant_is_nonzero;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:126:9
			VX_lzc #(
				.N(INT_MAN_WIDTH),
				.MODE(1)
			) lzc(
				.in_i(encoded_mant_s0[i * 32+:32]),
				.cnt_o(renorm_shamt_s0[i * 5+:5]),
				.valid_o(mant_is_nonzero)
			);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:134:9
			assign mant_is_zero_s0[i] = ~mant_is_nonzero;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:137:5
	wire [(LANES * 32) - 1:0] input_mant_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:138:5
	wire [(LANES * 9) - 1:0] input_exp_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:140:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk4
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:143:9
			assign input_mant_s0[i * 32+:32] = encoded_mant_s0[i * 32+:32] << renorm_shamt_s0[i * 5+:5];
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:146:9
			wire [8:0] fp_input_exp = (fmt_exponent_s0[i * 9+:9] + (FMT_SHIFT_COMPENSATION - EXP_BIAS)) - {1'b0, renorm_shamt_s0[i * 5+:5]};
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:147:9
			wire [8:0] int_input_exp = 31 - {1'b0, renorm_shamt_s0[i * 5+:5]};
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:149:9
			assign input_exp_s0[i * 9+:9] = (is_itof_s0 ? int_input_exp : fp_input_exp);
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:155:5
	wire valid_in_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:156:5
	wire [TAGW - 1:0] tag_in_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:157:5
	wire is_itof_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:158:5
	wire unsigned_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:159:5
	wire [2:0] rnd_mode_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:160:5
	wire [(LANES * 7) - 1:0] fp_clss_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:161:5
	wire [LANES - 1:0] input_sign_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:162:5
	wire [LANES - 1:0] mant_is_zero_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:163:5
	wire [(LANES * 32) - 1:0] input_mant_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:164:5
	wire [(LANES * 9) - 1:0] input_exp_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:166:5
	VX_pipe_register #(
		.DATAW(((1 + TAGW) + 5) + (LANES * 50)),
		.RESETW(1)
	) pipe_reg1(
		.clk(clk),
		.reset(reset),
		.enable(~stall),
		.data_in({valid_in_s0, tag_in_s0, is_itof_s0, unsigned_s0, rnd_mode_s0, fp_clss_s0, input_sign_s0, mant_is_zero_s0, input_mant_s0, input_exp_s0}),
		.data_out({valid_in_s1, tag_in_s1, is_itof_s1, unsigned_s1, rnd_mode_s1, fp_clss_s1, input_sign_s1, mant_is_zero_s1, input_mant_s1, input_exp_s1})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:179:5
	wire [(LANES * 65) - 1:0] destination_mant_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:180:5
	wire [(LANES * 9) - 1:0] final_exp_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:181:5
	wire [LANES - 1:0] of_before_round_s1;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:183:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk5
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:184:9
			reg [64:0] preshift_mant;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:185:9
			reg [5:0] denorm_shamt;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:186:9
			reg [8:0] final_exp;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:187:9
			reg of_before_round;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:189:9
			always @(*) begin
				// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:192:13
				final_exp = input_exp_s1[i * 9+:9] + EXP_BIAS;
				// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:193:13
				preshift_mant = {input_mant_s1[i * 32+:32], 33'b000000000000000000000000000000000};
				// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:194:13
				denorm_shamt = 0;
				// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:195:13
				of_before_round = 1'b0;
				// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:198:13
				if (is_itof_s1) begin
					begin
						// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:199:17
						if ($signed(input_exp_s1[i * 9+:9]) >= $signed(128)) begin
							// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:201:21
							final_exp = 254;
							// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:202:21
							preshift_mant = ~0;
							// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:203:21
							of_before_round = 1'b1;
						end
						else if ($signed(input_exp_s1[i * 9+:9]) < $signed(-150)) begin
							// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:206:21
							final_exp = 0;
							// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:207:21
							denorm_shamt = 25;
						end
						else if ($signed(input_exp_s1[i * 9+:9]) < $signed(1 - EXP_BIAS)) begin
							// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:210:21
							final_exp = 0;
							// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:211:21
							denorm_shamt = (1 - EXP_BIAS) - input_exp_s1[i * 9+:9];
						end
					end
				end
				else
					// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:214:17
					if ($signed(input_exp_s1[i * 9+:9]) >= $signed(31 + unsigned_s1)) begin
						// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:216:21
						denorm_shamt = 6'sd0;
						// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:217:21
						of_before_round = 1'b1;
					end
					else if ($signed(input_exp_s1[i * 9+:9]) < $signed(-1))
						// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:220:21
						denorm_shamt = 33;
					else
						// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:223:21
						denorm_shamt = 31 - input_exp_s1[i * 9+:9];
			end
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:229:9
			assign destination_mant_s1[i * 65+:65] = preshift_mant >> denorm_shamt;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:230:9
			assign final_exp_s1[i * 9+:9] = final_exp;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:231:9
			assign of_before_round_s1[i] = of_before_round;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:236:5
	wire valid_in_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:237:5
	wire [TAGW - 1:0] tag_in_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:238:5
	wire is_itof_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:239:5
	wire unsigned_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:240:5
	wire [2:0] rnd_mode_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:241:5
	wire [(LANES * 7) - 1:0] fp_clss_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:242:5
	wire [LANES - 1:0] mant_is_zero_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:243:5
	wire [LANES - 1:0] input_sign_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:244:5
	wire [(LANES * 65) - 1:0] destination_mant_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:245:5
	wire [(LANES * 9) - 1:0] final_exp_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:246:5
	wire [LANES - 1:0] of_before_round_s2;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:248:5
	VX_pipe_register #(
		.DATAW(((1 + TAGW) + 5) + (LANES * 84)),
		.RESETW(1)
	) pipe_reg2(
		.clk(clk),
		.reset(reset),
		.enable(~stall),
		.data_in({valid_in_s1, tag_in_s1, is_itof_s1, unsigned_s1, rnd_mode_s1, fp_clss_s1, mant_is_zero_s1, input_sign_s1, destination_mant_s1, final_exp_s1, of_before_round_s1}),
		.data_out({valid_in_s2, tag_in_s2, is_itof_s2, unsigned_s2, rnd_mode_s2, fp_clss_s2, mant_is_zero_s2, input_sign_s2, destination_mant_s2, final_exp_s2, of_before_round_s2})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:259:5
	wire [LANES - 1:0] rounded_sign;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:260:5
	wire [(LANES * 32) - 1:0] rounded_abs;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:261:5
	wire [(LANES * 2) - 1:0] fp_round_sticky_bits;
	wire [(LANES * 2) - 1:0] int_round_sticky_bits;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:265:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk6
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:266:9
			wire [22:0] final_mant;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:267:9
			wire [31:0] final_int;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:268:9
			wire [1:0] round_sticky_bits;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:269:9
			wire [31:0] fmt_pre_round_abs;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:270:9
			wire [31:0] pre_round_abs;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:273:9
			assign {final_mant, fp_round_sticky_bits[(i * 2) + 1]} = destination_mant_s2[(i * 65) + 63-:24];
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:274:9
			assign {final_int, int_round_sticky_bits[(i * 2) + 1]} = destination_mant_s2[(i * 65) + 64-:33];
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:277:9
			assign fp_round_sticky_bits[i * 2] = |destination_mant_s2[(i * 65) + 39-:40];
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:278:9
			assign int_round_sticky_bits[i * 2] = |destination_mant_s2[(i * 65) + 31-:32];
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:281:9
			assign round_sticky_bits = (is_itof_s2 ? fp_round_sticky_bits[i * 2+:2] : int_round_sticky_bits[i * 2+:2]);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:284:9
			assign fmt_pre_round_abs = {1'b0, final_exp_s2[(i * 9) + 7-:8], final_mant[22:0]};
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:287:9
			assign pre_round_abs = (is_itof_s2 ? fmt_pre_round_abs : final_int);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:290:9
			VX_fp_rounding #(.DAT_WIDTH(32)) fp_rounding(
				.abs_value_i(pre_round_abs),
				.sign_i(input_sign_s2[i]),
				.round_sticky_bits_i(round_sticky_bits),
				.rnd_mode_i(rnd_mode_s2),
				.effective_subtraction_i(1'b0),
				.abs_rounded_o(rounded_abs[i * 32+:32]),
				.sign_o(rounded_sign[i])
			);
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:306:5
	wire valid_in_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:307:5
	wire [TAGW - 1:0] tag_in_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:308:5
	wire is_itof_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:309:5
	wire unsigned_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:310:5
	wire [(LANES * 7) - 1:0] fp_clss_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:311:5
	wire [LANES - 1:0] mant_is_zero_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:312:5
	wire [LANES - 1:0] input_sign_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:313:5
	wire [LANES - 1:0] rounded_sign_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:314:5
	wire [(LANES * 32) - 1:0] rounded_abs_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:315:5
	wire [LANES - 1:0] of_before_round_s3;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:317:5
	VX_pipe_register #(
		.DATAW(((1 + TAGW) + 2) + (LANES * 43)),
		.RESETW(1)
	) pipe_reg3(
		.clk(clk),
		.reset(reset),
		.enable(~stall),
		.data_in({valid_in_s2, tag_in_s2, is_itof_s2, unsigned_s2, fp_clss_s2, mant_is_zero_s2, input_sign_s2, rounded_abs, rounded_sign, of_before_round_s2}),
		.data_out({valid_in_s3, tag_in_s3, is_itof_s3, unsigned_s3, fp_clss_s3, mant_is_zero_s3, input_sign_s3, rounded_abs_s3, rounded_sign_s3, of_before_round_s3})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:328:5
	wire [LANES - 1:0] of_after_round;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:329:5
	wire [LANES - 1:0] uf_after_round;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:330:5
	wire [(LANES * 32) - 1:0] fmt_result;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:331:5
	wire [(LANES * 32) - 1:0] rounded_int_res;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:332:5
	wire [LANES - 1:0] rounded_int_res_zero;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:334:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk7
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:336:9
			assign fmt_result[i * 32+:32] = (is_itof_s3 & mant_is_zero_s3[i] ? 0 : {rounded_sign_s3[i], rounded_abs_s3[(i * 32) + 30-:31]});
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:339:9
			assign uf_after_round[i] = rounded_abs_s3[(i * 32) + 30-:8] == 0;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:340:9
			assign of_after_round[i] = rounded_abs_s3[(i * 32) + 30-:8] == ~0;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:343:9
			assign rounded_int_res[i * 32+:32] = (rounded_sign_s3[i] ? -rounded_abs_s3[i * 32+:32] : rounded_abs_s3[i * 32+:32]);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:344:9
			assign rounded_int_res_zero[i] = rounded_int_res[i * 32+:32] == 0;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:349:5
	wire [(LANES * 32) - 1:0] fp_special_result;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:350:5
	wire [(LANES * 5) - 1:0] fp_special_status;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:351:5
	wire [LANES - 1:0] fp_result_is_special;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:353:5
	localparam [7:0] QNAN_EXPONENT = 255;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:354:5
	localparam [22:0] QNAN_MANTISSA = 4194304;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:356:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk8
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:358:9
			assign fp_result_is_special[i] = ~is_itof_s3 & (fp_clss_s3[(i * 7) + 5] | fp_clss_s3[(i * 7) + 2]);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:361:9
			assign fp_special_status[i * 5+:5] = (fp_clss_s3[i * 7] ? 5'h10 : 5'h00);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:364:9
			assign fp_special_result[i * 32+:32] = (fp_clss_s3[(i * 7) + 5] ? sv2v_cast_32(input_sign_s3) << 31 : {1'b0, QNAN_EXPONENT, QNAN_MANTISSA});
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:370:5
	reg [(LANES * 32) - 1:0] int_special_result;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:371:5
	wire [(LANES * 5) - 1:0] int_special_status;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:372:5
	wire [LANES - 1:0] int_result_is_special;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:374:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk9
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:376:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:377:13
				if (input_sign_s3[i] && !fp_clss_s3[(i * 7) + 2]) begin
					// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:378:17
					int_special_result[(i * 32) + 30-:31] = 0;
					// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:379:17
					int_special_result[(i * 32) + 31] = ~unsigned_s3;
				end
				else begin
					// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:381:17
					int_special_result[(i * 32) + 30-:31] = 33'sd2147483648 - 1;
					// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:382:17
					int_special_result[(i * 32) + 31] = unsigned_s3;
				end
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:387:9
			assign int_result_is_special[i] = ((fp_clss_s3[(i * 7) + 2] | fp_clss_s3[(i * 7) + 3]) | of_before_round_s3[i]) | ((input_sign_s3[i] & unsigned_s3) & ~rounded_int_res_zero[i]);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:393:9
			assign int_special_status[i * 5+:5] = 5'h10;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:398:5
	wire [(LANES * 5) - 1:0] tmp_fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:399:5
	wire [(LANES * 32) - 1:0] tmp_result;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:401:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk10
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:402:9
			wire [4:0] fp_regular_status;
			wire [4:0] int_regular_status;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:403:9
			wire [4:0] fp_status;
			wire [4:0] int_status;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:404:9
			wire [31:0] fp_result;
			wire [31:0] int_result;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:406:9
			wire inexact = (is_itof_s3 ? |fp_round_sticky_bits[i * 2+:2] : |fp_round_sticky_bits[i * 2+:2] | (~fp_clss_s3[(i * 7) + 3] & (of_before_round_s3[i] | of_after_round[i])));
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:409:9
			assign fp_regular_status[4] = is_itof_s3 & (of_before_round_s3[i] | of_after_round[i]);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:410:9
			assign fp_regular_status[3] = 1'b0;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:411:9
			assign fp_regular_status[2] = ~is_itof_s3 & (~fp_clss_s3[(i * 7) + 3] & (of_before_round_s3[i] | of_after_round[i]));
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:412:9
			assign fp_regular_status[1] = uf_after_round[i] & inexact;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:413:9
			assign fp_regular_status[0] = inexact;
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:415:9
			assign int_regular_status = (|int_round_sticky_bits[i * 2+:2] ? 5'h01 : 5'h00);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:417:9
			assign fp_result = (fp_result_is_special[i] ? fp_special_result[i * 32+:32] : fmt_result[i * 32+:32]);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:418:9
			assign int_result = (int_result_is_special[i] ? int_special_result[i * 32+:32] : rounded_int_res[i * 32+:32]);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:420:9
			assign fp_status = (fp_result_is_special[i] ? fp_special_status[i * 5+:5] : fp_regular_status);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:421:9
			assign int_status = (int_result_is_special[i] ? int_special_status[i * 5+:5] : int_regular_status);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:424:9
			assign tmp_result[i * 32+:32] = (is_itof_s3 ? fp_result : int_result);
			// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:425:9
			assign tmp_fflags[i * 5+:5] = (is_itof_s3 ? fp_status : int_status);
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:428:5
	assign stall = ~ready_out && valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:430:5
	VX_pipe_register #(
		.DATAW(((1 + TAGW) + (LANES * 32)) + (LANES * 5)),
		.RESETW(1)
	) pipe_reg4(
		.clk(clk),
		.reset(reset),
		.enable(!stall),
		.data_in({valid_in_s3, tag_in_s3, tmp_result, tmp_fflags}),
		.data_out({valid_out, tag_out, result, fflags})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:441:5
	assign ready_in = ~stall;
	// Trace: ../../rtl/fp_cores/VX_fp_cvt.sv:443:5
	assign has_fflags = 1'b1;
endmodule
module VX_fp_div (
	clk,
	reset,
	ready_in,
	valid_in,
	tag_in,
	frm,
	dataa,
	datab,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:4:15
	parameter TAGW = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:5:15
	parameter LANES = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:7:5
	input wire clk;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:8:5
	input wire reset;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:10:5
	output wire ready_in;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:11:5
	input wire valid_in;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:13:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:15:5
	input wire [2:0] frm;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:17:5
	input wire [(LANES * 32) - 1:0] dataa;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:18:5
	input wire [(LANES * 32) - 1:0] datab;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:19:5
	output wire [(LANES * 32) - 1:0] result;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:21:5
	output wire has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:22:5
	// removed localparam type fpu_types_fflags_t
	output wire [(LANES * 5) - 1:0] fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:24:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:26:5
	input wire ready_out;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:27:5
	output wire valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:29:5
	wire stall = ~ready_out && valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:30:5
	wire enable = ~stall;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:32:5
	genvar i;
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk1
			// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fp_div.sv:54:27
			wire fdiv_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fp_div.sv:54:60
			VX_reset_relay __fdiv_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(fdiv_reset)
			);
			// Trace: ../../rtl/fp_cores/VX_fp_div.sv:56:9
			
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:67:5
	VX_shift_register #(
		.DATAW(1 + TAGW),
		.DEPTH(15),
		.RESETW(1)
	) shift_reg(
		.clk(clk),
		.reset(reset),
		.enable(enable),
		.data_in({valid_in, tag_in}),
		.data_out({valid_out, tag_out})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:79:5
	assign ready_in = enable;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:82:5
	assign has_fflags = 0;
	// Trace: ../../rtl/fp_cores/VX_fp_div.sv:83:5
	assign fflags = 0;
endmodule
module VX_fp_fma (
	clk,
	reset,
	ready_in,
	valid_in,
	tag_in,
	frm,
	do_madd,
	do_sub,
	do_neg,
	dataa,
	datab,
	datac,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:4:15
	parameter TAGW = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:5:15
	parameter LANES = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:7:5
	input wire clk;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:8:5
	input wire reset;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:10:5
	output wire ready_in;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:11:5
	input wire valid_in;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:13:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:15:5
	input wire [2:0] frm;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:17:5
	input wire do_madd;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:18:5
	input wire do_sub;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:19:5
	input wire do_neg;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:21:5
	input wire [(LANES * 32) - 1:0] dataa;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:22:5
	input wire [(LANES * 32) - 1:0] datab;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:23:5
	input wire [(LANES * 32) - 1:0] datac;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:24:5
	output wire [(LANES * 32) - 1:0] result;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:26:5
	output wire has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:27:5
	// removed localparam type fpu_types_fflags_t
	output wire [(LANES * 5) - 1:0] fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:29:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:31:5
	input wire ready_out;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:32:5
	output wire valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:35:5
	wire stall = ~ready_out && valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:36:5
	wire enable = ~stall;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:38:5
	genvar i;
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk1
			// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:39:9
			reg [31:0] a;
			reg [31:0] b;
			reg [31:0] c;
			// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:41:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:42:13
				if (do_madd) begin
					// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:44:17
					a = (do_neg ? {~dataa[(i * 32) + 31], dataa[(i * 32) + 30-:31]} : dataa[i * 32+:32]);
					// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:45:17
					b = datab[i * 32+:32];
					// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:46:17
					c = (do_neg ^ do_sub ? {~datac[(i * 32) + 31], datac[(i * 32) + 30-:31]} : datac[i * 32+:32]);
				end
				else
					// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:48:17
					if (do_neg) begin
						// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:50:21
						a = dataa[i * 32+:32];
						// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:51:21
						b = datab[i * 32+:32];
						// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:52:21
						c = 0;
					end
					else begin
						// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:55:21
						a = 32'h3f800000;
						// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:56:21
						b = dataa[i * 32+:32];
						// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:57:21
						c = (do_sub ? {~datab[(i * 32) + 31], datab[(i * 32) + 30-:31]} : datab[i * 32+:32]);
					end
			// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fp_fma.sv:83:26
			wire fma_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fp_fma.sv:83:59
			VX_reset_relay __fma_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(fma_reset)
			);
			// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:85:9
			
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:97:5
	VX_shift_register #(
		.DATAW(1 + TAGW),
		.DEPTH(4),
		.RESETW(1)
	) shift_reg(
		.clk(clk),
		.reset(reset),
		.enable(enable),
		.data_in({valid_in, tag_in}),
		.data_out({valid_out, tag_out})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:109:5
	assign ready_in = enable;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:112:5
	assign has_fflags = 0;
	// Trace: ../../rtl/fp_cores/VX_fp_fma.sv:113:5
	assign fflags = 0;
endmodule
module VX_fp_ncomp (
	clk,
	reset,
	ready_in,
	valid_in,
	tag_in,
	op_type,
	frm,
	dataa,
	datab,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:7:15
	parameter TAGW = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:8:15
	parameter LANES = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:10:5
	input wire clk;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:11:5
	input wire reset;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:13:5
	output wire ready_in;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:14:5
	input wire valid_in;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:16:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:18:5
	input wire [3:0] op_type;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:19:5
	input wire [2:0] frm;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:21:5
	input wire [(LANES * 32) - 1:0] dataa;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:22:5
	input wire [(LANES * 32) - 1:0] datab;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:23:5
	output wire [(LANES * 32) - 1:0] result;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:25:5
	output wire has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:26:5
	// removed localparam type fpu_types_fflags_t
	output wire [(LANES * 5) - 1:0] fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:28:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:30:5
	input wire ready_out;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:31:5
	output wire valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:33:5
	localparam EXP_BITS = 8;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:34:5
	localparam MAN_BITS = 23;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:36:5
	localparam NEG_INF = 32'h00000001;
	localparam NEG_NORM = 32'h00000002;
	localparam NEG_SUBNORM = 32'h00000004;
	localparam NEG_ZERO = 32'h00000008;
	localparam POS_ZERO = 32'h00000010;
	localparam POS_SUBNORM = 32'h00000020;
	localparam POS_NORM = 32'h00000040;
	localparam POS_INF = 32'h00000080;
	localparam QUT_NAN = 32'h00000200;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:47:5
	wire [LANES - 1:0] a_sign;
	wire [LANES - 1:0] b_sign;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:48:5
	wire [(LANES * 8) - 1:0] a_exponent;
	wire [(LANES * 8) - 1:0] b_exponent;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:49:5
	wire [(LANES * 23) - 1:0] a_mantissa;
	wire [(LANES * 23) - 1:0] b_mantissa;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:50:5
	// removed localparam type fpu_types_fp_class_t
	wire [(LANES * 7) - 1:0] a_clss;
	wire [(LANES * 7) - 1:0] b_clss;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:51:5
	wire [LANES - 1:0] a_smaller;
	wire [LANES - 1:0] ab_equal;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:54:5
	genvar i;
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk1
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:55:9
			assign a_sign[i] = dataa[(i * 32) + 31];
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:56:9
			assign a_exponent[i * 8+:8] = dataa[(i * 32) + 30-:8];
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:57:9
			assign a_mantissa[i * 23+:23] = dataa[(i * 32) + 22-:23];
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:59:9
			assign b_sign[i] = datab[(i * 32) + 31];
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:60:9
			assign b_exponent[i * 8+:8] = datab[(i * 32) + 30-:8];
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:61:9
			assign b_mantissa[i * 23+:23] = datab[(i * 32) + 22-:23];
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:63:9
			VX_fp_class #(
				.EXP_BITS(EXP_BITS),
				.MAN_BITS(MAN_BITS)
			) fp_class_a(
				.exp_i(a_exponent[i * 8+:8]),
				.man_i(a_mantissa[i * 23+:23]),
				.clss_o(a_clss[i * 7+:7])
			);
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:72:9
			VX_fp_class #(
				.EXP_BITS(EXP_BITS),
				.MAN_BITS(MAN_BITS)
			) fp_class_b(
				.exp_i(b_exponent[i * 8+:8]),
				.man_i(b_mantissa[i * 23+:23]),
				.clss_o(b_clss[i * 7+:7])
			);
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:81:9
			assign a_smaller[i] = $signed(dataa[i * 32+:32]) < $signed(datab[i * 32+:32]);
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:82:9
			assign ab_equal[i] = (dataa[i * 32+:32] == datab[i * 32+:32]) | (a_clss[(i * 7) + 5] & b_clss[(i * 7) + 5]);
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:87:5
	wire valid_in_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:88:5
	wire [TAGW - 1:0] tag_in_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:89:5
	wire [3:0] op_type_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:90:5
	wire [2:0] frm_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:91:5
	wire [(LANES * 32) - 1:0] dataa_s0;
	wire [(LANES * 32) - 1:0] datab_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:92:5
	wire [LANES - 1:0] a_sign_s0;
	wire [LANES - 1:0] b_sign_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:93:5
	wire [(LANES * 8) - 1:0] a_exponent_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:94:5
	wire [(LANES * 23) - 1:0] a_mantissa_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:95:5
	wire [(LANES * 7) - 1:0] a_clss_s0;
	wire [(LANES * 7) - 1:0] b_clss_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:96:5
	wire [LANES - 1:0] a_smaller_s0;
	wire [LANES - 1:0] ab_equal_s0;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:98:5
	wire stall;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:100:5
	VX_pipe_register #(
		.DATAW(((1 + TAGW) + 7) + (LANES * 113)),
		.RESETW(1),
		.DEPTH(0)
	) pipe_reg0(
		.clk(clk),
		.reset(reset),
		.enable(!stall),
		.data_in({valid_in, tag_in, op_type, frm, dataa, datab, a_sign, b_sign, a_exponent, a_mantissa, a_clss, b_clss, a_smaller, ab_equal}),
		.data_out({valid_in_s0, tag_in_s0, op_type_s0, frm_s0, dataa_s0, datab_s0, a_sign_s0, b_sign_s0, a_exponent_s0, a_mantissa_s0, a_clss_s0, b_clss_s0, a_smaller_s0, ab_equal_s0})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:113:5
	reg [(LANES * 32) - 1:0] fclass_mask;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:114:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk2
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:115:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:116:13
				if (a_clss_s0[(i * 7) + 6])
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:117:17
					fclass_mask[i * 32+:32] = (a_sign_s0[i] ? NEG_NORM : POS_NORM);
				else if (a_clss_s0[(i * 7) + 3])
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:120:17
					fclass_mask[i * 32+:32] = (a_sign_s0[i] ? NEG_INF : POS_INF);
				else if (a_clss_s0[(i * 7) + 5])
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:123:17
					fclass_mask[i * 32+:32] = (a_sign_s0[i] ? NEG_ZERO : POS_ZERO);
				else if (a_clss_s0[(i * 7) + 4])
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:126:17
					fclass_mask[i * 32+:32] = (a_sign_s0[i] ? NEG_SUBNORM : POS_SUBNORM);
				else if (a_clss_s0[(i * 7) + 2])
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:129:17
					fclass_mask[i * 32+:32] = {22'h000000, a_clss_s0[(i * 7) + 1], a_clss_s0[i * 7], 8'h00};
				else
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:132:17
					fclass_mask[i * 32+:32] = QUT_NAN;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:138:5
	reg [(LANES * 32) - 1:0] fminmax_res;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:139:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk3
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:140:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:141:13
				if (a_clss_s0[(i * 7) + 2] && b_clss_s0[(i * 7) + 2])
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:142:17
					fminmax_res[i * 32+:32] = 32'h7fc00000;
				else if (a_clss_s0[(i * 7) + 2])
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:144:17
					fminmax_res[i * 32+:32] = datab_s0[i * 32+:32];
				else if (b_clss_s0[(i * 7) + 2])
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:146:17
					fminmax_res[i * 32+:32] = dataa_s0[i * 32+:32];
				else
					// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:148:17
					case (frm_s0)
						3:
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:149:24
							fminmax_res[i * 32+:32] = (a_smaller_s0[i] ? dataa_s0[i * 32+:32] : datab_s0[i * 32+:32]);
						4:
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:150:24
							fminmax_res[i * 32+:32] = (a_smaller_s0[i] ? datab_s0[i * 32+:32] : dataa_s0[i * 32+:32]);
						default:
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:151:24
							fminmax_res[i * 32+:32] = 1'sbx;
					endcase
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:158:5
	reg [(LANES * 32) - 1:0] fsgnj_res;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:159:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk4
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:160:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:161:13
				case (frm_s0)
					0:
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:162:20
						fsgnj_res[i * 32+:32] = {b_sign_s0[i], a_exponent_s0[i * 8+:8], a_mantissa_s0[i * 23+:23]};
					1:
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:163:20
						fsgnj_res[i * 32+:32] = {~b_sign_s0[i], a_exponent_s0[i * 8+:8], a_mantissa_s0[i * 23+:23]};
					2:
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:164:20
						fsgnj_res[i * 32+:32] = {a_sign_s0[i] ^ b_sign_s0[i], a_exponent_s0[i * 8+:8], a_mantissa_s0[i * 23+:23]};
					default:
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:165:20
						fsgnj_res[i * 32+:32] = 1'sbx;
				endcase
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:171:5
	reg [(LANES * 32) - 1:0] fcmp_res;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:172:5
	reg [(LANES * 5) - 1:0] fcmp_fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:173:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk5
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:174:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:175:13
				case (frm_s0)
					3'b000: begin
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:177:21
						fcmp_fflags[i * 5+:5] = 5'h00;
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:178:21
						if (a_clss_s0[(i * 7) + 2] || b_clss_s0[(i * 7) + 2]) begin
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:179:25
							fcmp_res[i * 32+:32] = 32'h00000000;
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:180:25
							fcmp_fflags[(i * 5) + 4] = 1'b1;
						end
						else
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:182:25
							fcmp_res[i * 32+:32] = {31'h00000000, a_smaller_s0[i] | ab_equal_s0[i]};
					end
					3'b001: begin
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:186:21
						fcmp_fflags[i * 5+:5] = 5'h00;
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:187:21
						if (a_clss_s0[(i * 7) + 2] || b_clss_s0[(i * 7) + 2]) begin
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:188:25
							fcmp_res[i * 32+:32] = 32'h00000000;
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:189:25
							fcmp_fflags[(i * 5) + 4] = 1'b1;
						end
						else
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:191:25
							fcmp_res[i * 32+:32] = {31'h00000000, a_smaller_s0[i] & ~ab_equal_s0[i]};
					end
					3'b010: begin
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:195:21
						fcmp_fflags[i * 5+:5] = 5'h00;
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:196:21
						if (a_clss_s0[(i * 7) + 2] || b_clss_s0[(i * 7) + 2]) begin
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:197:25
							fcmp_res[i * 32+:32] = 32'h00000000;
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:198:25
							fcmp_fflags[(i * 5) + 4] = a_clss_s0[i * 7] | b_clss_s0[i * 7];
						end
						else
							// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:200:25
							fcmp_res[i * 32+:32] = {31'h00000000, ab_equal_s0[i]};
					end
					default: begin
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:204:21
						fcmp_res[i * 32+:32] = 1'sbx;
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:205:21
						fcmp_fflags[i * 5+:5] = 1'sbx;
					end
				endcase
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:213:5
	reg [(LANES * 32) - 1:0] tmp_result;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:214:5
	reg [(LANES * 5) - 1:0] tmp_fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:216:5
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk6
			// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:217:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:218:13
				case (op_type_s0)
					4'h6: begin
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:220:21
						tmp_result[i * 32+:32] = fclass_mask[i * 32+:32];
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:221:21
						tmp_fflags[i * 5+:5] = 1'sbx;
					end
					4'ha: begin
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:224:21
						tmp_result[i * 32+:32] = fcmp_res[i * 32+:32];
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:225:21
						tmp_fflags[i * 5+:5] = fcmp_fflags[i * 5+:5];
					end
					default:
						// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:229:21
						case (frm_s0)
							0, 1, 2: begin
								// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:231:29
								tmp_result[i * 32+:32] = fsgnj_res[i * 32+:32];
								// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:232:29
								tmp_fflags[i * 5+:5] = 1'sbx;
							end
							3, 4: begin
								// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:235:29
								tmp_result[i * 32+:32] = fminmax_res[i * 32+:32];
								// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:236:29
								tmp_fflags[i * 5+:5] = 0;
								// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:237:29
								tmp_fflags[(i * 5) + 4] = a_clss_s0[i * 7] | b_clss_s0[i * 7];
							end
							default: begin
								// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:241:29
								tmp_result[i * 32+:32] = dataa_s0[i * 32+:32];
								// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:242:29
								tmp_fflags[i * 5+:5] = 1'sbx;
							end
						endcase
				endcase
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:250:5
	wire has_fflags_s0 = ((op_type_s0 == 4'he) && ((frm_s0 == 3) || (frm_s0 == 4))) || (op_type_s0 == 4'ha);
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:255:5
	assign stall = ~ready_out && valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:257:5
	VX_pipe_register #(
		.DATAW((((1 + TAGW) + (LANES * 32)) + 1) + (LANES * 5)),
		.RESETW(1)
	) pipe_reg1(
		.clk(clk),
		.reset(reset),
		.enable(!stall),
		.data_in({valid_in_s0, tag_in_s0, tmp_result, has_fflags_s0, tmp_fflags}),
		.data_out({valid_out, tag_out, result, has_fflags, fflags})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_ncomp.sv:268:5
	assign ready_in = ~stall;
endmodule
module VX_fp_rounding (
	abs_value_i,
	sign_i,
	round_sticky_bits_i,
	rnd_mode_i,
	effective_subtraction_i,
	abs_rounded_o,
	sign_o,
	exact_zero_o
);
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:7:15
	parameter DAT_WIDTH = 2;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:10:5
	input wire [DAT_WIDTH - 1:0] abs_value_i;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:11:5
	input wire sign_i;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:13:5
	input wire [1:0] round_sticky_bits_i;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:14:5
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:15:5
	input wire effective_subtraction_i;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:17:5
	output wire [DAT_WIDTH - 1:0] abs_rounded_o;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:18:5
	output wire sign_o;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:19:5
	output wire exact_zero_o;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:22:5
	reg round_up;
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:34:5
	always @(*)
		// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:35:9
		case (rnd_mode_i)
			3'b000:
				case (round_sticky_bits_i)
					2'b00, 2'b01:
						// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:39:30
						round_up = 1'b0;
					2'b10:
						// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:40:30
						round_up = abs_value_i[0];
					2'b11:
						// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:41:30
						round_up = 1'b1;
					default:
						// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:42:30
						round_up = 1'bx;
				endcase
			3'b001:
				// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:44:28
				round_up = 1'b0;
			3'b010:
				// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:45:28
				round_up = |round_sticky_bits_i & sign_i;
			3'b011:
				// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:46:28
				round_up = |round_sticky_bits_i & ~sign_i;
			3'b100:
				// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:47:28
				round_up = round_sticky_bits_i[1];
			default:
				// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:48:23
				round_up = 1'bx;
		endcase
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:53:5
	function automatic [DAT_WIDTH - 1:0] sv2v_cast_8455B;
		input reg [DAT_WIDTH - 1:0] inp;
		sv2v_cast_8455B = inp;
	endfunction
	assign abs_rounded_o = abs_value_i + sv2v_cast_8455B(round_up);
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:56:5
	assign exact_zero_o = (abs_value_i == 0) && (round_sticky_bits_i == 0);
	// Trace: ../../rtl/fp_cores/VX_fp_rounding.sv:60:5
	assign sign_o = (exact_zero_o && effective_subtraction_i ? rnd_mode_i == 3'b010 : sign_i);
endmodule
module VX_fp_sqrt (
	clk,
	reset,
	ready_in,
	valid_in,
	tag_in,
	frm,
	dataa,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:4:15
	parameter TAGW = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:5:15
	parameter LANES = 1;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:7:5
	input wire clk;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:8:5
	input wire reset;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:10:5
	output wire ready_in;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:11:5
	input wire valid_in;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:13:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:15:5
	input wire [2:0] frm;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:17:5
	input wire [(LANES * 32) - 1:0] dataa;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:18:5
	output wire [(LANES * 32) - 1:0] result;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:20:5
	output wire has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:21:5
	// removed localparam type fpu_types_fflags_t
	output wire [(LANES * 5) - 1:0] fflags;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:23:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:25:5
	input wire ready_out;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:26:5
	output wire valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:28:5
	wire stall = ~ready_out && valid_out;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:29:5
	wire enable = ~stall;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:31:5
	genvar i;
	generate
		for (i = 0; i < LANES; i = i + 1) begin : genblk1
			// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fp_sqrt.sv:53:28
			wire fsqrt_reset;
			// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fp_sqrt.sv:53:61
			VX_reset_relay __fsqrt_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(fsqrt_reset)
			);
			// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:55:9
			
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:65:5
	VX_shift_register #(
		.DATAW(1 + TAGW),
		.DEPTH(10),
		.RESETW(1)
	) shift_reg(
		.clk(clk),
		.reset(reset),
		.enable(enable),
		.data_in({valid_in, tag_in}),
		.data_out({valid_out, tag_out})
	);
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:77:5
	assign ready_in = enable;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:80:5
	assign has_fflags = 0;
	// Trace: ../../rtl/fp_cores/VX_fp_sqrt.sv:81:5
	assign fflags = 0;
endmodule
module VX_fpu_dpi (
	clk,
	reset,
	valid_in,
	ready_in,
	tag_in,
	op_type,
	frm,
	dataa,
	datab,
	datac,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:4:15
	parameter TAGW = 1;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:6:5
	input wire clk;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:7:5
	input wire reset;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:9:5
	input wire valid_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:10:5
	output wire ready_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:12:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:14:5
	input wire [3:0] op_type;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:15:5
	input wire [2:0] frm;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:17:5
	input wire [63:0] dataa;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:18:5
	input wire [63:0] datab;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:19:5
	input wire [63:0] datac;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:20:5
	output wire [63:0] result;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:22:5
	output wire has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:23:5
	// removed localparam type fpu_types_fflags_t
	output wire [9:0] fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:25:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:27:5
	input wire ready_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:28:5
	output wire valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:30:5
	localparam FPU_FMA = 0;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:31:5
	localparam FPU_DIV = 1;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:32:5
	localparam FPU_SQRT = 2;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:33:5
	localparam FPU_CVT = 3;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:34:5
	localparam FPU_NCP = 4;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:35:5
	localparam NUM_FPC = 5;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:36:5
	localparam FPC_BITS = 3;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:38:5
	wire [4:0] per_core_ready_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:39:5
	wire [319:0] per_core_result;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:40:5
	wire [(5 * TAGW) - 1:0] per_core_tag_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:41:5
	reg [4:0] per_core_ready_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:42:5
	wire [4:0] per_core_valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:44:5
	wire [4:0] per_core_has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:45:5
	wire [49:0] per_core_fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:47:5
	reg [2:0] core_select;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:49:5
	reg is_fadd;
	reg is_fsub;
	reg is_fmul;
	reg is_fmadd;
	reg is_fmsub;
	reg is_fnmadd;
	reg is_fnmsub;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:50:5
	reg is_itof;
	reg is_utof;
	reg is_ftoi;
	reg is_ftou;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:51:5
	reg is_fclss;
	reg is_flt;
	reg is_fle;
	reg is_feq;
	reg is_fmin;
	reg is_fmax;
	reg is_fsgnj;
	reg is_fsgnjn;
	reg is_fsgnjx;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:53:5
	always @(*) begin
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:54:9
		is_fadd = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:55:9
		is_fsub = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:56:9
		is_fmul = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:57:9
		is_fmadd = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:58:9
		is_fmsub = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:59:9
		is_fnmadd = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:60:9
		is_fnmsub = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:61:9
		is_itof = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:62:9
		is_utof = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:63:9
		is_ftoi = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:64:9
		is_ftou = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:65:9
		is_fclss = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:66:9
		is_flt = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:67:9
		is_fle = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:68:9
		is_feq = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:69:9
		is_fmin = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:70:9
		is_fmax = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:71:9
		is_fsgnj = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:72:9
		is_fsgnjn = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:73:9
		is_fsgnjx = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:75:9
		case (op_type)
			4'h0: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:76:36
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:76:59
				is_fadd = 1;
			end
			4'h4: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:77:36
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:77:59
				is_fsub = 1;
			end
			4'h8: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:78:36
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:78:59
				is_fmul = 1;
			end
			4'h3: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:79:36
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:79:59
				is_fmadd = 1;
			end
			4'h7: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:80:36
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:80:59
				is_fmsub = 1;
			end
			4'hf: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:81:36
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:81:59
				is_fnmadd = 1;
			end
			4'hb: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:82:36
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:82:59
				is_fnmsub = 1;
			end
			4'hc:
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:83:36
				core_select = FPU_DIV;
			4'h2:
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:84:36
				core_select = FPU_SQRT;
			4'h1: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:85:36
				core_select = FPU_CVT;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:85:59
				is_ftoi = 1;
			end
			4'h5: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:86:36
				core_select = FPU_CVT;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:86:59
				is_ftou = 1;
			end
			4'h9: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:87:36
				core_select = FPU_CVT;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:87:59
				is_itof = 1;
			end
			4'hd: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:88:36
				core_select = FPU_CVT;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:88:59
				is_utof = 1;
			end
			4'h6: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:89:36
				core_select = FPU_NCP;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:89:59
				is_fclss = 1;
			end
			4'ha: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:90:36
				core_select = FPU_NCP;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:91:29
				is_fle = frm == 0;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:92:29
				is_flt = frm == 1;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:93:29
				is_feq = frm == 2;
			end
			default: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:95:30
				core_select = FPU_NCP;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:96:29
				is_fsgnj = frm == 0;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:97:29
				is_fsgnjn = frm == 1;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:98:29
				is_fsgnjx = frm == 2;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:99:29
				is_fmin = frm == 3;
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:100:29
				is_fmax = frm == 4;
			end
		endcase
	end
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:105:5
	generate
		if (1) begin : fma
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:108:9
			wire [63:0] result_fma;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:109:9
			wire [63:0] result_fadd;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:110:9
			wire [63:0] result_fsub;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:111:9
			wire [63:0] result_fmul;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:112:9
			wire [63:0] result_fmadd;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:113:9
			wire [63:0] result_fmsub;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:114:9
			wire [63:0] result_fnmadd;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:115:9
			wire [63:0] result_fnmsub;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:117:9
			wire [9:0] fflags_fma;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:118:9
			wire [9:0] fflags_fadd;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:119:9
			wire [9:0] fflags_fsub;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:120:9
			wire [9:0] fflags_fmul;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:121:9
			wire [9:0] fflags_fmadd;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:122:9
			wire [9:0] fflags_fmsub;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:123:9
			wire [9:0] fflags_fnmadd;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:124:9
			wire [9:0] fflags_fnmsub;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:126:9
			wire fma_valid = valid_in && (core_select == FPU_FMA);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:127:9
			wire fma_ready = per_core_ready_out[FPU_FMA] || ~per_core_valid_out[FPU_FMA];
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:129:9
			wire fma_fire = fma_valid && fma_ready;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:131:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:132:13
				begin : sv2v_autoblock_1
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:132:18
					integer i;
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:132:18
					for (i = 0; i < 2; i = i + 1)
						begin
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:133:17
							dpi_fadd(fma_fire, dataa[i * 32+:32], datab[i * 32+:32], frm, result_fadd[i * 32+:32], fflags_fadd[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:134:17
							dpi_fsub(fma_fire, dataa[i * 32+:32], datab[i * 32+:32], frm, result_fsub[i * 32+:32], fflags_fsub[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:135:17
							dpi_fmul(fma_fire, dataa[i * 32+:32], datab[i * 32+:32], frm, result_fmul[i * 32+:32], fflags_fmul[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:136:17
							dpi_fmadd(fma_fire, dataa[i * 32+:32], datab[i * 32+:32], datac[i * 32+:32], frm, result_fmadd[i * 32+:32], fflags_fmadd[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:137:17
							dpi_fmsub(fma_fire, dataa[i * 32+:32], datab[i * 32+:32], datac[i * 32+:32], frm, result_fmsub[i * 32+:32], fflags_fmsub[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:138:17
							dpi_fnmadd(fma_fire, dataa[i * 32+:32], datab[i * 32+:32], datac[i * 32+:32], frm, result_fnmadd[i * 32+:32], fflags_fnmadd[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:139:17
							dpi_fnmsub(fma_fire, dataa[i * 32+:32], datab[i * 32+:32], datac[i * 32+:32], frm, result_fnmsub[i * 32+:32], fflags_fnmsub[i * 5+:5]);
						end
				end
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:143:9
			assign result_fma = (is_fadd ? result_fadd : (is_fsub ? result_fsub : (is_fmul ? result_fmul : (is_fmadd ? result_fmadd : (is_fmsub ? result_fmsub : (is_fnmadd ? result_fnmadd : (is_fnmsub ? result_fnmsub : 0)))))));
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:152:9
			assign fflags_fma = (is_fadd ? fflags_fadd : (is_fsub ? fflags_fsub : (is_fmul ? fflags_fmul : (is_fmadd ? fflags_fmadd : (is_fmsub ? fflags_fmsub : (is_fnmadd ? fflags_fnmadd : (is_fnmsub ? fflags_fnmsub : 0)))))));
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:161:9
			VX_shift_register #(
				.DATAW((1 + TAGW) + 74),
				.DEPTH(4),
				.RESETW(1)
			) shift_reg(
				.clk(clk),
				.reset(reset),
				.enable(fma_ready),
				.data_in({fma_valid, tag_in, result_fma, fflags_fma}),
				.data_out({per_core_valid_out[FPU_FMA], per_core_tag_out[0+:TAGW], per_core_result[0+:64], per_core_fflags[0+:10]})
			);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:173:9
			assign per_core_has_fflags[FPU_FMA] = 1;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:174:9
			assign per_core_ready_in[FPU_FMA] = fma_ready;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:179:5
	generate
		if (1) begin : fdiv
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:182:9
			wire [63:0] result_fdiv;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:183:9
			wire [9:0] fflags_fdiv;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:185:9
			wire fdiv_valid = valid_in && (core_select == FPU_DIV);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:186:9
			wire fdiv_ready = per_core_ready_out[FPU_DIV] || ~per_core_valid_out[FPU_DIV];
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:188:9
			wire fdiv_fire = fdiv_valid && fdiv_ready;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:190:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:191:13
				begin : sv2v_autoblock_2
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:191:18
					integer i;
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:191:18
					for (i = 0; i < 2; i = i + 1)
						begin
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:192:17
							dpi_fdiv(fdiv_fire, dataa[i * 32+:32], datab[i * 32+:32], frm, result_fdiv[i * 32+:32], fflags_fdiv[i * 5+:5]);
						end
				end
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:196:9
			VX_shift_register #(
				.DATAW((1 + TAGW) + 74),
				.DEPTH(15),
				.RESETW(1)
			) shift_reg(
				.clk(clk),
				.reset(reset),
				.enable(fdiv_ready),
				.data_in({fdiv_valid, tag_in, result_fdiv, fflags_fdiv}),
				.data_out({per_core_valid_out[FPU_DIV], per_core_tag_out[FPU_DIV * TAGW+:TAGW], per_core_result[64+:64], per_core_fflags[10+:10]})
			);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:208:9
			assign per_core_has_fflags[FPU_DIV] = 1;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:209:9
			assign per_core_ready_in[FPU_DIV] = fdiv_ready;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:214:5
	generate
		if (1) begin : fsqrt
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:217:9
			wire [63:0] result_fsqrt;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:218:9
			wire [9:0] fflags_fsqrt;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:220:9
			wire fsqrt_valid = valid_in && (core_select == FPU_SQRT);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:221:9
			wire fsqrt_ready = per_core_ready_out[FPU_SQRT] || ~per_core_valid_out[FPU_SQRT];
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:223:9
			wire fsqrt_fire = fsqrt_valid && fsqrt_ready;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:225:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:226:13
				begin : sv2v_autoblock_3
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:226:18
					integer i;
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:226:18
					for (i = 0; i < 2; i = i + 1)
						begin
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:227:17
							dpi_fsqrt(fsqrt_fire, dataa[i * 32+:32], frm, result_fsqrt[i * 32+:32], fflags_fsqrt[i * 5+:5]);
						end
				end
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:231:9
			VX_shift_register #(
				.DATAW((1 + TAGW) + 74),
				.DEPTH(10),
				.RESETW(1)
			) shift_reg(
				.clk(clk),
				.reset(reset),
				.enable(fsqrt_ready),
				.data_in({fsqrt_valid, tag_in, result_fsqrt, fflags_fsqrt}),
				.data_out({per_core_valid_out[FPU_SQRT], per_core_tag_out[FPU_SQRT * TAGW+:TAGW], per_core_result[128+:64], per_core_fflags[20+:10]})
			);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:243:9
			assign per_core_has_fflags[FPU_SQRT] = 1;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:244:9
			assign per_core_ready_in[FPU_SQRT] = fsqrt_ready;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:249:5
	generate
		if (1) begin : fcvt
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:252:9
			wire [63:0] result_fcvt;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:253:9
			wire [63:0] result_itof;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:254:9
			wire [63:0] result_utof;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:255:9
			wire [63:0] result_ftoi;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:256:9
			wire [63:0] result_ftou;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:258:9
			wire [9:0] fflags_fcvt;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:259:9
			wire [9:0] fflags_itof;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:260:9
			wire [9:0] fflags_utof;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:261:9
			wire [9:0] fflags_ftoi;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:262:9
			wire [9:0] fflags_ftou;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:264:9
			wire fcvt_valid = valid_in && (core_select == FPU_CVT);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:265:9
			wire fcvt_ready = per_core_ready_out[FPU_CVT] || ~per_core_valid_out[FPU_CVT];
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:267:9
			wire fcvt_fire = fcvt_valid && fcvt_ready;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:269:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:270:13
				begin : sv2v_autoblock_4
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:270:18
					integer i;
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:270:18
					for (i = 0; i < 2; i = i + 1)
						begin
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:271:17
							dpi_itof(fcvt_fire, dataa[i * 32+:32], frm, result_itof[i * 32+:32], fflags_itof[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:272:17
							dpi_utof(fcvt_fire, dataa[i * 32+:32], frm, result_utof[i * 32+:32], fflags_utof[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:273:17
							dpi_ftoi(fcvt_fire, dataa[i * 32+:32], frm, result_ftoi[i * 32+:32], fflags_ftoi[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:274:17
							dpi_ftou(fcvt_fire, dataa[i * 32+:32], frm, result_ftou[i * 32+:32], fflags_ftou[i * 5+:5]);
						end
				end
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:278:9
			assign result_fcvt = (is_itof ? result_itof : (is_utof ? result_utof : (is_ftoi ? result_ftoi : (is_ftou ? result_ftou : 0))));
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:284:9
			assign fflags_fcvt = (is_itof ? fflags_itof : (is_utof ? fflags_utof : (is_ftoi ? fflags_ftoi : (is_ftou ? fflags_ftou : 0))));
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:290:9
			VX_shift_register #(
				.DATAW((1 + TAGW) + 74),
				.DEPTH(5),
				.RESETW(1)
			) shift_reg(
				.clk(clk),
				.reset(reset),
				.enable(fcvt_ready),
				.data_in({fcvt_valid, tag_in, result_fcvt, fflags_fcvt}),
				.data_out({per_core_valid_out[FPU_CVT], per_core_tag_out[FPU_CVT * TAGW+:TAGW], per_core_result[192+:64], per_core_fflags[30+:10]})
			);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:302:9
			assign per_core_has_fflags[FPU_CVT] = 1;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:303:9
			assign per_core_ready_in[FPU_CVT] = fcvt_ready;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:308:5
	generate
		if (1) begin : fncp
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:311:9
			wire [63:0] result_fncp;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:312:9
			wire [63:0] result_fclss;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:313:9
			wire [63:0] result_flt;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:314:9
			wire [63:0] result_fle;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:315:9
			wire [63:0] result_feq;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:316:9
			wire [63:0] result_fmin;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:317:9
			wire [63:0] result_fmax;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:318:9
			wire [63:0] result_fsgnj;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:319:9
			wire [63:0] result_fsgnjn;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:320:9
			wire [63:0] result_fsgnjx;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:321:9
			reg [63:0] result_fmv;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:323:9
			wire [9:0] fflags_fncp;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:324:9
			wire [9:0] fflags_flt;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:325:9
			wire [9:0] fflags_fle;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:326:9
			wire [9:0] fflags_feq;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:327:9
			wire [9:0] fflags_fmin;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:328:9
			wire [9:0] fflags_fmax;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:330:9
			wire fncp_valid = valid_in && (core_select == FPU_NCP);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:331:9
			wire fncp_ready = per_core_ready_out[FPU_NCP] || ~per_core_valid_out[FPU_NCP];
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:333:9
			wire fncp_fire = fncp_valid && fncp_ready;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:335:9
			always @(*)
				// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:336:13
				begin : sv2v_autoblock_5
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:336:18
					integer i;
					// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:336:18
					for (i = 0; i < 2; i = i + 1)
						begin
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:337:17
							dpi_fclss(fncp_fire, dataa[i * 32+:32], result_fclss[i * 32+:32]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:338:17
							dpi_flt(fncp_fire, dataa[i * 32+:32], datab[i * 32+:32], result_flt[i * 32+:32], fflags_flt[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:339:17
							dpi_fle(fncp_fire, dataa[i * 32+:32], datab[i * 32+:32], result_fle[i * 32+:32], fflags_fle[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:340:17
							dpi_feq(fncp_fire, dataa[i * 32+:32], datab[i * 32+:32], result_feq[i * 32+:32], fflags_feq[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:341:17
							dpi_fmin(fncp_fire, dataa[i * 32+:32], datab[i * 32+:32], result_fmin[i * 32+:32], fflags_fmin[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:342:17
							dpi_fmax(fncp_fire, dataa[i * 32+:32], datab[i * 32+:32], result_fmax[i * 32+:32], fflags_fmax[i * 5+:5]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:343:17
							dpi_fsgnj(fncp_fire, dataa[i * 32+:32], datab[i * 32+:32], result_fsgnj[i * 32+:32]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:344:17
							dpi_fsgnjn(fncp_fire, dataa[i * 32+:32], datab[i * 32+:32], result_fsgnjn[i * 32+:32]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:345:17
							dpi_fsgnjx(fncp_fire, dataa[i * 32+:32], datab[i * 32+:32], result_fsgnjx[i * 32+:32]);
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:346:17
							result_fmv[i * 32+:32] = dataa[i * 32+:32];
						end
				end
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:350:9
			assign result_fncp = (is_fclss ? result_fclss : (is_flt ? result_flt : (is_fle ? result_fle : (is_feq ? result_feq : (is_fmin ? result_fmin : (is_fmax ? result_fmax : (is_fsgnj ? result_fsgnj : (is_fsgnjn ? result_fsgnjn : (is_fsgnjx ? result_fsgnjx : result_fmv)))))))));
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:361:9
			wire has_fflags_fncp = (((is_flt || is_fle) || is_feq) || is_fmin) || is_fmax;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:363:9
			assign fflags_fncp = (is_flt ? fflags_flt : (is_fle ? fflags_fle : (is_feq ? fflags_feq : (is_fmin ? fflags_fmin : (is_fmax ? fflags_fmax : 0)))));
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:370:9
			VX_shift_register #(
				.DATAW((1 + TAGW) + 75),
				.DEPTH(2),
				.RESETW(1)
			) shift_reg(
				.clk(clk),
				.reset(reset),
				.enable(fncp_ready),
				.data_in({fncp_valid, tag_in, has_fflags_fncp, result_fncp, fflags_fncp}),
				.data_out({per_core_valid_out[FPU_NCP], per_core_tag_out[FPU_NCP * TAGW+:TAGW], per_core_has_fflags[FPU_NCP], per_core_result[256+:64], per_core_fflags[40+:10]})
			);
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:382:9
			assign per_core_ready_in[FPU_NCP] = fncp_ready;
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:389:5
	reg has_fflags_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:390:5
	reg [9:0] fflags_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:391:5
	reg [63:0] result_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:392:5
	reg [TAGW - 1:0] tag_out_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:394:5
	always @(*) begin : sv2v_autoblock_6
		reg [0:1] _sv2v_jump;
		_sv2v_jump = 2'b00;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:395:9
		per_core_ready_out = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:396:9
		has_fflags_n = 1'sbx;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:397:9
		fflags_n = 1'sbx;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:398:9
		result_n = 1'sbx;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:399:9
		tag_out_n = 1'sbx;
		// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:400:9
		begin : sv2v_autoblock_7
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:400:14
			integer i;
			// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:400:14
			begin : sv2v_autoblock_8
				integer _sv2v_value_on_break;
				for (i = 0; i < NUM_FPC; i = i + 1)
					if (_sv2v_jump < 2'b10) begin
						_sv2v_jump = 2'b00;
						// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:401:13
						if (per_core_valid_out[i]) begin
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:402:17
							has_fflags_n = per_core_has_fflags[i];
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:403:17
							fflags_n = per_core_fflags[5 * (i * 2)+:10];
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:404:17
							result_n = per_core_result[32 * (i * 2)+:64];
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:405:17
							tag_out_n = per_core_tag_out[i * TAGW+:TAGW];
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:406:17
							per_core_ready_out[i] = ready_out;
							// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:407:17
							_sv2v_jump = 2'b10;
						end
						_sv2v_value_on_break = i;
					end
				if (!(_sv2v_jump < 2'b10))
					i = _sv2v_value_on_break;
				if (_sv2v_jump != 2'b11)
					_sv2v_jump = 2'b00;
			end
		end
	end
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:412:5
	assign valid_out = |per_core_valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:413:5
	assign has_fflags = has_fflags_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:414:5
	assign tag_out = tag_out_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:415:5
	assign result = result_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:416:5
	assign fflags = fflags_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_dpi.sv:418:5
	assign ready_in = per_core_ready_in[core_select];
endmodule
module VX_fpu_fpga (
	clk,
	reset,
	valid_in,
	ready_in,
	tag_in,
	op_type,
	frm,
	dataa,
	datab,
	datac,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:4:15
	parameter TAGW = 4;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:6:5
	input wire clk;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:7:5
	input wire reset;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:9:5
	input wire valid_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:10:5
	output wire ready_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:12:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:14:5
	input wire [3:0] op_type;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:15:5
	input wire [2:0] frm;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:17:5
	input wire [63:0] dataa;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:18:5
	input wire [63:0] datab;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:19:5
	input wire [63:0] datac;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:20:5
	output wire [63:0] result;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:22:5
	output wire has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:23:5
	// removed localparam type fpu_types_fflags_t
	output wire [9:0] fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:25:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:27:5
	input wire ready_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:28:5
	output wire valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:30:5
	localparam FPU_FMA = 0;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:31:5
	localparam FPU_DIV = 1;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:32:5
	localparam FPU_SQRT = 2;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:33:5
	localparam FPU_CVT = 3;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:34:5
	localparam FPU_NCP = 4;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:35:5
	localparam NUM_FPC = 5;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:36:5
	localparam FPC_BITS = 3;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:38:5
	wire [4:0] per_core_ready_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:39:5
	wire [319:0] per_core_result;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:40:5
	wire [(5 * TAGW) - 1:0] per_core_tag_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:41:5
	reg [4:0] per_core_ready_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:42:5
	wire [4:0] per_core_valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:44:5
	wire [4:0] per_core_has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:45:5
	wire [49:0] per_core_fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:47:5
	reg [2:0] core_select;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:48:5
	reg do_madd;
	reg do_sub;
	reg do_neg;
	reg is_itof;
	reg is_signed;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:50:5
	always @(*) begin
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:51:9
		do_madd = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:52:9
		do_sub = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:53:9
		do_neg = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:54:9
		is_itof = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:55:9
		is_signed = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:56:9
		case (op_type)
			4'h0:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:57:37
				core_select = FPU_FMA;
			4'h4: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:58:37
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:58:60
				do_sub = 1;
			end
			4'h8: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:59:37
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:59:60
				do_neg = 1;
			end
			4'h3: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:60:37
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:60:60
				do_madd = 1;
			end
			4'h7: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:61:37
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:61:60
				do_madd = 1;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:61:73
				do_sub = 1;
			end
			4'hf: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:62:37
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:62:60
				do_madd = 1;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:62:73
				do_neg = 1;
			end
			4'hb: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:63:37
				core_select = FPU_FMA;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:63:60
				do_madd = 1;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:63:73
				do_sub = 1;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:63:85
				do_neg = 1;
			end
			4'hc:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:64:37
				core_select = FPU_DIV;
			4'h2:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:65:37
				core_select = FPU_SQRT;
			4'h1: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:66:37
				core_select = FPU_CVT;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:66:60
				is_signed = 1;
			end
			4'h5:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:67:37
				core_select = FPU_CVT;
			4'h9: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:68:37
				core_select = FPU_CVT;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:68:60
				is_itof = 1;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:68:73
				is_signed = 1;
			end
			4'hd: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:69:37
				core_select = FPU_CVT;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:69:60
				is_itof = 1;
			end
			default:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:70:32
				core_select = FPU_NCP;
		endcase
	end
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:74:22
	wire fma_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:74:55
	VX_reset_relay __fma_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(fma_reset)
	);
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:75:22
	wire div_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:75:55
	VX_reset_relay __div_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(div_reset)
	);
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:76:23
	wire sqrt_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:76:56
	VX_reset_relay __sqrt_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(sqrt_reset)
	);
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:77:22
	wire cvt_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:77:55
	VX_reset_relay __cvt_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(cvt_reset)
	);
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:78:22
	wire ncp_reset;
	// Trace: macro expansion of RESET_RELAY at ../../rtl/fp_cores/VX_fpu_fpga.sv:78:55
	VX_reset_relay __ncp_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(ncp_reset)
	);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:80:5
	VX_fp_fma #(
		.TAGW(TAGW),
		.LANES(2)
	) fp_fma(
		.clk(clk),
		.reset(fma_reset),
		.valid_in(valid_in && (core_select == FPU_FMA)),
		.ready_in(per_core_ready_in[FPU_FMA]),
		.tag_in(tag_in),
		.frm(frm),
		.do_madd(do_madd),
		.do_sub(do_sub),
		.do_neg(do_neg),
		.dataa(dataa),
		.datab(datab),
		.datac(datac),
		.has_fflags(per_core_has_fflags[FPU_FMA]),
		.fflags(per_core_fflags[0+:10]),
		.result(per_core_result[0+:64]),
		.tag_out(per_core_tag_out[0+:TAGW]),
		.ready_out(per_core_ready_out[FPU_FMA]),
		.valid_out(per_core_valid_out[FPU_FMA])
	);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:104:5
	VX_fp_div #(
		.TAGW(TAGW),
		.LANES(2)
	) fp_div(
		.clk(clk),
		.reset(div_reset),
		.valid_in(valid_in && (core_select == FPU_DIV)),
		.ready_in(per_core_ready_in[FPU_DIV]),
		.tag_in(tag_in),
		.frm(frm),
		.dataa(dataa),
		.datab(datab),
		.has_fflags(per_core_has_fflags[FPU_DIV]),
		.fflags(per_core_fflags[10+:10]),
		.result(per_core_result[64+:64]),
		.tag_out(per_core_tag_out[FPU_DIV * TAGW+:TAGW]),
		.ready_out(per_core_ready_out[FPU_DIV]),
		.valid_out(per_core_valid_out[FPU_DIV])
	);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:124:5
	VX_fp_sqrt #(
		.TAGW(TAGW),
		.LANES(2)
	) fp_sqrt(
		.clk(clk),
		.reset(sqrt_reset),
		.valid_in(valid_in && (core_select == FPU_SQRT)),
		.ready_in(per_core_ready_in[FPU_SQRT]),
		.tag_in(tag_in),
		.frm(frm),
		.dataa(dataa),
		.has_fflags(per_core_has_fflags[FPU_SQRT]),
		.fflags(per_core_fflags[20+:10]),
		.result(per_core_result[128+:64]),
		.tag_out(per_core_tag_out[FPU_SQRT * TAGW+:TAGW]),
		.ready_out(per_core_ready_out[FPU_SQRT]),
		.valid_out(per_core_valid_out[FPU_SQRT])
	);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:143:5
	VX_fp_cvt #(
		.TAGW(TAGW),
		.LANES(2)
	) fp_cvt(
		.clk(clk),
		.reset(cvt_reset),
		.valid_in(valid_in && (core_select == FPU_CVT)),
		.ready_in(per_core_ready_in[FPU_CVT]),
		.tag_in(tag_in),
		.frm(frm),
		.is_itof(is_itof),
		.is_signed(is_signed),
		.dataa(dataa),
		.has_fflags(per_core_has_fflags[FPU_CVT]),
		.fflags(per_core_fflags[30+:10]),
		.result(per_core_result[192+:64]),
		.tag_out(per_core_tag_out[FPU_CVT * TAGW+:TAGW]),
		.ready_out(per_core_ready_out[FPU_CVT]),
		.valid_out(per_core_valid_out[FPU_CVT])
	);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:164:5
	VX_fp_ncomp #(
		.TAGW(TAGW),
		.LANES(2)
	) fp_ncomp(
		.clk(clk),
		.reset(ncp_reset),
		.valid_in(valid_in && (core_select == FPU_NCP)),
		.ready_in(per_core_ready_in[FPU_NCP]),
		.tag_in(tag_in),
		.op_type(op_type),
		.frm(frm),
		.dataa(dataa),
		.datab(datab),
		.result(per_core_result[256+:64]),
		.has_fflags(per_core_has_fflags[FPU_NCP]),
		.fflags(per_core_fflags[40+:10]),
		.tag_out(per_core_tag_out[FPU_NCP * TAGW+:TAGW]),
		.ready_out(per_core_ready_out[FPU_NCP]),
		.valid_out(per_core_valid_out[FPU_NCP])
	);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:185:5
	reg has_fflags_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:186:5
	reg [9:0] fflags_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:187:5
	reg [63:0] result_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:188:5
	reg [TAGW - 1:0] tag_out_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:190:5
	always @(*) begin : sv2v_autoblock_1
		reg [0:1] _sv2v_jump;
		_sv2v_jump = 2'b00;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:191:9
		per_core_ready_out = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:192:9
		has_fflags_n = 1'sbx;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:193:9
		fflags_n = 1'sbx;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:194:9
		result_n = 1'sbx;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:195:9
		tag_out_n = 1'sbx;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:196:9
		begin : sv2v_autoblock_2
			// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:196:14
			integer i;
			// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:196:14
			begin : sv2v_autoblock_3
				integer _sv2v_value_on_break;
				for (i = 0; i < NUM_FPC; i = i + 1)
					if (_sv2v_jump < 2'b10) begin
						_sv2v_jump = 2'b00;
						// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:197:13
						if (per_core_valid_out[i]) begin
							// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:198:17
							has_fflags_n = per_core_has_fflags[i];
							// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:199:17
							fflags_n = per_core_fflags[5 * (i * 2)+:10];
							// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:200:17
							result_n = per_core_result[32 * (i * 2)+:64];
							// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:201:17
							tag_out_n = per_core_tag_out[i * TAGW+:TAGW];
							// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:202:17
							per_core_ready_out[i] = ready_out;
							// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:203:17
							_sv2v_jump = 2'b10;
						end
						_sv2v_value_on_break = i;
					end
				if (!(_sv2v_jump < 2'b10))
					i = _sv2v_value_on_break;
				if (_sv2v_jump != 2'b11)
					_sv2v_jump = 2'b00;
			end
		end
	end
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:208:5
	assign valid_out = |per_core_valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:209:5
	assign has_fflags = has_fflags_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:210:5
	assign tag_out = tag_out_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:211:5
	assign result = result_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:212:5
	assign fflags = fflags_n;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpga.sv:214:5
	assign ready_in = per_core_ready_in[core_select];
endmodule
// removed package "fpnew_pkg"
// removed package "defs_div_sqrt_mvp"
module VX_fpu_fpnew (
	clk,
	reset,
	valid_in,
	ready_in,
	tag_in,
	op_type,
	frm,
	dataa,
	datab,
	datac,
	result,
	has_fflags,
	fflags,
	tag_out,
	ready_out,
	valid_out
);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:7:15
	parameter TAGW = 1;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:8:15
	parameter FMULADD = 1;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:9:15
	parameter FDIVSQRT = 1;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:10:15
	parameter FNONCOMP = 1;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:11:15
	parameter FCONV = 1;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:13:5
	input wire clk;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:14:5
	input wire reset;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:16:5
	input wire valid_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:17:5
	output wire ready_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:19:5
	input wire [TAGW - 1:0] tag_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:21:5
	input wire [3:0] op_type;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:22:5
	input wire [2:0] frm;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:24:5
	input wire [63:0] dataa;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:25:5
	input wire [63:0] datab;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:26:5
	input wire [63:0] datac;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:27:5
	output wire [63:0] result;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:29:5
	output wire has_fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:30:5
	// removed localparam type fpu_types_fflags_t
	output wire [9:0] fflags;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:32:5
	output wire [TAGW - 1:0] tag_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:34:5
	input wire ready_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:35:5
	output wire valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:37:5
	// removed localparam type fpnew_pkg_unit_type_t
	localparam UNIT_FMULADD = (FMULADD ? 2'd1 : 2'd0);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:38:5
	localparam UNIT_FDIVSQRT = (FDIVSQRT ? 2'd2 : 2'd0);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:39:5
	localparam UNIT_FNONCOMP = (FNONCOMP ? 2'd1 : 2'd0);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:40:5
	localparam UNIT_FCONV = (FCONV ? 2'd2 : 2'd0);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:42:5
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	localparam FOP_BITS = fpnew_pkg_OP_BITS;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:43:5
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam FMTF_BITS = 3;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:44:5
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	localparam FMTI_BITS = 2;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:46:5
	localparam FPU_DPATHW = 32'd32;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:48:5
	// removed localparam type fpnew_pkg_fmt_logic_t
	// removed localparam type fpnew_pkg_ifmt_logic_t
	// removed localparam type fpnew_pkg_fpu_features_t
	localparam [42:0] FPU_FEATURES = {FPU_DPATHW, 11'b01100000010};
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:56:5
	// removed localparam type fpnew_pkg_pipe_config_t
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unit_types_t
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unsigned_t
	// removed localparam type fpnew_pkg_fpu_implementation_t
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_CDC93;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_CDC93 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_15FEF;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_15FEF = inp;
	endfunction
	localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] FPU_IMPLEMENTATION = {sv2v_cast_CDC93({160'h0000000400000000000000000000000000000000, {fpnew_pkg_NUM_FP_FORMATS {32'd32}}, {fpnew_pkg_NUM_FP_FORMATS {32'd2}}, {fpnew_pkg_NUM_FP_FORMATS {32'd5}}}), sv2v_cast_15FEF({{fpnew_pkg_NUM_FP_FORMATS {UNIT_FMULADD}}, {fpnew_pkg_NUM_FP_FORMATS {UNIT_FDIVSQRT}}, {fpnew_pkg_NUM_FP_FORMATS {UNIT_FNONCOMP}}, {fpnew_pkg_NUM_FP_FORMATS {UNIT_FCONV}}}), 2'd3};
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:68:5
	wire fpu_ready_in;
	wire fpu_valid_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:69:5
	wire fpu_ready_out;
	wire fpu_valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:71:5
	reg [TAGW - 1:0] fpu_tag_in;
	reg [TAGW - 1:0] fpu_tag_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:73:5
	reg [191:0] fpu_operands;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:75:5
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	wire [2:0] fpu_src_fmt = sv2v_cast_0BC43('d0);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:76:5
	wire [2:0] fpu_dst_fmt = sv2v_cast_0BC43('d0);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:77:5
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	wire [1:0] fpu_int_fmt = sv2v_cast_87CC5(2);
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:79:5
	wire [63:0] fpu_result;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:80:5
	// removed localparam type fpnew_pkg_status_t
	wire [9:0] fpu_status;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:82:5
	reg [3:0] fpu_op;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:83:5
	reg [2:0] fpu_rnd;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:84:5
	reg fpu_op_mod;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:85:5
	reg fpu_has_fflags;
	reg fpu_has_fflags_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:87:5
	// removed localparam type fpnew_pkg_operation_e
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	always @(*) begin
		// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:88:9
		fpu_op = sv2v_cast_A53F3(6);
		// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:89:9
		fpu_rnd = frm;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:90:9
		fpu_op_mod = 0;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:91:9
		fpu_has_fflags = 1;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:92:9
		fpu_operands[0+:64] = dataa;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:93:9
		fpu_operands[64+:64] = datab;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:94:9
		fpu_operands[128+:64] = datac;
		// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:96:9
		case (op_type)
			4'h0: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:98:21
				fpu_op = sv2v_cast_A53F3(2);
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:99:21
				fpu_operands[64+:64] = dataa;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:100:21
				fpu_operands[128+:64] = datab;
			end
			4'h4: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:103:21
				fpu_op = sv2v_cast_A53F3(2);
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:104:21
				fpu_operands[64+:64] = dataa;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:105:21
				fpu_operands[128+:64] = datab;
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:106:21
				fpu_op_mod = 1;
			end
			4'h8:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:108:36
				fpu_op = sv2v_cast_A53F3(3);
			4'hc:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:109:36
				fpu_op = sv2v_cast_A53F3(4);
			4'h2:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:110:36
				fpu_op = sv2v_cast_A53F3(5);
			4'h3:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:111:36
				fpu_op = sv2v_cast_A53F3(0);
			4'h7: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:112:36
				fpu_op = sv2v_cast_A53F3(0);
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:112:64
				fpu_op_mod = 1;
			end
			4'hf: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:113:36
				fpu_op = sv2v_cast_A53F3(1);
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:113:64
				fpu_op_mod = 1;
			end
			4'hb:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:114:36
				fpu_op = sv2v_cast_A53F3(1);
			4'h1:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:115:36
				fpu_op = sv2v_cast_A53F3(11);
			4'h5: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:116:36
				fpu_op = sv2v_cast_A53F3(11);
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:116:61
				fpu_op_mod = 1;
			end
			4'h9:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:117:36
				fpu_op = sv2v_cast_A53F3(12);
			4'hd: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:118:36
				fpu_op = sv2v_cast_A53F3(12);
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:118:61
				fpu_op_mod = 1;
			end
			4'h6: begin
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:119:36
				fpu_op = sv2v_cast_A53F3(9);
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:119:66
				fpu_has_fflags = 0;
			end
			4'ha:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:120:36
				fpu_op = sv2v_cast_A53F3(8);
			4'he:
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:122:17
				case (frm)
					0: begin
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:123:32
						fpu_op = sv2v_cast_A53F3(6);
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:123:60
						fpu_rnd = 3'b000;
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:123:85
						fpu_has_fflags = 0;
					end
					1: begin
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:124:32
						fpu_op = sv2v_cast_A53F3(6);
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:124:60
						fpu_rnd = 3'b001;
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:124:85
						fpu_has_fflags = 0;
					end
					2: begin
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:125:32
						fpu_op = sv2v_cast_A53F3(6);
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:125:60
						fpu_rnd = 3'b010;
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:125:85
						fpu_has_fflags = 0;
					end
					3: begin
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:126:32
						fpu_op = sv2v_cast_A53F3(7);
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:126:60
						fpu_rnd = 3'b000;
					end
					4: begin
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:127:32
						fpu_op = sv2v_cast_A53F3(7);
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:127:60
						fpu_rnd = 3'b001;
					end
					default: begin
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:128:32
						fpu_op = sv2v_cast_A53F3(6);
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:128:60
						fpu_rnd = 3'b011;
						// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:128:85
						fpu_has_fflags = 0;
					end
				endcase
			default:
				;
		endcase
	end
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:135:5
	genvar i;
	// removed localparam type fpnew_pkg_roundmode_e
	generate
		for (i = 0; i < 2; i = i + 1) begin : genblk1
			if (0 == i) begin : genblk1
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:137:13
				// rewrote reg-to-output bindings
				wire [(0 + TAGW) + 1:1] sv2v_tmp_fpnew_core_tag_o;
				always @(*) {fpu_tag_out, fpu_has_fflags_out} = sv2v_tmp_fpnew_core_tag_o;
				fpnew_top_3ED0B_1EC5F #(
					.TagType_TAGW(TAGW),
					.Features(FPU_FEATURES),
					.Implementation(FPU_IMPLEMENTATION)
				) fpnew_core(
					.clk_i(clk),
					.rst_ni(1'b1),
					.operands_i({fpu_operands[128+:32], fpu_operands[64+:32], fpu_operands[0+:32]}),
					.rnd_mode_i(fpu_rnd),
					.op_i(sv2v_cast_A53F3(fpu_op)),
					.op_mod_i(fpu_op_mod),
					.src_fmt_i(sv2v_cast_0BC43(fpu_src_fmt)),
					.dst_fmt_i(sv2v_cast_0BC43(fpu_dst_fmt)),
					.int_fmt_i(sv2v_cast_87CC5(fpu_int_fmt)),
					.vectorial_op_i(1'b0),
					.tag_i({fpu_tag_in, fpu_has_fflags}),
					.in_valid_i(fpu_valid_in),
					.in_ready_o(fpu_ready_in),
					.flush_i(reset),
					.result_o(fpu_result[0+:32]),
					.status_o(fpu_status[0+:5]),
					.tag_o(sv2v_tmp_fpnew_core_tag_o),
					.out_valid_o(fpu_valid_out),
					.out_ready_i(fpu_ready_out)
				);
			end
			else begin : genblk1
				// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:164:13
				fpnew_top_FF541 #(
					.Features(FPU_FEATURES),
					.Implementation(FPU_IMPLEMENTATION)
				) fpnew_core(
					.clk_i(clk),
					.rst_ni(1'b1),
					.operands_i({fpu_operands[(4 + i) * 32+:32], fpu_operands[(2 + i) * 32+:32], fpu_operands[(0 + i) * 32+:32]}),
					.rnd_mode_i(fpu_rnd),
					.op_i(sv2v_cast_A53F3(fpu_op)),
					.op_mod_i(fpu_op_mod),
					.src_fmt_i(sv2v_cast_0BC43(fpu_src_fmt)),
					.dst_fmt_i(sv2v_cast_0BC43(fpu_dst_fmt)),
					.int_fmt_i(sv2v_cast_87CC5(fpu_int_fmt)),
					.vectorial_op_i(1'b0),
					.tag_i(1'b0),
					.in_valid_i(fpu_valid_in),
					.flush_i(reset),
					.result_o(fpu_result[i * 32+:32]),
					.status_o(fpu_status[i * 5+:5]),
					.out_ready_i(fpu_ready_out)
				);
			end
		end
	endgenerate
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:193:5
	assign fpu_valid_in = valid_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:194:5
	assign ready_in = fpu_ready_in;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:196:5
	wire [TAGW:1] sv2v_tmp_14562;
	assign sv2v_tmp_14562 = tag_in;
	always @(*) fpu_tag_in = sv2v_tmp_14562;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:197:5
	assign tag_out = fpu_tag_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:199:5
	assign result = fpu_result;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:201:5
	assign has_fflags = fpu_has_fflags_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:202:5
	assign fflags = fpu_status;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:204:5
	assign valid_out = fpu_valid_out;
	// Trace: ../../rtl/fp_cores/VX_fpu_fpnew.sv:205:5
	assign fpu_ready_out = ready_out;
endmodule
// removed package "ahb_pkg"
module fpnew_cast_multi_35196_62023 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// removed localparam type TagType_TagType_TagType_TagType_TAGW_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:18:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:20:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:21:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:22:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:23:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:25:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:306:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:307:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:310:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:86:45
		input reg [1:0] ifmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:87:5
		case (ifmt)
			sv2v_cast_87CC5(0): fpnew_pkg_int_width = 8;
			sv2v_cast_87CC5(1): fpnew_pkg_int_width = 16;
			sv2v_cast_87CC5(2): fpnew_pkg_int_width = 32;
			sv2v_cast_87CC5(3): fpnew_pkg_int_width = 64;
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:94:9
				$fatal(1, "Invalid INT format supplied");
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:98:9
				fpnew_pkg_int_width = sv2v_cast_87CC5(0);
			end
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:353:49
		input reg [0:3] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:354:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:5
			begin : sv2v_autoblock_2
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:10
				reg signed [31:0] ifmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:356:7
						if (cfg[ifmt])
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:356:22
							res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)));
					end
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_maximum(fpnew_pkg_max_fp_width(FpFmtConfig), fpnew_pkg_max_int_width(IntFmtConfig));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:27:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:29:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:30:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:32:3
	input wire [WIDTH - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:33:3
	input wire [4:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:34:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:35:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:36:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:37:3
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:38:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:39:3
	input wire [1:0] int_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:40:3
	input wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:41:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:43:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:44:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:45:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:47:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:48:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:49:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:50:3
	output wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:51:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:53:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:54:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:56:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:62:3
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:63:3
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:65:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:338:49
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:339:5
		reg [63:0] res;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:340:5
			res = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:5
			begin : sv2v_autoblock_3
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:10
				reg [31:0] fmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:343:9
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt))));
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:344:9
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:67:3
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:68:3
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:69:3
	localparam [31:0] SUPER_BIAS = (2 ** (SUPER_EXP_BITS - 1)) - 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:72:3
	localparam [31:0] INT_MAN_WIDTH = fpnew_pkg_maximum(SUPER_MAN_BITS + 1, MAX_INT_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:74:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(INT_MAN_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:77:3
	localparam [31:0] INT_EXP_WIDTH = fpnew_pkg_maximum($clog2(MAX_INT_WIDTH), fpnew_pkg_maximum(SUPER_EXP_BITS, $clog2(SUPER_BIAS + SUPER_MAN_BITS))) + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:80:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:85:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:90:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:100:3
	wire [WIDTH - 1:0] operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:101:3
	wire [4:0] is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:102:3
	wire op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:103:3
	wire [2:0] src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:104:3
	wire [2:0] dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:105:3
	wire [1:0] int_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:108:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * WIDTH) + ((NUM_INP_REGS * WIDTH) - 1) : ((NUM_INP_REGS + 1) * WIDTH) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * WIDTH : 0)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:109:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)] inp_pipe_is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:110:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:111:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:112:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:113:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:114:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:115:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] inp_pipe_int_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:116:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:117:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:118:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:120:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:123:3
	wire [WIDTH * 1:1] sv2v_tmp_6E45B;
	assign sv2v_tmp_6E45B = operands_i;
	always @(*) inp_pipe_operands_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6E45B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:124:3
	wire [5:1] sv2v_tmp_C47E1;
	assign sv2v_tmp_C47E1 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS] = sv2v_tmp_C47E1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:125:3
	wire [3:1] sv2v_tmp_45ED9;
	assign sv2v_tmp_45ED9 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_45ED9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:126:3
	wire [4:1] sv2v_tmp_AD1FB;
	assign sv2v_tmp_AD1FB = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_AD1FB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:127:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:128:3
	wire [3:1] sv2v_tmp_CB295;
	assign sv2v_tmp_CB295 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_CB295;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:129:3
	wire [3:1] sv2v_tmp_6AF63;
	assign sv2v_tmp_6AF63 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_6AF63;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:130:3
	wire [2:1] sv2v_tmp_CA55F;
	assign sv2v_tmp_CA55F = int_fmt_i;
	always @(*) inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_CA55F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:131:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_BF46E;
	assign sv2v_tmp_BF46E = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_BF46E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:132:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_929AB;
	assign sv2v_tmp_929AB = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_929AB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:133:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:135:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:137:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] sv2v_cast_5B742;
		input reg [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] inp;
		sv2v_cast_5B742 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:139:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:143:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:145:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:145:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:145:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:145:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:147:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:149:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:149:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:149:183
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:149:291
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * WIDTH+:WIDTH] : inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:150:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:150:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:150:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:150:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS+:NUM_FORMATS] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:151:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:151:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:151:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:151:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:152:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:152:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:152:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:152:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:153:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:153:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:153:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:153:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:154:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:154:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:154:207
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:154:315
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:155:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:155:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:155:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:155:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:156:96
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:156:152
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:156:208
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_87CC5(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:156:316
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= (reg_ena ? inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] : inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:157:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:157:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:157:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:157:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:158:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:158:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:158:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:158:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:161:3
	assign operands_q = inp_pipe_operands_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:162:3
	assign is_boxed_q = inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:163:3
	assign op_mod_q = inp_pipe_op_mod_q[NUM_INP_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:164:3
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:165:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:166:3
	assign int_fmt_q = inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:171:3
	wire src_is_int;
	wire dst_is_int;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:173:3
	assign src_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(12);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:174:3
	assign dst_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(11);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:176:3
	wire [INT_MAN_WIDTH - 1:0] encoded_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:178:3
	wire [4:0] fmt_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:179:3
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:180:3
	wire [(NUM_FORMATS * INT_MAN_WIDTH) - 1:0] fmt_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:181:3
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_shift_compensation;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:183:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [39:0] info;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:185:3
	reg [(NUM_INT_FORMATS * INT_MAN_WIDTH) - 1:0] ifmt_input_val;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:186:3
	wire int_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:187:3
	wire [INT_MAN_WIDTH - 1:0] int_value;
	wire [INT_MAN_WIDTH - 1:0] int_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:190:3
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [0:0] sv2v_cast_1_signed;
		input reg signed [0:0] inp;
		sv2v_cast_1_signed = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : fmt_init_inputs
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:192:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:193:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:194:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:198:7
				fpnew_classifier #(
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.NumOperands(1)
				) i_fpnew_classifier(
					.operands_i(operands_q[FP_WIDTH - 1:0]),
					.is_boxed_i(is_boxed_q[fmt]),
					.info_o(info[fmt * 8+:8])
				);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:207:7
				assign fmt_sign[fmt] = operands_q[FP_WIDTH - 1];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:208:7
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed({1'b0, operands_q[MAN_BITS+:EXP_BITS]});
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:209:7
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {info[(fmt * 8) + 7], operands_q[MAN_BITS - 1:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:211:7
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed((INT_MAN_WIDTH - 1) - MAN_BITS);
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:213:7
				assign info[fmt * 8+:8] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:214:7
				assign fmt_sign[fmt] = fpnew_pkg_DONT_CARE;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:215:7
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:216:7
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:217:7
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:222:3
	genvar ifmt;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	generate
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_sign_extend_int
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:224:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:227:7
				always @(*) begin : sign_ext_input
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:229:9
					ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {sv2v_cast_1(operands_q[INT_WIDTH - 1] & ~op_mod_q)}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:230:9
					ifmt_input_val[(ifmt * INT_MAN_WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = operands_q[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:233:7
				wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_5B946;
				assign sv2v_tmp_5B946 = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_5B946;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:238:3
	assign int_value = ifmt_input_val[int_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:239:3
	assign int_sign = int_value[INT_MAN_WIDTH - 1] & ~op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:240:3
	assign int_mantissa = (int_sign ? $unsigned(-int_value) : int_value);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:243:3
	assign encoded_mant = (src_is_int ? int_mantissa : fmt_mantissa[src_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:248:3
	wire signed [INT_EXP_WIDTH - 1:0] src_bias;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:249:3
	wire signed [INT_EXP_WIDTH - 1:0] src_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:250:3
	wire signed [INT_EXP_WIDTH - 1:0] src_subnormal;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:251:3
	wire signed [INT_EXP_WIDTH - 1:0] src_offset;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:253:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:334:40
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:335:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	assign src_bias = $signed(fpnew_pkg_bias(src_fmt_q));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:254:3
	assign src_exp = fmt_exponent[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:255:3
	assign src_subnormal = $signed({1'b0, info[(src_fmt_q * 8) + 6]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:256:3
	assign src_offset = fmt_shift_compensation[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:258:3
	wire input_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:259:3
	wire signed [INT_EXP_WIDTH - 1:0] input_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:260:3
	wire [INT_MAN_WIDTH - 1:0] input_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:261:3
	wire mant_is_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:263:3
	wire signed [INT_EXP_WIDTH - 1:0] fp_input_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:264:3
	wire signed [INT_EXP_WIDTH - 1:0] int_input_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:267:3
	wire [LZC_RESULT_WIDTH - 1:0] renorm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:268:3
	wire [LZC_RESULT_WIDTH:0] renorm_shamt_sgn;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:271:3
	lzc #(
		.WIDTH(INT_MAN_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(encoded_mant),
		.cnt_o(renorm_shamt),
		.empty_o(mant_is_zero)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:279:3
	assign renorm_shamt_sgn = $signed({1'b0, renorm_shamt});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:282:3
	assign input_sign = (src_is_int ? int_sign : fmt_sign[src_fmt_q]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:284:3
	assign input_mant = encoded_mant << renorm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:286:3
	assign fp_input_exp = $signed((((src_exp + src_subnormal) - src_bias) - renorm_shamt_sgn) + src_offset);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:288:3
	assign int_input_exp = $signed((INT_MAN_WIDTH - 1) - renorm_shamt_sgn);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:290:3
	assign input_exp = (src_is_int ? int_input_exp : fp_input_exp);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:292:3
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:295:3
	assign destination_exp = input_exp + $signed(fpnew_pkg_bias(dst_fmt_q));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:301:3
	wire input_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:302:3
	wire signed [INT_EXP_WIDTH - 1:0] input_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:303:3
	wire [INT_MAN_WIDTH - 1:0] input_mant_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:304:3
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:305:3
	wire src_is_int_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:306:3
	wire dst_is_int_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:307:3
	wire [7:0] info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:308:3
	wire mant_is_zero_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:309:3
	wire op_mod_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:310:3
	wire [2:0] rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:311:3
	wire [2:0] src_fmt_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:312:3
	wire [2:0] dst_fmt_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:313:3
	wire [1:0] int_fmt_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:317:3
	reg [0:NUM_MID_REGS] mid_pipe_input_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:318:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_input_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:319:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_MAN_WIDTH) + ((NUM_MID_REGS * INT_MAN_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_MAN_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_MAN_WIDTH : 0)] mid_pipe_input_mant_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:320:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_dest_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:321:3
	reg [0:NUM_MID_REGS] mid_pipe_src_is_int_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:322:3
	reg [0:NUM_MID_REGS] mid_pipe_dst_is_int_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:323:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 8) + ((NUM_MID_REGS * 8) - 1) : ((NUM_MID_REGS + 1) * 8) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 8 : 0)] mid_pipe_info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:324:3
	reg [0:NUM_MID_REGS] mid_pipe_mant_zero_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:325:3
	reg [0:NUM_MID_REGS] mid_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:326:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:327:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:328:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:329:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] mid_pipe_int_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:330:3
	reg [(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_MID_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_MID_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_MID_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_MID_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] mid_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:331:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:332:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:334:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:337:3
	wire [1:1] sv2v_tmp_3DFAC;
	assign sv2v_tmp_3DFAC = input_sign;
	always @(*) mid_pipe_input_sign_q[0] = sv2v_tmp_3DFAC;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:338:3
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_9AB08;
	assign sv2v_tmp_9AB08 = input_exp;
	always @(*) mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_9AB08;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:339:3
	wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_3BE44;
	assign sv2v_tmp_3BE44 = input_mant;
	always @(*) mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_3BE44;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:340:3
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_F626F;
	assign sv2v_tmp_F626F = destination_exp;
	always @(*) mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_F626F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:341:3
	wire [1:1] sv2v_tmp_3D9F8;
	assign sv2v_tmp_3D9F8 = src_is_int;
	always @(*) mid_pipe_src_is_int_q[0] = sv2v_tmp_3D9F8;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:342:3
	wire [1:1] sv2v_tmp_4E95C;
	assign sv2v_tmp_4E95C = dst_is_int;
	always @(*) mid_pipe_dst_is_int_q[0] = sv2v_tmp_4E95C;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:343:3
	wire [8:1] sv2v_tmp_48E57;
	assign sv2v_tmp_48E57 = info[src_fmt_q * 8+:8];
	always @(*) mid_pipe_info_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 8+:8] = sv2v_tmp_48E57;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:344:3
	wire [1:1] sv2v_tmp_4351A;
	assign sv2v_tmp_4351A = mant_is_zero;
	always @(*) mid_pipe_mant_zero_q[0] = sv2v_tmp_4351A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:345:3
	wire [1:1] sv2v_tmp_88AB6;
	assign sv2v_tmp_88AB6 = op_mod_q;
	always @(*) mid_pipe_op_mod_q[0] = sv2v_tmp_88AB6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:346:3
	wire [3:1] sv2v_tmp_32E16;
	assign sv2v_tmp_32E16 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_32E16;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:347:3
	wire [3:1] sv2v_tmp_DE9EA;
	assign sv2v_tmp_DE9EA = src_fmt_q;
	always @(*) mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_DE9EA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:348:3
	wire [3:1] sv2v_tmp_FC1E4;
	assign sv2v_tmp_FC1E4 = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_FC1E4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:349:3
	wire [2:1] sv2v_tmp_2AE08;
	assign sv2v_tmp_2AE08 = int_fmt_q;
	always @(*) mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_2AE08;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:350:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_B21BC;
	assign sv2v_tmp_B21BC = inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	always @(*) mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_B21BC;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:351:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_BB372;
	assign sv2v_tmp_BB372 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_BB372;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:352:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:354:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:357:3
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:359:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:363:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:365:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:365:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:365:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:365:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:367:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:369:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:369:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:369:187
					mid_pipe_input_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:369:295
					mid_pipe_input_sign_q[i + 1] <= (reg_ena ? mid_pipe_input_sign_q[i] : mid_pipe_input_sign_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:370:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:370:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:370:187
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:370:295
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= (reg_ena ? mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH] : mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:371:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:371:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:371:187
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:371:295
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= (reg_ena ? mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_MAN_WIDTH+:INT_MAN_WIDTH] : mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:372:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:372:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:372:187
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:372:295
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= (reg_ena ? mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH] : mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:373:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:373:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:373:187
					mid_pipe_src_is_int_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:373:295
					mid_pipe_src_is_int_q[i + 1] <= (reg_ena ? mid_pipe_src_is_int_q[i] : mid_pipe_src_is_int_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:374:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:374:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:374:187
					mid_pipe_dst_is_int_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:374:295
					mid_pipe_dst_is_int_q[i + 1] <= (reg_ena ? mid_pipe_dst_is_int_q[i] : mid_pipe_dst_is_int_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:375:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:375:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:375:187
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:375:295
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= (reg_ena ? mid_pipe_info_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 8+:8] : mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:376:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:376:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:376:187
					mid_pipe_mant_zero_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:376:295
					mid_pipe_mant_zero_q[i + 1] <= (reg_ena ? mid_pipe_mant_zero_q[i] : mid_pipe_mant_zero_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:377:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:377:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:377:187
					mid_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:377:295
					mid_pipe_op_mod_q[i + 1] <= (reg_ena ? mid_pipe_op_mod_q[i] : mid_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:378:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:378:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:378:199
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:378:307
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:379:99
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:379:155
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:379:211
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:379:319
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:380:99
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:380:155
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:380:211
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:380:319
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:381:100
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:381:156
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:381:212
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_87CC5(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:381:320
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= (reg_ena ? mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] : mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:382:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:382:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:382:197
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:382:305
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:383:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:383:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:383:197
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:383:305
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:386:3
	assign input_sign_q = mid_pipe_input_sign_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:387:3
	assign input_exp_q = mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:388:3
	assign input_mant_q = mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:389:3
	assign destination_exp_q = mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:390:3
	assign src_is_int_q = mid_pipe_src_is_int_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:391:3
	assign dst_is_int_q = mid_pipe_dst_is_int_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:392:3
	assign info_q = mid_pipe_info_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 8+:8];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:393:3
	assign mant_is_zero_q = mid_pipe_mant_zero_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:394:3
	assign op_mod_q2 = mid_pipe_op_mod_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:395:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:396:3
	assign src_fmt_q2 = mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:397:3
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:398:3
	assign int_fmt_q2 = mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:403:3
	reg [INT_EXP_WIDTH - 1:0] final_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:405:3
	reg [2 * INT_MAN_WIDTH:0] preshift_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:406:3
	wire [2 * INT_MAN_WIDTH:0] destination_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:407:3
	wire [SUPER_MAN_BITS - 1:0] final_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:408:3
	wire [MAX_INT_WIDTH - 1:0] final_int;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:410:3
	reg [$clog2(INT_MAN_WIDTH + 1) - 1:0] denorm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:412:3
	wire [1:0] fp_round_sticky_bits;
	wire [1:0] int_round_sticky_bits;
	wire [1:0] round_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:413:3
	reg of_before_round;
	reg uf_before_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:417:3
	always @(*) begin : cast_value
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:419:5
		final_exp = $unsigned(destination_exp_q);
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:420:5
		preshift_mant = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:421:5
		denorm_shamt = SUPER_MAN_BITS - fpnew_pkg_man_bits(dst_fmt_q2);
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:422:5
		of_before_round = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:423:5
		uf_before_round = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:426:5
		preshift_mant = input_mant_q << (INT_MAN_WIDTH + 1);
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:429:5
		if (dst_is_int_q) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:431:7
			denorm_shamt = $unsigned((MAX_INT_WIDTH - 1) - input_exp_q);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:433:7
			if (input_exp_q >= $signed((fpnew_pkg_int_width(int_fmt_q2) - 1) + op_mod_q2)) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:434:9
				denorm_shamt = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:435:9
				of_before_round = 1'b1;
			end
			else if (input_exp_q < -1) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:438:9
				denorm_shamt = MAX_INT_WIDTH + 1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:439:9
				uf_before_round = 1'b1;
			end
		end
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:444:7
			if ((destination_exp_q >= ($signed(2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1)) || (~src_is_int_q && info_q[4])) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:446:9
				final_exp = $unsigned((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 2);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:447:9
				preshift_mant = 1'sb1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:448:9
				of_before_round = 1'b1;
			end
			else if ((destination_exp_q < 1) && (destination_exp_q >= -$signed(fpnew_pkg_man_bits(dst_fmt_q2)))) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:452:9
				final_exp = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:453:9
				denorm_shamt = $unsigned((denorm_shamt + 1) - destination_exp_q);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:454:9
				uf_before_round = 1'b1;
			end
			else if (destination_exp_q < -$signed(fpnew_pkg_man_bits(dst_fmt_q2))) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:457:9
				final_exp = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:458:9
				denorm_shamt = $unsigned((denorm_shamt + 2) + fpnew_pkg_man_bits(dst_fmt_q2));
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:459:9
				uf_before_round = 1'b1;
			end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:464:3
	localparam NUM_FP_STICKY = ((2 * INT_MAN_WIDTH) - SUPER_MAN_BITS) - 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:465:3
	localparam NUM_INT_STICKY = (2 * INT_MAN_WIDTH) - MAX_INT_WIDTH;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:468:3
	assign destination_mant = preshift_mant >> denorm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:470:3
	assign {final_mant, fp_round_sticky_bits[1]} = destination_mant[(2 * INT_MAN_WIDTH) - 1-:SUPER_MAN_BITS + 1];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:472:3
	assign {final_int, int_round_sticky_bits[1]} = destination_mant[2 * INT_MAN_WIDTH-:MAX_INT_WIDTH + 1];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:474:3
	assign fp_round_sticky_bits[0] = |{destination_mant[NUM_FP_STICKY - 1:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:475:3
	assign int_round_sticky_bits[0] = |{destination_mant[NUM_INT_STICKY - 1:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:478:3
	assign round_sticky_bits = (dst_is_int_q ? int_round_sticky_bits : fp_round_sticky_bits);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:483:3
	wire [WIDTH - 1:0] pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:484:3
	wire of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:485:3
	wire uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:487:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:488:3
	reg [4:0] fmt_of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:489:3
	reg [4:0] fmt_uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:491:3
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:493:3
	wire rounded_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:494:3
	wire [WIDTH - 1:0] rounded_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:495:3
	wire result_true_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:497:3
	wire [WIDTH - 1:0] rounded_int_res;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:498:3
	wire rounded_int_res_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:502:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_res_assemble
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:504:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:505:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:508:7
				always @(*) begin : assemble_result
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:509:9
					fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = {final_exp[EXP_BITS - 1:0], final_mant[MAN_BITS - 1:0]};
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:512:7
				wire [WIDTH * 1:1] sv2v_tmp_C33E0;
				assign sv2v_tmp_C33E0 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = sv2v_tmp_C33E0;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:517:3
	generate
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_int_res_sign_ext
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:519:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:522:7
				always @(*) begin : assemble_result
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:524:9
					ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = {WIDTH {final_int[INT_WIDTH - 1]}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:525:9
					ifmt_pre_round_abs[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = final_int[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:528:7
				wire [WIDTH * 1:1] sv2v_tmp_F6FA8;
				assign sv2v_tmp_F6FA8 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = sv2v_tmp_F6FA8;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:533:3
	assign pre_round_abs = (dst_is_int_q ? ifmt_pre_round_abs[int_fmt_q2 * WIDTH+:WIDTH] : fmt_pre_round_abs[dst_fmt_q2 * WIDTH+:WIDTH]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:535:3
	fpnew_rounding #(.AbsWidth(WIDTH)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(input_sign_q),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(1'b0),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_true_zero)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:548:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:551:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_sign_inject
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:553:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:554:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:555:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:558:7
				always @(*) begin : post_process
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:560:9
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:561:9
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:564:9
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:565:9
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = (src_is_int_q & mant_is_zero_q ? {FP_WIDTH * 1 {1'sb0}} : {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]});
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:570:7
				wire [1:1] sv2v_tmp_4A747;
				assign sv2v_tmp_4A747 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4A747;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:571:7
				wire [1:1] sv2v_tmp_90681;
				assign sv2v_tmp_90681 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_90681;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:572:7
				wire [WIDTH * 1:1] sv2v_tmp_649FB;
				assign sv2v_tmp_649FB = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_649FB;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:577:3
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:578:3
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:581:3
	assign rounded_int_res = (rounded_sign ? $unsigned(-rounded_abs) : rounded_abs);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:582:3
	assign rounded_int_res_zero = rounded_int_res == {WIDTH {1'sb0}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:587:3
	wire [WIDTH - 1:0] fp_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:588:3
	wire [4:0] fp_special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:589:3
	wire fp_result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:591:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:594:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_special_results
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:596:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:597:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:598:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:600:5
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:601:5
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:604:7
				always @(*) begin : special_results
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:605:9
					reg [FP_WIDTH - 1:0] special_res;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:606:9
					special_res = (info_q[5] ? input_sign_q << (FP_WIDTH - 1) : {1'b0, QNAN_EXPONENT, QNAN_MANTISSA});
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:611:9
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:612:9
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:615:7
				wire [WIDTH * 1:1] sv2v_tmp_B718F;
				assign sv2v_tmp_B718F = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_B718F;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:620:3
	assign fp_result_is_special = ~src_is_int_q & ((info_q[5] | info_q[3]) | ~info_q[0]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:625:3
	assign fp_special_status = {info_q[2], 4'b0000};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:628:3
	assign fp_special_result = fmt_special_result[dst_fmt_q2 * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:633:3
	wire [WIDTH - 1:0] int_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:634:3
	wire [4:0] int_special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:635:3
	wire int_result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:637:3
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:640:3
	generate
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_special_results_int
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:642:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:645:7
				always @(*) begin : special_results
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:646:9
					reg [INT_WIDTH - 1:0] special_res;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:649:9
					special_res[INT_WIDTH - 2:0] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:650:9
					special_res[INT_WIDTH - 1] = op_mod_q2;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:653:9
					if (input_sign_q && !info_q[3])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:654:11
						special_res = ~special_res;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:657:9
					ifmt_special_result[ifmt * WIDTH+:WIDTH] = {WIDTH {special_res[INT_WIDTH - 1]}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:658:9
					ifmt_special_result[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:661:7
				wire [WIDTH * 1:1] sv2v_tmp_99B6D;
				assign sv2v_tmp_99B6D = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_special_result[ifmt * WIDTH+:WIDTH] = sv2v_tmp_99B6D;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:666:3
	assign int_result_is_special = (((info_q[3] | info_q[4]) | of_before_round) | ~info_q[0]) | ((input_sign_q & op_mod_q2) & ~rounded_int_res_zero);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:671:3
	assign int_special_status = 5'b10000;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:674:3
	assign int_special_result = ifmt_special_result[int_fmt_q2 * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:679:3
	wire [4:0] int_regular_status;
	wire [4:0] fp_regular_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:681:3
	wire [WIDTH - 1:0] fp_result;
	wire [WIDTH - 1:0] int_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:682:3
	wire [4:0] fp_status;
	wire [4:0] int_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:684:3
	assign fp_regular_status[4] = src_is_int_q & (of_before_round | of_after_round);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:685:3
	assign fp_regular_status[3] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:686:3
	assign fp_regular_status[2] = ~src_is_int_q & (~info_q[4] & (of_before_round | of_after_round));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:687:3
	assign fp_regular_status[1] = uf_after_round & fp_regular_status[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:688:3
	assign fp_regular_status[0] = (src_is_int_q ? |fp_round_sticky_bits : |fp_round_sticky_bits | (~info_q[4] & (of_before_round | of_after_round)));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:690:3
	assign int_regular_status = {4'b0000, |int_round_sticky_bits};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:692:3
	assign fp_result = (fp_result_is_special ? fp_special_result : fmt_result[dst_fmt_q2 * WIDTH+:WIDTH]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:693:3
	assign fp_status = (fp_result_is_special ? fp_special_status : fp_regular_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:694:3
	assign int_result = (int_result_is_special ? int_special_result : rounded_int_res);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:695:3
	assign int_status = (int_result_is_special ? int_special_status : int_regular_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:698:3
	wire [WIDTH - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:699:3
	wire [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:700:3
	wire extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:703:3
	assign result_d = (dst_is_int_q ? int_result : fp_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:704:3
	assign status_d = (dst_is_int_q ? int_status : fp_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:707:3
	assign extension_bit = (dst_is_int_q ? int_result[WIDTH - 1] : 1'b1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:713:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:714:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:715:3
	reg [0:NUM_OUT_REGS] out_pipe_ext_bit_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:716:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:717:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:718:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:720:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:723:3
	wire [WIDTH * 1:1] sv2v_tmp_4086F;
	assign sv2v_tmp_4086F = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_4086F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:724:3
	wire [5:1] sv2v_tmp_B7C45;
	assign sv2v_tmp_B7C45 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_B7C45;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:725:3
	wire [1:1] sv2v_tmp_8F736;
	assign sv2v_tmp_8F736 = extension_bit;
	always @(*) out_pipe_ext_bit_q[0] = sv2v_tmp_8F736;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:726:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_F9425;
	assign sv2v_tmp_F9425 = mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_F9425;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:727:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_3D161;
	assign sv2v_tmp_3D161 = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_3D161;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:728:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:730:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:732:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:734:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:738:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:740:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:740:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:740:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:740:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:742:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:744:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:744:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:744:181
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:744:289
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:745:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:745:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:745:181
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:745:289
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:746:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:746:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:746:181
					out_pipe_ext_bit_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:746:289
					out_pipe_ext_bit_q[i + 1] <= (reg_ena ? out_pipe_ext_bit_q[i] : out_pipe_ext_bit_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:747:79
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:747:135
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:747:191
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:747:299
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:748:79
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:748:135
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:748:191
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:748:299
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:751:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:753:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:754:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:755:3
	assign extension_bit_o = out_pipe_ext_bit_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:756:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:757:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:758:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:759:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_cast_multi_7061A_0B31A (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:18:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:20:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:21:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:22:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:23:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:25:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:306:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:307:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:310:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:86:45
		input reg [1:0] ifmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:87:5
		case (ifmt)
			sv2v_cast_87CC5(0): fpnew_pkg_int_width = 8;
			sv2v_cast_87CC5(1): fpnew_pkg_int_width = 16;
			sv2v_cast_87CC5(2): fpnew_pkg_int_width = 32;
			sv2v_cast_87CC5(3): fpnew_pkg_int_width = 64;
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:94:9
				$fatal(1, "Invalid INT format supplied");
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:98:9
				fpnew_pkg_int_width = sv2v_cast_87CC5(0);
			end
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:353:49
		input reg [0:3] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:354:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:5
			begin : sv2v_autoblock_2
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:10
				reg signed [31:0] ifmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:356:7
						if (cfg[ifmt])
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:356:22
							res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)));
					end
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_maximum(fpnew_pkg_max_fp_width(FpFmtConfig), fpnew_pkg_max_int_width(IntFmtConfig));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:27:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:29:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:30:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:32:3
	input wire [WIDTH - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:33:3
	input wire [4:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:34:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:35:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:36:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:37:3
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:38:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:39:3
	input wire [1:0] int_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:40:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:41:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:43:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:44:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:45:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:47:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:48:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:49:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:50:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:51:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:53:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:54:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:56:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:62:3
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:63:3
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:65:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:338:49
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:339:5
		reg [63:0] res;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:340:5
			res = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:5
			begin : sv2v_autoblock_3
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:10
				reg [31:0] fmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:343:9
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt))));
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:344:9
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:67:3
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:68:3
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:69:3
	localparam [31:0] SUPER_BIAS = (2 ** (SUPER_EXP_BITS - 1)) - 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:72:3
	localparam [31:0] INT_MAN_WIDTH = fpnew_pkg_maximum(SUPER_MAN_BITS + 1, MAX_INT_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:74:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(INT_MAN_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:77:3
	localparam [31:0] INT_EXP_WIDTH = fpnew_pkg_maximum($clog2(MAX_INT_WIDTH), fpnew_pkg_maximum(SUPER_EXP_BITS, $clog2(SUPER_BIAS + SUPER_MAN_BITS))) + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:80:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:85:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:90:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:100:3
	wire [WIDTH - 1:0] operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:101:3
	wire [4:0] is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:102:3
	wire op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:103:3
	wire [2:0] src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:104:3
	wire [2:0] dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:105:3
	wire [1:0] int_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:108:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * WIDTH) + ((NUM_INP_REGS * WIDTH) - 1) : ((NUM_INP_REGS + 1) * WIDTH) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * WIDTH : 0)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:109:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)] inp_pipe_is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:110:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:111:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:112:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:113:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:114:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:115:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] inp_pipe_int_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:116:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:117:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:118:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:120:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:123:3
	wire [WIDTH * 1:1] sv2v_tmp_6E45B;
	assign sv2v_tmp_6E45B = operands_i;
	always @(*) inp_pipe_operands_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6E45B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:124:3
	wire [5:1] sv2v_tmp_C47E1;
	assign sv2v_tmp_C47E1 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS] = sv2v_tmp_C47E1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:125:3
	wire [3:1] sv2v_tmp_45ED9;
	assign sv2v_tmp_45ED9 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_45ED9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:126:3
	wire [4:1] sv2v_tmp_AD1FB;
	assign sv2v_tmp_AD1FB = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_AD1FB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:127:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:128:3
	wire [3:1] sv2v_tmp_CB295;
	assign sv2v_tmp_CB295 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_CB295;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:129:3
	wire [3:1] sv2v_tmp_6AF63;
	assign sv2v_tmp_6AF63 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_6AF63;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:130:3
	wire [2:1] sv2v_tmp_CA55F;
	assign sv2v_tmp_CA55F = int_fmt_i;
	always @(*) inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_CA55F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:131:3
	wire [1:1] sv2v_tmp_76699;
	assign sv2v_tmp_76699 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_76699;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:132:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_90A49;
	assign sv2v_tmp_90A49 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_90A49;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:133:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:135:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:137:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:139:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:143:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:145:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:145:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:145:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:145:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:147:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:149:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:149:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:149:183
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:149:291
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * WIDTH+:WIDTH] : inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:150:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:150:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:150:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:150:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS+:NUM_FORMATS] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:151:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:151:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:151:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:151:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:152:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:152:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:152:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:152:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:153:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:153:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:153:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:153:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:154:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:154:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:154:207
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:154:315
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:155:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:155:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:155:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:155:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:156:96
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:156:152
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:156:208
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_87CC5(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:156:316
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= (reg_ena ? inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] : inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:157:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:157:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:157:193
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:157:301
					inp_pipe_tag_q[i + 1] <= (reg_ena ? inp_pipe_tag_q[i] : inp_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:158:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:158:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:158:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:158:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:161:3
	assign operands_q = inp_pipe_operands_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:162:3
	assign is_boxed_q = inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:163:3
	assign op_mod_q = inp_pipe_op_mod_q[NUM_INP_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:164:3
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:165:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:166:3
	assign int_fmt_q = inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:171:3
	wire src_is_int;
	wire dst_is_int;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:173:3
	assign src_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(12);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:174:3
	assign dst_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(11);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:176:3
	wire [INT_MAN_WIDTH - 1:0] encoded_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:178:3
	wire [4:0] fmt_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:179:3
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:180:3
	wire [(NUM_FORMATS * INT_MAN_WIDTH) - 1:0] fmt_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:181:3
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_shift_compensation;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:183:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [39:0] info;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:185:3
	reg [(NUM_INT_FORMATS * INT_MAN_WIDTH) - 1:0] ifmt_input_val;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:186:3
	wire int_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:187:3
	wire [INT_MAN_WIDTH - 1:0] int_value;
	wire [INT_MAN_WIDTH - 1:0] int_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:190:3
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [0:0] sv2v_cast_1_signed;
		input reg signed [0:0] inp;
		sv2v_cast_1_signed = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : fmt_init_inputs
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:192:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:193:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:194:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:198:7
				fpnew_classifier #(
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.NumOperands(1)
				) i_fpnew_classifier(
					.operands_i(operands_q[FP_WIDTH - 1:0]),
					.is_boxed_i(is_boxed_q[fmt]),
					.info_o(info[fmt * 8+:8])
				);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:207:7
				assign fmt_sign[fmt] = operands_q[FP_WIDTH - 1];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:208:7
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed({1'b0, operands_q[MAN_BITS+:EXP_BITS]});
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:209:7
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {info[(fmt * 8) + 7], operands_q[MAN_BITS - 1:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:211:7
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed((INT_MAN_WIDTH - 1) - MAN_BITS);
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:213:7
				assign info[fmt * 8+:8] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:214:7
				assign fmt_sign[fmt] = fpnew_pkg_DONT_CARE;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:215:7
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:216:7
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:217:7
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:222:3
	genvar ifmt;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	generate
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_sign_extend_int
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:224:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:227:7
				always @(*) begin : sign_ext_input
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:229:9
					ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {sv2v_cast_1(operands_q[INT_WIDTH - 1] & ~op_mod_q)}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:230:9
					ifmt_input_val[(ifmt * INT_MAN_WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = operands_q[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:233:7
				wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_5B946;
				assign sv2v_tmp_5B946 = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_5B946;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:238:3
	assign int_value = ifmt_input_val[int_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:239:3
	assign int_sign = int_value[INT_MAN_WIDTH - 1] & ~op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:240:3
	assign int_mantissa = (int_sign ? $unsigned(-int_value) : int_value);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:243:3
	assign encoded_mant = (src_is_int ? int_mantissa : fmt_mantissa[src_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:248:3
	wire signed [INT_EXP_WIDTH - 1:0] src_bias;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:249:3
	wire signed [INT_EXP_WIDTH - 1:0] src_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:250:3
	wire signed [INT_EXP_WIDTH - 1:0] src_subnormal;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:251:3
	wire signed [INT_EXP_WIDTH - 1:0] src_offset;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:253:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:334:40
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:335:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	assign src_bias = $signed(fpnew_pkg_bias(src_fmt_q));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:254:3
	assign src_exp = fmt_exponent[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:255:3
	assign src_subnormal = $signed({1'b0, info[(src_fmt_q * 8) + 6]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:256:3
	assign src_offset = fmt_shift_compensation[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:258:3
	wire input_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:259:3
	wire signed [INT_EXP_WIDTH - 1:0] input_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:260:3
	wire [INT_MAN_WIDTH - 1:0] input_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:261:3
	wire mant_is_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:263:3
	wire signed [INT_EXP_WIDTH - 1:0] fp_input_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:264:3
	wire signed [INT_EXP_WIDTH - 1:0] int_input_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:267:3
	wire [LZC_RESULT_WIDTH - 1:0] renorm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:268:3
	wire [LZC_RESULT_WIDTH:0] renorm_shamt_sgn;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:271:3
	lzc #(
		.WIDTH(INT_MAN_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(encoded_mant),
		.cnt_o(renorm_shamt),
		.empty_o(mant_is_zero)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:279:3
	assign renorm_shamt_sgn = $signed({1'b0, renorm_shamt});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:282:3
	assign input_sign = (src_is_int ? int_sign : fmt_sign[src_fmt_q]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:284:3
	assign input_mant = encoded_mant << renorm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:286:3
	assign fp_input_exp = $signed((((src_exp + src_subnormal) - src_bias) - renorm_shamt_sgn) + src_offset);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:288:3
	assign int_input_exp = $signed((INT_MAN_WIDTH - 1) - renorm_shamt_sgn);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:290:3
	assign input_exp = (src_is_int ? int_input_exp : fp_input_exp);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:292:3
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:295:3
	assign destination_exp = input_exp + $signed(fpnew_pkg_bias(dst_fmt_q));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:301:3
	wire input_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:302:3
	wire signed [INT_EXP_WIDTH - 1:0] input_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:303:3
	wire [INT_MAN_WIDTH - 1:0] input_mant_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:304:3
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:305:3
	wire src_is_int_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:306:3
	wire dst_is_int_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:307:3
	wire [7:0] info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:308:3
	wire mant_is_zero_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:309:3
	wire op_mod_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:310:3
	wire [2:0] rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:311:3
	wire [2:0] src_fmt_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:312:3
	wire [2:0] dst_fmt_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:313:3
	wire [1:0] int_fmt_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:317:3
	reg [0:NUM_MID_REGS] mid_pipe_input_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:318:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_input_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:319:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_MAN_WIDTH) + ((NUM_MID_REGS * INT_MAN_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_MAN_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_MAN_WIDTH : 0)] mid_pipe_input_mant_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:320:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_dest_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:321:3
	reg [0:NUM_MID_REGS] mid_pipe_src_is_int_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:322:3
	reg [0:NUM_MID_REGS] mid_pipe_dst_is_int_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:323:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 8) + ((NUM_MID_REGS * 8) - 1) : ((NUM_MID_REGS + 1) * 8) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 8 : 0)] mid_pipe_info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:324:3
	reg [0:NUM_MID_REGS] mid_pipe_mant_zero_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:325:3
	reg [0:NUM_MID_REGS] mid_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:326:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:327:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:328:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:329:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] mid_pipe_int_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:330:3
	reg [0:NUM_MID_REGS] mid_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:331:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:332:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:334:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:337:3
	wire [1:1] sv2v_tmp_3DFAC;
	assign sv2v_tmp_3DFAC = input_sign;
	always @(*) mid_pipe_input_sign_q[0] = sv2v_tmp_3DFAC;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:338:3
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_9AB08;
	assign sv2v_tmp_9AB08 = input_exp;
	always @(*) mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_9AB08;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:339:3
	wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_3BE44;
	assign sv2v_tmp_3BE44 = input_mant;
	always @(*) mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_3BE44;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:340:3
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_F626F;
	assign sv2v_tmp_F626F = destination_exp;
	always @(*) mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_F626F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:341:3
	wire [1:1] sv2v_tmp_3D9F8;
	assign sv2v_tmp_3D9F8 = src_is_int;
	always @(*) mid_pipe_src_is_int_q[0] = sv2v_tmp_3D9F8;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:342:3
	wire [1:1] sv2v_tmp_4E95C;
	assign sv2v_tmp_4E95C = dst_is_int;
	always @(*) mid_pipe_dst_is_int_q[0] = sv2v_tmp_4E95C;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:343:3
	wire [8:1] sv2v_tmp_48E57;
	assign sv2v_tmp_48E57 = info[src_fmt_q * 8+:8];
	always @(*) mid_pipe_info_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 8+:8] = sv2v_tmp_48E57;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:344:3
	wire [1:1] sv2v_tmp_4351A;
	assign sv2v_tmp_4351A = mant_is_zero;
	always @(*) mid_pipe_mant_zero_q[0] = sv2v_tmp_4351A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:345:3
	wire [1:1] sv2v_tmp_88AB6;
	assign sv2v_tmp_88AB6 = op_mod_q;
	always @(*) mid_pipe_op_mod_q[0] = sv2v_tmp_88AB6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:346:3
	wire [3:1] sv2v_tmp_32E16;
	assign sv2v_tmp_32E16 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_32E16;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:347:3
	wire [3:1] sv2v_tmp_DE9EA;
	assign sv2v_tmp_DE9EA = src_fmt_q;
	always @(*) mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_DE9EA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:348:3
	wire [3:1] sv2v_tmp_FC1E4;
	assign sv2v_tmp_FC1E4 = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_FC1E4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:349:3
	wire [2:1] sv2v_tmp_2AE08;
	assign sv2v_tmp_2AE08 = int_fmt_q;
	always @(*) mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_2AE08;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:350:3
	wire [1:1] sv2v_tmp_44BCE;
	assign sv2v_tmp_44BCE = inp_pipe_tag_q[NUM_INP_REGS];
	always @(*) mid_pipe_tag_q[0] = sv2v_tmp_44BCE;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:351:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_FBD8C;
	assign sv2v_tmp_FBD8C = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_FBD8C;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:352:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:354:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:357:3
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:359:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:363:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:365:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:365:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:365:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:365:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:367:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:369:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:369:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:369:187
					mid_pipe_input_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:369:295
					mid_pipe_input_sign_q[i + 1] <= (reg_ena ? mid_pipe_input_sign_q[i] : mid_pipe_input_sign_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:370:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:370:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:370:187
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:370:295
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= (reg_ena ? mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH] : mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:371:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:371:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:371:187
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:371:295
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= (reg_ena ? mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_MAN_WIDTH+:INT_MAN_WIDTH] : mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:372:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:372:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:372:187
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:372:295
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= (reg_ena ? mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH] : mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:373:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:373:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:373:187
					mid_pipe_src_is_int_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:373:295
					mid_pipe_src_is_int_q[i + 1] <= (reg_ena ? mid_pipe_src_is_int_q[i] : mid_pipe_src_is_int_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:374:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:374:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:374:187
					mid_pipe_dst_is_int_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:374:295
					mid_pipe_dst_is_int_q[i + 1] <= (reg_ena ? mid_pipe_dst_is_int_q[i] : mid_pipe_dst_is_int_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:375:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:375:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:375:187
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:375:295
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= (reg_ena ? mid_pipe_info_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 8+:8] : mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:376:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:376:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:376:187
					mid_pipe_mant_zero_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:376:295
					mid_pipe_mant_zero_q[i + 1] <= (reg_ena ? mid_pipe_mant_zero_q[i] : mid_pipe_mant_zero_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:377:75
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:377:131
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:377:187
					mid_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:377:295
					mid_pipe_op_mod_q[i + 1] <= (reg_ena ? mid_pipe_op_mod_q[i] : mid_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:378:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:378:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:378:199
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:378:307
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:379:99
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:379:155
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:379:211
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:379:319
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:380:99
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:380:155
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:380:211
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:380:319
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:381:100
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:381:156
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:381:212
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_87CC5(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:381:320
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= (reg_ena ? mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] : mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:382:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:382:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:382:197
					mid_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:382:305
					mid_pipe_tag_q[i + 1] <= (reg_ena ? mid_pipe_tag_q[i] : mid_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:383:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:383:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:383:197
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:383:305
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:386:3
	assign input_sign_q = mid_pipe_input_sign_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:387:3
	assign input_exp_q = mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:388:3
	assign input_mant_q = mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:389:3
	assign destination_exp_q = mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:390:3
	assign src_is_int_q = mid_pipe_src_is_int_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:391:3
	assign dst_is_int_q = mid_pipe_dst_is_int_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:392:3
	assign info_q = mid_pipe_info_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 8+:8];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:393:3
	assign mant_is_zero_q = mid_pipe_mant_zero_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:394:3
	assign op_mod_q2 = mid_pipe_op_mod_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:395:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:396:3
	assign src_fmt_q2 = mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:397:3
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:398:3
	assign int_fmt_q2 = mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:403:3
	reg [INT_EXP_WIDTH - 1:0] final_exp;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:405:3
	reg [2 * INT_MAN_WIDTH:0] preshift_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:406:3
	wire [2 * INT_MAN_WIDTH:0] destination_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:407:3
	wire [SUPER_MAN_BITS - 1:0] final_mant;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:408:3
	wire [MAX_INT_WIDTH - 1:0] final_int;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:410:3
	reg [$clog2(INT_MAN_WIDTH + 1) - 1:0] denorm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:412:3
	wire [1:0] fp_round_sticky_bits;
	wire [1:0] int_round_sticky_bits;
	wire [1:0] round_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:413:3
	reg of_before_round;
	reg uf_before_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:417:3
	always @(*) begin : cast_value
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:419:5
		final_exp = $unsigned(destination_exp_q);
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:420:5
		preshift_mant = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:421:5
		denorm_shamt = SUPER_MAN_BITS - fpnew_pkg_man_bits(dst_fmt_q2);
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:422:5
		of_before_round = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:423:5
		uf_before_round = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:426:5
		preshift_mant = input_mant_q << (INT_MAN_WIDTH + 1);
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:429:5
		if (dst_is_int_q) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:431:7
			denorm_shamt = $unsigned((MAX_INT_WIDTH - 1) - input_exp_q);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:433:7
			if (input_exp_q >= $signed((fpnew_pkg_int_width(int_fmt_q2) - 1) + op_mod_q2)) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:434:9
				denorm_shamt = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:435:9
				of_before_round = 1'b1;
			end
			else if (input_exp_q < -1) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:438:9
				denorm_shamt = MAX_INT_WIDTH + 1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:439:9
				uf_before_round = 1'b1;
			end
		end
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:444:7
			if ((destination_exp_q >= ($signed(2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1)) || (~src_is_int_q && info_q[4])) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:446:9
				final_exp = $unsigned((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 2);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:447:9
				preshift_mant = 1'sb1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:448:9
				of_before_round = 1'b1;
			end
			else if ((destination_exp_q < 1) && (destination_exp_q >= -$signed(fpnew_pkg_man_bits(dst_fmt_q2)))) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:452:9
				final_exp = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:453:9
				denorm_shamt = $unsigned((denorm_shamt + 1) - destination_exp_q);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:454:9
				uf_before_round = 1'b1;
			end
			else if (destination_exp_q < -$signed(fpnew_pkg_man_bits(dst_fmt_q2))) begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:457:9
				final_exp = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:458:9
				denorm_shamt = $unsigned((denorm_shamt + 2) + fpnew_pkg_man_bits(dst_fmt_q2));
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:459:9
				uf_before_round = 1'b1;
			end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:464:3
	localparam NUM_FP_STICKY = ((2 * INT_MAN_WIDTH) - SUPER_MAN_BITS) - 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:465:3
	localparam NUM_INT_STICKY = (2 * INT_MAN_WIDTH) - MAX_INT_WIDTH;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:468:3
	assign destination_mant = preshift_mant >> denorm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:470:3
	assign {final_mant, fp_round_sticky_bits[1]} = destination_mant[(2 * INT_MAN_WIDTH) - 1-:SUPER_MAN_BITS + 1];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:472:3
	assign {final_int, int_round_sticky_bits[1]} = destination_mant[2 * INT_MAN_WIDTH-:MAX_INT_WIDTH + 1];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:474:3
	assign fp_round_sticky_bits[0] = |{destination_mant[NUM_FP_STICKY - 1:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:475:3
	assign int_round_sticky_bits[0] = |{destination_mant[NUM_INT_STICKY - 1:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:478:3
	assign round_sticky_bits = (dst_is_int_q ? int_round_sticky_bits : fp_round_sticky_bits);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:483:3
	wire [WIDTH - 1:0] pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:484:3
	wire of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:485:3
	wire uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:487:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:488:3
	reg [4:0] fmt_of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:489:3
	reg [4:0] fmt_uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:491:3
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:493:3
	wire rounded_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:494:3
	wire [WIDTH - 1:0] rounded_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:495:3
	wire result_true_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:497:3
	wire [WIDTH - 1:0] rounded_int_res;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:498:3
	wire rounded_int_res_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:502:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_res_assemble
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:504:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:505:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:508:7
				always @(*) begin : assemble_result
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:509:9
					fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = {final_exp[EXP_BITS - 1:0], final_mant[MAN_BITS - 1:0]};
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:512:7
				wire [WIDTH * 1:1] sv2v_tmp_C33E0;
				assign sv2v_tmp_C33E0 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = sv2v_tmp_C33E0;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:517:3
	generate
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_int_res_sign_ext
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:519:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:522:7
				always @(*) begin : assemble_result
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:524:9
					ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = {WIDTH {final_int[INT_WIDTH - 1]}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:525:9
					ifmt_pre_round_abs[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = final_int[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:528:7
				wire [WIDTH * 1:1] sv2v_tmp_F6FA8;
				assign sv2v_tmp_F6FA8 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = sv2v_tmp_F6FA8;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:533:3
	assign pre_round_abs = (dst_is_int_q ? ifmt_pre_round_abs[int_fmt_q2 * WIDTH+:WIDTH] : fmt_pre_round_abs[dst_fmt_q2 * WIDTH+:WIDTH]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:535:3
	fpnew_rounding #(.AbsWidth(WIDTH)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(input_sign_q),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(1'b0),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_true_zero)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:548:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:551:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_sign_inject
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:553:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:554:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:555:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:558:7
				always @(*) begin : post_process
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:560:9
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:561:9
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:564:9
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:565:9
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = (src_is_int_q & mant_is_zero_q ? {FP_WIDTH * 1 {1'sb0}} : {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]});
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:570:7
				wire [1:1] sv2v_tmp_4A747;
				assign sv2v_tmp_4A747 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4A747;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:571:7
				wire [1:1] sv2v_tmp_90681;
				assign sv2v_tmp_90681 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_90681;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:572:7
				wire [WIDTH * 1:1] sv2v_tmp_649FB;
				assign sv2v_tmp_649FB = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_649FB;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:577:3
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:578:3
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:581:3
	assign rounded_int_res = (rounded_sign ? $unsigned(-rounded_abs) : rounded_abs);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:582:3
	assign rounded_int_res_zero = rounded_int_res == {WIDTH {1'sb0}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:587:3
	wire [WIDTH - 1:0] fp_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:588:3
	wire [4:0] fp_special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:589:3
	wire fp_result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:591:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:594:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_special_results
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:596:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:597:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:598:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:600:5
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:601:5
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:604:7
				always @(*) begin : special_results
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:605:9
					reg [FP_WIDTH - 1:0] special_res;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:606:9
					special_res = (info_q[5] ? input_sign_q << (FP_WIDTH - 1) : {1'b0, QNAN_EXPONENT, QNAN_MANTISSA});
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:611:9
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:612:9
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:615:7
				wire [WIDTH * 1:1] sv2v_tmp_B718F;
				assign sv2v_tmp_B718F = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_B718F;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:620:3
	assign fp_result_is_special = ~src_is_int_q & ((info_q[5] | info_q[3]) | ~info_q[0]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:625:3
	assign fp_special_status = {info_q[2], 4'b0000};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:628:3
	assign fp_special_result = fmt_special_result[dst_fmt_q2 * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:633:3
	wire [WIDTH - 1:0] int_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:634:3
	wire [4:0] int_special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:635:3
	wire int_result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:637:3
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:640:3
	generate
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_special_results_int
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:642:5
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:645:7
				always @(*) begin : special_results
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:646:9
					reg [INT_WIDTH - 1:0] special_res;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:649:9
					special_res[INT_WIDTH - 2:0] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:650:9
					special_res[INT_WIDTH - 1] = op_mod_q2;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:653:9
					if (input_sign_q && !info_q[3])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:654:11
						special_res = ~special_res;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:657:9
					ifmt_special_result[ifmt * WIDTH+:WIDTH] = {WIDTH {special_res[INT_WIDTH - 1]}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:658:9
					ifmt_special_result[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:661:7
				wire [WIDTH * 1:1] sv2v_tmp_99B6D;
				assign sv2v_tmp_99B6D = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_special_result[ifmt * WIDTH+:WIDTH] = sv2v_tmp_99B6D;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:666:3
	assign int_result_is_special = (((info_q[3] | info_q[4]) | of_before_round) | ~info_q[0]) | ((input_sign_q & op_mod_q2) & ~rounded_int_res_zero);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:671:3
	assign int_special_status = 5'b10000;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:674:3
	assign int_special_result = ifmt_special_result[int_fmt_q2 * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:679:3
	wire [4:0] int_regular_status;
	wire [4:0] fp_regular_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:681:3
	wire [WIDTH - 1:0] fp_result;
	wire [WIDTH - 1:0] int_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:682:3
	wire [4:0] fp_status;
	wire [4:0] int_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:684:3
	assign fp_regular_status[4] = src_is_int_q & (of_before_round | of_after_round);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:685:3
	assign fp_regular_status[3] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:686:3
	assign fp_regular_status[2] = ~src_is_int_q & (~info_q[4] & (of_before_round | of_after_round));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:687:3
	assign fp_regular_status[1] = uf_after_round & fp_regular_status[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:688:3
	assign fp_regular_status[0] = (src_is_int_q ? |fp_round_sticky_bits : |fp_round_sticky_bits | (~info_q[4] & (of_before_round | of_after_round)));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:690:3
	assign int_regular_status = {4'b0000, |int_round_sticky_bits};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:692:3
	assign fp_result = (fp_result_is_special ? fp_special_result : fmt_result[dst_fmt_q2 * WIDTH+:WIDTH]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:693:3
	assign fp_status = (fp_result_is_special ? fp_special_status : fp_regular_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:694:3
	assign int_result = (int_result_is_special ? int_special_result : rounded_int_res);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:695:3
	assign int_status = (int_result_is_special ? int_special_status : int_regular_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:698:3
	wire [WIDTH - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:699:3
	wire [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:700:3
	wire extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:703:3
	assign result_d = (dst_is_int_q ? int_result : fp_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:704:3
	assign status_d = (dst_is_int_q ? int_status : fp_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:707:3
	assign extension_bit = (dst_is_int_q ? int_result[WIDTH - 1] : 1'b1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:713:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:714:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:715:3
	reg [0:NUM_OUT_REGS] out_pipe_ext_bit_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:716:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:717:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:718:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:720:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:723:3
	wire [WIDTH * 1:1] sv2v_tmp_4086F;
	assign sv2v_tmp_4086F = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_4086F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:724:3
	wire [5:1] sv2v_tmp_B7C45;
	assign sv2v_tmp_B7C45 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_B7C45;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:725:3
	wire [1:1] sv2v_tmp_8F736;
	assign sv2v_tmp_8F736 = extension_bit;
	always @(*) out_pipe_ext_bit_q[0] = sv2v_tmp_8F736;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:726:3
	wire [1:1] sv2v_tmp_DF7DA;
	assign sv2v_tmp_DF7DA = mid_pipe_tag_q[NUM_MID_REGS];
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_DF7DA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:727:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_F4B7F;
	assign sv2v_tmp_F4B7F = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_F4B7F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:728:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:730:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:732:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:734:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:738:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:740:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:740:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:740:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:740:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:742:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:744:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:744:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:744:181
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:744:289
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:745:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:745:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:745:181
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:745:289
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:746:69
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:746:125
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:746:181
					out_pipe_ext_bit_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:746:289
					out_pipe_ext_bit_q[i + 1] <= (reg_ena ? out_pipe_ext_bit_q[i] : out_pipe_ext_bit_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:747:79
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:747:135
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:747:191
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:747:299
					out_pipe_tag_q[i + 1] <= (reg_ena ? out_pipe_tag_q[i] : out_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:748:79
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:748:135
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:748:191
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:748:299
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:751:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:753:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:754:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:755:3
	assign extension_bit_o = out_pipe_ext_bit_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:756:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:757:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:758:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_cast_multi.sv:759:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_classifier (
	operands_i,
	is_boxed_i,
	info_o
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:15:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:16:13
	parameter [31:0] NumOperands = 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:18:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:20:3
	input wire [(NumOperands * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:21:3
	input wire [NumOperands - 1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:22:3
	// removed localparam type fpnew_pkg_fp_info_t
	output reg [(NumOperands * 8) - 1:0] info_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:25:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:26:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:29:3
	// removed localparam type fp_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:36:3
	genvar op;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (op = 0; op < sv2v_cast_32_signed(NumOperands); op = op + 1) begin : gen_num_values
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:38:5
			reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] value;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:39:5
			reg is_boxed;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:40:5
			reg is_normal;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:41:5
			reg is_inf;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:42:5
			reg is_nan;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:43:5
			reg is_signalling;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:44:5
			reg is_quiet;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:45:5
			reg is_zero;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:46:5
			reg is_subnormal;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:51:5
			always @(*) begin : classify_input
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:52:7
				value = operands_i[op * WIDTH+:WIDTH];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:53:7
				is_boxed = is_boxed_i[op];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:54:7
				is_normal = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] != {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] != {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}});
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:55:7
				is_zero = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && (value[MAN_BITS - 1-:MAN_BITS] == {MAN_BITS * 1 {1'sb0}});
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:56:7
				is_subnormal = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && !is_zero;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:57:7
				is_inf = is_boxed && ((value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}}) && (value[MAN_BITS - 1-:MAN_BITS] == {MAN_BITS * 1 {1'sb0}}));
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:58:7
				is_nan = !is_boxed || ((value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}}) && (value[MAN_BITS - 1-:MAN_BITS] != {MAN_BITS * 1 {1'sb0}}));
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:59:7
				is_signalling = (is_boxed && is_nan) && (value[(MAN_BITS - 1) - ((MAN_BITS - 1) - (MAN_BITS - 1))] == 1'b0);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:60:7
				is_quiet = is_nan && !is_signalling;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:62:7
				info_o[(op * 8) + 7] = is_normal;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:63:7
				info_o[(op * 8) + 6] = is_subnormal;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:64:7
				info_o[(op * 8) + 5] = is_zero;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:65:7
				info_o[(op * 8) + 4] = is_inf;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:66:7
				info_o[(op * 8) + 3] = is_nan;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:67:7
				info_o[(op * 8) + 2] = is_signalling;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:68:7
				info_o[(op * 8) + 1] = is_quiet;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_classifier.sv:69:7
				info_o[op * 8] = is_boxed;
			end
		end
	endgenerate
endmodule
module fpnew_divsqrt_multi_CBA5B_DFE5F (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	dst_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// removed localparam type TagType_TagType_TagType_TagType_TAGW_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:19:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:20:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:21:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:22:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:24:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:306:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:307:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:310:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:25:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:27:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:28:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:30:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:31:3
	input wire [9:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:32:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:33:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:34:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:35:3
	input wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:36:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:38:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:39:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:40:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:42:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:43:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:44:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:45:3
	output wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:46:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:48:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:49:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:51:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:58:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:63:3
	localparam NUM_OUT_REGS = ((PipeConfig == 2'd1) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:73:3
	wire [(2 * WIDTH) - 1:0] operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:74:3
	wire [2:0] rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:75:3
	wire [3:0] op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:76:3
	wire [2:0] dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:77:3
	wire in_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:80:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:81:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:82:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:83:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:84:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:85:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:86:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:88:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:91:3
	wire [2 * WIDTH:1] sv2v_tmp_83757;
	assign sv2v_tmp_83757 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_83757;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:92:3
	wire [3:1] sv2v_tmp_857E9;
	assign sv2v_tmp_857E9 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_857E9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:93:3
	wire [4:1] sv2v_tmp_4BFFB;
	assign sv2v_tmp_4BFFB = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_4BFFB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:94:3
	wire [3:1] sv2v_tmp_54055;
	assign sv2v_tmp_54055 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_54055;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:95:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_43752;
	assign sv2v_tmp_43752 = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_43752;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:96:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_3BDAF;
	assign sv2v_tmp_3BDAF = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_3BDAF;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:97:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:99:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:101:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] sv2v_cast_5B742;
		input reg [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] inp;
		sv2v_cast_5B742 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:103:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:107:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:109:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:109:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:109:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:109:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:111:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:113:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:113:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:113:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:113:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:114:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:114:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:114:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:114:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:115:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:115:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:115:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:115:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:116:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:116:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:116:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:116:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:117:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:117:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:117:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:117:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:118:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:118:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:118:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:118:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:121:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:122:3
	assign rnd_mode_q = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:123:3
	assign op_q = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:124:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:125:3
	assign in_valid_q = inp_pipe_valid_q[NUM_INP_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:130:3
	reg [1:0] divsqrt_fmt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:131:3
	reg [127:0] divsqrt_operands;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:132:3
	reg input_is_fp8;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:135:3
	always @(*) begin : translate_fmt
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:136:5
		case (dst_fmt_q)
			sv2v_cast_0BC43('d0):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:137:27
				divsqrt_fmt = 2'b00;
			sv2v_cast_0BC43('d1):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:138:27
				divsqrt_fmt = 2'b01;
			sv2v_cast_0BC43('d2):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:139:27
				divsqrt_fmt = 2'b10;
			sv2v_cast_0BC43('d4):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:140:27
				divsqrt_fmt = 2'b11;
			default:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:141:27
				divsqrt_fmt = 2'b10;
		endcase
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:145:5
		input_is_fp8 = FpFmtConfig[sv2v_cast_0BC43('d3)] & (dst_fmt_q == sv2v_cast_0BC43('d3));
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:148:5
		divsqrt_operands[0+:64] = (input_is_fp8 ? operands_q[0+:WIDTH] << 8 : operands_q[0+:WIDTH]);
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:149:5
		divsqrt_operands[64+:64] = (input_is_fp8 ? operands_q[WIDTH+:WIDTH] << 8 : operands_q[WIDTH+:WIDTH]);
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:155:3
	reg in_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:156:3
	wire div_valid;
	wire sqrt_valid;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:157:3
	wire unit_ready;
	wire unit_done;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:158:3
	wire op_starting;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:159:3
	reg out_valid;
	wire out_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:160:3
	reg hold_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:161:3
	reg data_is_held;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:162:3
	reg unit_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:164:3
	// removed localparam type fsm_state_e
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:165:3
	reg [1:0] state_q;
	reg [1:0] state_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:168:3
	assign inp_pipe_ready[NUM_INP_REGS] = in_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:171:3
	assign div_valid = ((in_valid_q & (op_q == sv2v_cast_A53F3(4))) & in_ready) & ~flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:172:3
	assign sqrt_valid = ((in_valid_q & (op_q != sv2v_cast_A53F3(4))) & in_ready) & ~flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:173:3
	assign op_starting = div_valid | sqrt_valid;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:176:3
	always @(*) begin : flag_fsm
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:178:5
		in_ready = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:179:5
		out_valid = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:180:5
		hold_result = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:181:5
		data_is_held = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:182:5
		unit_busy = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:183:5
		state_d = state_q;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:185:5
		case (state_q)
			2'd0: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:188:9
				in_ready = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:189:9
				if (in_valid_q && unit_ready)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:190:11
					state_d = 2'd1;
			end
			2'd1: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:195:9
				unit_busy = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:197:9
				if (unit_done) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:198:11
					out_valid = 1'b1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:200:11
					if (out_ready) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:201:13
						state_d = 2'd0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:202:13
						if (in_valid_q && unit_ready) begin
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:203:15
							in_ready = 1'b1;
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:204:15
							state_d = 2'd1;
						end
					end
					else begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:208:13
						hold_result = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:209:13
						state_d = 2'd2;
					end
				end
			end
			2'd2: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:215:9
				unit_busy = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:216:9
				data_is_held = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:217:9
				out_valid = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:219:9
				if (out_ready) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:220:11
					state_d = 2'd0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:221:11
					if (in_valid_q && unit_ready) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:222:13
						in_ready = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:223:13
						state_d = 2'd1;
					end
				end
			end
			default:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:228:16
				state_d = 2'd0;
		endcase
		if (flush_i) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:233:7
			unit_busy = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:234:7
			out_valid = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:235:7
			state_d = 2'd0;
		end
	end
	// Trace: macro expansion of FF at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:240:30
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:240:86
		if (!rst_ni)
			// Trace: macro expansion of FF at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:240:142
			state_q <= 2'd0;
		else
			// Trace: macro expansion of FF at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:240:250
			state_q <= state_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:243:3
	reg result_is_fp8_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:244:3
	reg [TagType_TagType_TagType_TagType_TAGW + 1:0] result_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:245:3
	reg [AuxType_AUX_BITS - 1:0] result_aux_q;
	// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:248:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:248:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:248:182
			result_is_fp8_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:248:290
			result_is_fp8_q <= (op_starting ? input_is_fp8 : result_is_fp8_q);
	// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:249:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:249:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:249:182
			result_tag_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:249:290
			result_tag_q <= (op_starting ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : result_tag_q);
	// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:250:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:250:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:250:182
			result_aux_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:250:290
			result_aux_q <= (op_starting ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : result_aux_q);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:255:3
	wire [63:0] unit_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:256:3
	wire [WIDTH - 1:0] adjusted_result;
	reg [WIDTH - 1:0] held_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:257:3
	wire [4:0] unit_status;
	reg [4:0] held_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:259:3
	// removed localparam type sv2v_uu_i_divsqrt_lei_Precision_ctl_SI
	localparam [5:0] sv2v_uu_i_divsqrt_lei_ext_Precision_ctl_SI_0 = 1'sb0;
	div_sqrt_top_mvp i_divsqrt_lei(
		.Clk_CI(clk_i),
		.Rst_RBI(rst_ni),
		.Div_start_SI(div_valid),
		.Sqrt_start_SI(sqrt_valid),
		.Operand_a_DI(divsqrt_operands[0+:64]),
		.Operand_b_DI(divsqrt_operands[64+:64]),
		.RM_SI(rnd_mode_q),
		.Precision_ctl_SI(sv2v_uu_i_divsqrt_lei_ext_Precision_ctl_SI_0),
		.Format_sel_SI(divsqrt_fmt),
		.Kill_SI(flush_i),
		.Result_DO(unit_result),
		.Fflags_SO(unit_status),
		.Ready_SO(unit_ready),
		.Done_SO(unit_done)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:277:3
	assign adjusted_result = (result_is_fp8_q ? unit_result >> 8 : unit_result);
	// Trace: macro expansion of FFLNR at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:280:58
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:280:100
		held_result_q <= (hold_result ? adjusted_result : held_result_q);
	// Trace: macro expansion of FFLNR at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:281:58
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:281:100
		held_status_q <= (hold_result ? unit_status : held_status_q);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:286:3
	wire [WIDTH - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:287:3
	wire [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:289:3
	assign result_d = (data_is_held ? held_result_q : adjusted_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:290:3
	assign status_d = (data_is_held ? held_status_q : unit_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:296:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:297:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:298:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:299:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:300:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:302:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:305:3
	wire [WIDTH * 1:1] sv2v_tmp_6C30D;
	assign sv2v_tmp_6C30D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6C30D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:306:3
	wire [5:1] sv2v_tmp_2ED07;
	assign sv2v_tmp_2ED07 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_2ED07;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:307:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_D5B68;
	assign sv2v_tmp_D5B68 = result_tag_q;
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_D5B68;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:308:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_62781;
	assign sv2v_tmp_62781 = result_aux_q;
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_62781;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:309:3
	wire [1:1] sv2v_tmp_D06FD;
	assign sv2v_tmp_D06FD = out_valid;
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_D06FD;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:311:3
	assign out_ready = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:313:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:315:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:319:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:321:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:321:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:321:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:321:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:323:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:325:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:325:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:325:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:325:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:326:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:326:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:326:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:326:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:327:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:327:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:327:189
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:327:297
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:328:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:328:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:328:189
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:328:297
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:331:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:333:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:334:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:335:3
	assign extension_bit_o = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:336:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:337:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:338:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:339:3
	assign busy_o = |{inp_pipe_valid_q, unit_busy, out_pipe_valid_q};
endmodule
module fpnew_divsqrt_multi_EA2AD_2C8BD (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	dst_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:19:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:20:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:21:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:22:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:24:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:306:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:307:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:310:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:25:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:27:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:28:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:30:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:31:3
	input wire [9:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:32:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:33:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:34:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:35:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:36:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:38:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:39:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:40:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:42:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:43:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:44:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:45:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:46:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:48:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:49:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:51:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:58:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:63:3
	localparam NUM_OUT_REGS = ((PipeConfig == 2'd1) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:73:3
	wire [(2 * WIDTH) - 1:0] operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:74:3
	wire [2:0] rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:75:3
	wire [3:0] op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:76:3
	wire [2:0] dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:77:3
	wire in_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:80:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:81:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:82:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:83:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:84:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:85:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:86:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:88:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:91:3
	wire [2 * WIDTH:1] sv2v_tmp_83757;
	assign sv2v_tmp_83757 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_83757;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:92:3
	wire [3:1] sv2v_tmp_857E9;
	assign sv2v_tmp_857E9 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_857E9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:93:3
	wire [4:1] sv2v_tmp_4BFFB;
	assign sv2v_tmp_4BFFB = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_4BFFB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:94:3
	wire [3:1] sv2v_tmp_54055;
	assign sv2v_tmp_54055 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_54055;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:95:3
	wire [1:1] sv2v_tmp_76699;
	assign sv2v_tmp_76699 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_76699;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:96:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_D1879;
	assign sv2v_tmp_D1879 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_D1879;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:97:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:99:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:101:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:103:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:107:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:109:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:109:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:109:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:109:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:111:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:113:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:113:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:113:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:113:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:114:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:114:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:114:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:114:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:115:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:115:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:115:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:115:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:116:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:116:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:116:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:116:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:117:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:117:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:117:193
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:117:301
					inp_pipe_tag_q[i + 1] <= (reg_ena ? inp_pipe_tag_q[i] : inp_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:118:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:118:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:118:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:118:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:121:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:122:3
	assign rnd_mode_q = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:123:3
	assign op_q = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:124:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:125:3
	assign in_valid_q = inp_pipe_valid_q[NUM_INP_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:130:3
	reg [1:0] divsqrt_fmt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:131:3
	reg [127:0] divsqrt_operands;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:132:3
	reg input_is_fp8;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:135:3
	always @(*) begin : translate_fmt
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:136:5
		case (dst_fmt_q)
			sv2v_cast_0BC43('d0):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:137:27
				divsqrt_fmt = 2'b00;
			sv2v_cast_0BC43('d1):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:138:27
				divsqrt_fmt = 2'b01;
			sv2v_cast_0BC43('d2):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:139:27
				divsqrt_fmt = 2'b10;
			sv2v_cast_0BC43('d4):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:140:27
				divsqrt_fmt = 2'b11;
			default:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:141:27
				divsqrt_fmt = 2'b10;
		endcase
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:145:5
		input_is_fp8 = FpFmtConfig[sv2v_cast_0BC43('d3)] & (dst_fmt_q == sv2v_cast_0BC43('d3));
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:148:5
		divsqrt_operands[0+:64] = (input_is_fp8 ? operands_q[0+:WIDTH] << 8 : operands_q[0+:WIDTH]);
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:149:5
		divsqrt_operands[64+:64] = (input_is_fp8 ? operands_q[WIDTH+:WIDTH] << 8 : operands_q[WIDTH+:WIDTH]);
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:155:3
	reg in_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:156:3
	wire div_valid;
	wire sqrt_valid;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:157:3
	wire unit_ready;
	wire unit_done;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:158:3
	wire op_starting;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:159:3
	reg out_valid;
	wire out_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:160:3
	reg hold_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:161:3
	reg data_is_held;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:162:3
	reg unit_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:164:3
	// removed localparam type fsm_state_e
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:165:3
	reg [1:0] state_q;
	reg [1:0] state_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:168:3
	assign inp_pipe_ready[NUM_INP_REGS] = in_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:171:3
	assign div_valid = ((in_valid_q & (op_q == sv2v_cast_A53F3(4))) & in_ready) & ~flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:172:3
	assign sqrt_valid = ((in_valid_q & (op_q != sv2v_cast_A53F3(4))) & in_ready) & ~flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:173:3
	assign op_starting = div_valid | sqrt_valid;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:176:3
	always @(*) begin : flag_fsm
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:178:5
		in_ready = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:179:5
		out_valid = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:180:5
		hold_result = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:181:5
		data_is_held = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:182:5
		unit_busy = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:183:5
		state_d = state_q;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:185:5
		case (state_q)
			2'd0: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:188:9
				in_ready = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:189:9
				if (in_valid_q && unit_ready)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:190:11
					state_d = 2'd1;
			end
			2'd1: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:195:9
				unit_busy = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:197:9
				if (unit_done) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:198:11
					out_valid = 1'b1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:200:11
					if (out_ready) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:201:13
						state_d = 2'd0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:202:13
						if (in_valid_q && unit_ready) begin
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:203:15
							in_ready = 1'b1;
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:204:15
							state_d = 2'd1;
						end
					end
					else begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:208:13
						hold_result = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:209:13
						state_d = 2'd2;
					end
				end
			end
			2'd2: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:215:9
				unit_busy = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:216:9
				data_is_held = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:217:9
				out_valid = 1'b1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:219:9
				if (out_ready) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:220:11
					state_d = 2'd0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:221:11
					if (in_valid_q && unit_ready) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:222:13
						in_ready = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:223:13
						state_d = 2'd1;
					end
				end
			end
			default:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:228:16
				state_d = 2'd0;
		endcase
		if (flush_i) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:233:7
			unit_busy = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:234:7
			out_valid = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:235:7
			state_d = 2'd0;
		end
	end
	// Trace: macro expansion of FF at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:240:30
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FF at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:240:86
		if (!rst_ni)
			// Trace: macro expansion of FF at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:240:142
			state_q <= 2'd0;
		else
			// Trace: macro expansion of FF at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:240:250
			state_q <= state_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:243:3
	reg result_is_fp8_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:244:3
	reg result_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:245:3
	reg [AuxType_AUX_BITS - 1:0] result_aux_q;
	// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:248:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:248:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:248:182
			result_is_fp8_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:248:290
			result_is_fp8_q <= (op_starting ? input_is_fp8 : result_is_fp8_q);
	// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:249:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:249:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:249:182
			result_tag_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:249:290
			result_tag_q <= (op_starting ? inp_pipe_tag_q[NUM_INP_REGS] : result_tag_q);
	// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:250:70
	always @(posedge clk_i or negedge rst_ni)
		// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:250:126
		if (!rst_ni)
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:250:182
			result_aux_q <= 1'sb0;
		else
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:250:290
			result_aux_q <= (op_starting ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : result_aux_q);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:255:3
	wire [63:0] unit_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:256:3
	wire [WIDTH - 1:0] adjusted_result;
	reg [WIDTH - 1:0] held_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:257:3
	wire [4:0] unit_status;
	reg [4:0] held_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:259:3
	// removed localparam type sv2v_uu_i_divsqrt_lei_Precision_ctl_SI
	localparam [5:0] sv2v_uu_i_divsqrt_lei_ext_Precision_ctl_SI_0 = 1'sb0;
	div_sqrt_top_mvp i_divsqrt_lei(
		.Clk_CI(clk_i),
		.Rst_RBI(rst_ni),
		.Div_start_SI(div_valid),
		.Sqrt_start_SI(sqrt_valid),
		.Operand_a_DI(divsqrt_operands[0+:64]),
		.Operand_b_DI(divsqrt_operands[64+:64]),
		.RM_SI(rnd_mode_q),
		.Precision_ctl_SI(sv2v_uu_i_divsqrt_lei_ext_Precision_ctl_SI_0),
		.Format_sel_SI(divsqrt_fmt),
		.Kill_SI(flush_i),
		.Result_DO(unit_result),
		.Fflags_SO(unit_status),
		.Ready_SO(unit_ready),
		.Done_SO(unit_done)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:277:3
	assign adjusted_result = (result_is_fp8_q ? unit_result >> 8 : unit_result);
	// Trace: macro expansion of FFLNR at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:280:58
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:280:100
		held_result_q <= (hold_result ? adjusted_result : held_result_q);
	// Trace: macro expansion of FFLNR at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:281:58
	always @(posedge clk_i)
		// Trace: macro expansion of FFLNR at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:281:100
		held_status_q <= (hold_result ? unit_status : held_status_q);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:286:3
	wire [WIDTH - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:287:3
	wire [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:289:3
	assign result_d = (data_is_held ? held_result_q : adjusted_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:290:3
	assign status_d = (data_is_held ? held_status_q : unit_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:296:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:297:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:298:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:299:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:300:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:302:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:305:3
	wire [WIDTH * 1:1] sv2v_tmp_6C30D;
	assign sv2v_tmp_6C30D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6C30D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:306:3
	wire [5:1] sv2v_tmp_2ED07;
	assign sv2v_tmp_2ED07 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_2ED07;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:307:3
	wire [1:1] sv2v_tmp_0F1D1;
	assign sv2v_tmp_0F1D1 = result_tag_q;
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_0F1D1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:308:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_46FBB;
	assign sv2v_tmp_46FBB = result_aux_q;
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_46FBB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:309:3
	wire [1:1] sv2v_tmp_D06FD;
	assign sv2v_tmp_D06FD = out_valid;
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_D06FD;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:311:3
	assign out_ready = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:313:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:315:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:319:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:321:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:321:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:321:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:321:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:323:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:325:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:325:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:325:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:325:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:326:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:326:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:326:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:326:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:327:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:327:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:327:189
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:327:297
					out_pipe_tag_q[i + 1] <= (reg_ena ? out_pipe_tag_q[i] : out_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:328:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:328:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:328:189
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:328:297
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:331:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:333:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:334:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:335:3
	assign extension_bit_o = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:336:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:337:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:338:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_divsqrt_multi.sv:339:3
	assign busy_o = |{inp_pipe_valid_q, unit_busy, out_pipe_valid_q};
endmodule
module fpnew_fma_141C6 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:18:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:19:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:20:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:21:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:23:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:25:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:26:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:28:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:29:3
	input wire [2:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:30:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:31:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:32:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:33:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:34:3
	input wire aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:36:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:37:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:38:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:40:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:41:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:42:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:43:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:44:3
	output wire aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:46:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:47:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:49:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:55:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:56:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:57:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:334:40
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:335:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	localparam [31:0] BIAS = fpnew_pkg_bias(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:59:3
	localparam [31:0] PRECISION_BITS = MAN_BITS + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:61:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:62:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:66:3
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	localparam [31:0] EXP_WIDTH = $unsigned(fpnew_pkg_maximum(EXP_BITS + 2, LZC_RESULT_WIDTH));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:68:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 3);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:70:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:75:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:80:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:89:3
	// removed localparam type fp_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:99:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:100:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:101:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:102:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:103:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:104:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:105:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:106:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:108:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:111:3
	wire [3 * WIDTH:1] sv2v_tmp_BC8B9;
	assign sv2v_tmp_BC8B9 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_BC8B9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:112:3
	wire [3:1] sv2v_tmp_FE389;
	assign sv2v_tmp_FE389 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_FE389;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:113:3
	wire [3:1] sv2v_tmp_E1339;
	assign sv2v_tmp_E1339 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_E1339;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:114:3
	wire [4:1] sv2v_tmp_CBA8F;
	assign sv2v_tmp_CBA8F = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_CBA8F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:115:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:116:3
	wire [1:1] sv2v_tmp_76699;
	assign sv2v_tmp_76699 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_76699;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:117:3
	wire [1:1] sv2v_tmp_8D189;
	assign sv2v_tmp_8D189 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_8D189;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:118:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:120:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:122:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:124:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:128:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:130:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:130:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:130:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:130:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:132:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:134:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:134:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:134:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:134:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:135:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:135:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:135:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:135:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:136:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:136:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:136:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:136:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:137:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:137:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:137:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:137:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:138:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:138:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:138:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:138:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:139:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:139:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:139:193
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:139:301
					inp_pipe_tag_q[i + 1] <= (reg_ena ? inp_pipe_tag_q[i] : inp_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:140:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:140:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:140:193
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:140:301
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:146:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [23:0] info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:149:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(3)
	) i_class_inputs(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3]),
		.info_o(info_q)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:158:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:159:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:173:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_91364;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_91364 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_60B87;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_60B87 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_F33EE;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_F33EE = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_14681;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_14681 = inp;
	endfunction
	always @(*) begin : op_select
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:176:5
		operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:177:5
		operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:178:5
		operand_c = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:179:5
		info_a = info_q[0+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:180:5
		info_b = info_q[8+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:181:5
		info_c = info_q[16+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:184:5
		operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] = operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:186:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(0):
				;
			sv2v_cast_A53F3(1):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:188:26
				operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] = ~operand_a[1 + (EXP_BITS + (MAN_BITS - 1))];
			sv2v_cast_A53F3(2): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:190:9
				operand_a = {1'b0, sv2v_cast_91364(BIAS), sv2v_cast_60B87(1'sb0)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:191:9
				info_a = 8'b10000001;
			end
			sv2v_cast_A53F3(3): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:194:9
				operand_c = {1'b1, sv2v_cast_F33EE(1'sb0), sv2v_cast_60B87(1'sb0)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:195:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:198:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:199:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:200:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:201:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:202:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:203:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:211:3
	wire any_operand_inf;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:212:3
	wire any_operand_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:213:3
	wire signalling_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:214:3
	wire effective_subtraction;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:215:3
	wire tentative_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:218:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:219:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:220:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:222:3
	assign effective_subtraction = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]) ^ operand_c[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:224:3
	assign tentative_sign = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:229:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:230:3
	reg [4:0] special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:231:3
	reg result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:233:3
	always @(*) begin : special_cases
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:235:5
		special_result = {1'b0, sv2v_cast_F33EE(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:236:5
		special_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:237:5
		result_is_special = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:243:5
		if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:244:7
			result_is_special = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:245:7
			special_status[4] = 1'b1;
		end
		else if (any_operand_nan) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:248:7
			result_is_special = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:249:7
			special_status[4] = signalling_nan;
		end
		else if (any_operand_inf) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:252:7
			result_is_special = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:254:7
			if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:255:9
				special_status[4] = 1'b1;
			else if (info_a[4] || info_b[4])
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:259:9
				special_result = {operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_F33EE(1'sb1), sv2v_cast_60B87(1'sb0)};
			else if (info_c[4])
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:263:9
				special_result = {operand_c[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_F33EE(1'sb1), sv2v_cast_60B87(1'sb0)};
		end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:271:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:272:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:273:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:276:3
	assign exponent_a = $signed({1'b0, operand_a[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:277:3
	assign exponent_b = $signed({1'b0, operand_b[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:278:3
	assign exponent_c = $signed({1'b0, operand_c[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:282:3
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:284:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(BIAS) : $signed((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - $signed(BIAS)));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:290:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:292:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:295:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:297:3
	always @(*) begin : addend_shift_amount
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:299:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:300:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:303:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:306:7
			addend_shamt = 0;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:312:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:313:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:314:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:317:3
	assign mantissa_a = {info_a[7], operand_a[MAN_BITS - 1-:MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:318:3
	assign mantissa_b = {info_b[7], operand_b[MAN_BITS - 1-:MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:319:3
	assign mantissa_c = {info_c[7], operand_c[MAN_BITS - 1-:MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:322:3
	assign product = mantissa_a * mantissa_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:327:3
	assign product_shifted = product << 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:332:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:333:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:334:3
	wire sticky_before_add;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:335:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:336:3
	wire inject_carry_in;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:346:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:349:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:353:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:354:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:359:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:360:3
	wire sum_carry;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:361:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:362:3
	wire final_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:365:3
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:366:3
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:369:3
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:372:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:380:3
	wire effective_subtraction_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:381:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:382:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:383:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:384:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:385:3
	wire sticky_before_add_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:386:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:387:3
	wire final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:388:3
	wire [2:0] rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:389:3
	wire result_is_special_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:390:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:391:3
	wire [4:0] special_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:393:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:394:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:395:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:396:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:397:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:398:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:399:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:400:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:401:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:402:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:403:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:404:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:405:3
	reg [0:NUM_MID_REGS] mid_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:406:3
	reg [0:NUM_MID_REGS] mid_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:407:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:409:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:412:3
	wire [1:1] sv2v_tmp_56A72;
	assign sv2v_tmp_56A72 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_56A72;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:413:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_2D21E;
	assign sv2v_tmp_2D21E = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_2D21E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:414:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_00793;
	assign sv2v_tmp_00793 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_00793;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:415:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_B4C85;
	assign sv2v_tmp_B4C85 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_B4C85;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:416:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_83404;
	assign sv2v_tmp_83404 = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_83404;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:417:3
	wire [1:1] sv2v_tmp_6F5F7;
	assign sv2v_tmp_6F5F7 = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6F5F7;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:418:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_CEAB3;
	assign sv2v_tmp_CEAB3 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_CEAB3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:419:3
	wire [1:1] sv2v_tmp_D7BD0;
	assign sv2v_tmp_D7BD0 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_D7BD0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:420:3
	wire [3:1] sv2v_tmp_A74E2;
	assign sv2v_tmp_A74E2 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_A74E2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:421:3
	wire [1:1] sv2v_tmp_7DEC5;
	assign sv2v_tmp_7DEC5 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_7DEC5;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:422:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_4A83E;
	assign sv2v_tmp_4A83E = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_4A83E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:423:3
	wire [5:1] sv2v_tmp_EC01B;
	assign sv2v_tmp_EC01B = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_EC01B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:424:3
	wire [1:1] sv2v_tmp_44BCE;
	assign sv2v_tmp_44BCE = inp_pipe_tag_q[NUM_INP_REGS];
	always @(*) mid_pipe_tag_q[0] = sv2v_tmp_44BCE;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:425:3
	wire [1:1] sv2v_tmp_CDA0E;
	assign sv2v_tmp_CDA0E = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) mid_pipe_aux_q[0] = sv2v_tmp_CDA0E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:426:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:428:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:431:3
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:433:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:437:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:439:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:439:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:439:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:439:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:441:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:443:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:443:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:443:189
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:443:297
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:444:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:444:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:444:189
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:444:297
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:445:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:445:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:445:189
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:445:297
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:446:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:446:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:446:189
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:446:297
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:447:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:447:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:447:189
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:447:297
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:448:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:448:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:448:189
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:448:297
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:449:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:449:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:449:189
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:449:297
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:450:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:450:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:450:189
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:450:297
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:451:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:451:145
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:451:201
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:451:309
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:452:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:452:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:452:189
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:452:297
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:453:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:453:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:453:189
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:453:297
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:454:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:454:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:454:189
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:454:297
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:455:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:455:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:455:199
					mid_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:455:307
					mid_pipe_tag_q[i + 1] <= (reg_ena ? mid_pipe_tag_q[i] : mid_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:456:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:456:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:456:199
					mid_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:456:307
					mid_pipe_aux_q[i + 1] <= (reg_ena ? mid_pipe_aux_q[i] : mid_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:459:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:460:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:461:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:462:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:463:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:464:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:465:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:466:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:467:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:468:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:469:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:470:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:475:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:476:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:477:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:478:3
	wire lzc_zeroes;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:480:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:481:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:483:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:484:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:485:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:486:3
	wire sticky_after_norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:488:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:490:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:493:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:502:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:505:3
	always @(*) begin : norm_shift_amount
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:507:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:509:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:511:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:512:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:516:9
					norm_shamt = $unsigned(($signed(PRECISION_BITS) + 2) + exponent_product_q);
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:517:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:521:7
			norm_shamt = addend_shamt_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:522:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:527:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:531:3
	always @(*) begin : small_norm
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:533:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:534:5
		final_exponent = normalized_exponent;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:537:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:538:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:539:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:545:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:546:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:549:7
			final_exponent = 1'sb0;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:554:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:559:3
	wire pre_round_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:560:3
	wire [EXP_BITS - 1:0] pre_round_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:561:3
	wire [MAN_BITS - 1:0] pre_round_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:562:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:563:3
	wire [1:0] round_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:565:3
	wire of_before_round;
	wire of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:566:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:567:3
	wire result_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:569:3
	wire rounded_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:570:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] rounded_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:573:3
	assign of_before_round = final_exponent >= ((2 ** EXP_BITS) - 1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:574:3
	assign uf_before_round = final_exponent == 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:577:3
	assign pre_round_sign = final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:578:3
	assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : $unsigned(final_exponent[EXP_BITS - 1:0]));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:579:3
	assign pre_round_mantissa = (of_before_round ? {MAN_BITS {1'sb1}} : final_mantissa[MAN_BITS:1]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:580:3
	assign pre_round_abs = {pre_round_exponent, pre_round_mantissa};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:583:3
	assign round_sticky_bits = (of_before_round ? 2'b11 : {final_mantissa[0], sticky_after_norm});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:586:3
	fpnew_rounding #(.AbsWidth(EXP_BITS + MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:600:3
	assign uf_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:601:3
	assign of_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:606:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:607:3
	wire [4:0] regular_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:610:3
	assign regular_result = {rounded_sign, rounded_abs};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:611:3
	assign regular_status[4] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:612:3
	assign regular_status[3] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:613:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:614:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:615:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:618:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:619:3
	wire [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:622:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:623:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:629:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:630:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:631:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:632:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:633:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:635:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:638:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_0252C;
	assign sv2v_tmp_0252C = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_0252C;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:639:3
	wire [5:1] sv2v_tmp_2A843;
	assign sv2v_tmp_2A843 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_2A843;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:640:3
	wire [1:1] sv2v_tmp_DF7DA;
	assign sv2v_tmp_DF7DA = mid_pipe_tag_q[NUM_MID_REGS];
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_DF7DA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:641:3
	wire [1:1] sv2v_tmp_9E262;
	assign sv2v_tmp_9E262 = mid_pipe_aux_q[NUM_MID_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_9E262;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:642:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:644:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:646:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:648:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:652:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:654:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:654:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:654:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:654:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:656:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:658:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:658:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:658:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:658:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:659:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:659:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:659:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:659:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:660:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:660:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:660:189
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:660:297
					out_pipe_tag_q[i + 1] <= (reg_ena ? out_pipe_tag_q[i] : out_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:661:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:661:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:661:189
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:661:297
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:664:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:666:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:667:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:668:3
	assign extension_bit_o = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:669:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:670:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:671:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:672:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_fma_1D182_0A4E9 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TagType_TagType_TagType_TAGW_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:18:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:19:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:20:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:21:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:23:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:25:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:26:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:28:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:29:3
	input wire [2:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:30:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:31:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:32:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:33:3
	input wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:34:3
	input wire aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:36:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:37:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:38:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:40:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:41:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:42:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:43:3
	output wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:44:3
	output wire aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:46:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:47:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:49:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:55:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:56:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:57:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:334:40
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:335:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	localparam [31:0] BIAS = fpnew_pkg_bias(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:59:3
	localparam [31:0] PRECISION_BITS = MAN_BITS + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:61:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:62:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:66:3
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	localparam [31:0] EXP_WIDTH = $unsigned(fpnew_pkg_maximum(EXP_BITS + 2, LZC_RESULT_WIDTH));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:68:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 3);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:70:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:75:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:80:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:89:3
	// removed localparam type fp_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:99:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:100:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:101:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:102:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:103:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:104:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:105:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:106:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:108:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:111:3
	wire [3 * WIDTH:1] sv2v_tmp_BC8B9;
	assign sv2v_tmp_BC8B9 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_BC8B9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:112:3
	wire [3:1] sv2v_tmp_FE389;
	assign sv2v_tmp_FE389 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_FE389;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:113:3
	wire [3:1] sv2v_tmp_E1339;
	assign sv2v_tmp_E1339 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_E1339;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:114:3
	wire [4:1] sv2v_tmp_CBA8F;
	assign sv2v_tmp_CBA8F = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_CBA8F;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:115:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:116:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_35336;
	assign sv2v_tmp_35336 = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_35336;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:117:3
	wire [1:1] sv2v_tmp_8D189;
	assign sv2v_tmp_8D189 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_8D189;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:118:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:120:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:122:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] sv2v_cast_5B742;
		input reg [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] inp;
		sv2v_cast_5B742 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:124:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:128:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:130:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:130:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:130:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:130:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:132:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:134:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:134:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:134:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:134:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:135:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:135:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:135:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:135:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:136:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:136:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:136:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:136:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:137:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:137:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:137:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:137:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:138:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:138:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:138:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:138:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:139:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:139:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:139:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:139:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:140:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:140:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:140:193
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:140:301
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:146:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [23:0] info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:149:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(3)
	) i_class_inputs(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3]),
		.info_o(info_q)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:158:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:159:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:173:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_91364;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_91364 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_60B87;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_60B87 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_F33EE;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_F33EE = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_14681;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_14681 = inp;
	endfunction
	always @(*) begin : op_select
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:176:5
		operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:177:5
		operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:178:5
		operand_c = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:179:5
		info_a = info_q[0+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:180:5
		info_b = info_q[8+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:181:5
		info_c = info_q[16+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:184:5
		operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] = operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:186:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(0):
				;
			sv2v_cast_A53F3(1):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:188:26
				operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] = ~operand_a[1 + (EXP_BITS + (MAN_BITS - 1))];
			sv2v_cast_A53F3(2): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:190:9
				operand_a = {1'b0, sv2v_cast_91364(BIAS), sv2v_cast_60B87(1'sb0)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:191:9
				info_a = 8'b10000001;
			end
			sv2v_cast_A53F3(3): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:194:9
				operand_c = {1'b1, sv2v_cast_F33EE(1'sb0), sv2v_cast_60B87(1'sb0)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:195:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:198:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:199:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:200:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:201:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:202:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:203:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:211:3
	wire any_operand_inf;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:212:3
	wire any_operand_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:213:3
	wire signalling_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:214:3
	wire effective_subtraction;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:215:3
	wire tentative_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:218:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:219:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:220:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:222:3
	assign effective_subtraction = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]) ^ operand_c[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:224:3
	assign tentative_sign = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:229:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:230:3
	reg [4:0] special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:231:3
	reg result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:233:3
	always @(*) begin : special_cases
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:235:5
		special_result = {1'b0, sv2v_cast_F33EE(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:236:5
		special_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:237:5
		result_is_special = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:243:5
		if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:244:7
			result_is_special = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:245:7
			special_status[4] = 1'b1;
		end
		else if (any_operand_nan) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:248:7
			result_is_special = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:249:7
			special_status[4] = signalling_nan;
		end
		else if (any_operand_inf) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:252:7
			result_is_special = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:254:7
			if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:255:9
				special_status[4] = 1'b1;
			else if (info_a[4] || info_b[4])
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:259:9
				special_result = {operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_F33EE(1'sb1), sv2v_cast_60B87(1'sb0)};
			else if (info_c[4])
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:263:9
				special_result = {operand_c[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_F33EE(1'sb1), sv2v_cast_60B87(1'sb0)};
		end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:271:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:272:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:273:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:276:3
	assign exponent_a = $signed({1'b0, operand_a[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:277:3
	assign exponent_b = $signed({1'b0, operand_b[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:278:3
	assign exponent_c = $signed({1'b0, operand_c[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:282:3
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:284:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(BIAS) : $signed((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - $signed(BIAS)));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:290:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:292:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:295:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:297:3
	always @(*) begin : addend_shift_amount
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:299:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:300:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:303:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:306:7
			addend_shamt = 0;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:312:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:313:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:314:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:317:3
	assign mantissa_a = {info_a[7], operand_a[MAN_BITS - 1-:MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:318:3
	assign mantissa_b = {info_b[7], operand_b[MAN_BITS - 1-:MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:319:3
	assign mantissa_c = {info_c[7], operand_c[MAN_BITS - 1-:MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:322:3
	assign product = mantissa_a * mantissa_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:327:3
	assign product_shifted = product << 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:332:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:333:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:334:3
	wire sticky_before_add;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:335:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:336:3
	wire inject_carry_in;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:346:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:349:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:353:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:354:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:359:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:360:3
	wire sum_carry;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:361:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:362:3
	wire final_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:365:3
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:366:3
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:369:3
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:372:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:380:3
	wire effective_subtraction_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:381:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:382:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:383:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:384:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:385:3
	wire sticky_before_add_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:386:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:387:3
	wire final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:388:3
	wire [2:0] rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:389:3
	wire result_is_special_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:390:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:391:3
	wire [4:0] special_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:393:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:394:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:395:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:396:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:397:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:398:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:399:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:400:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:401:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:402:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:403:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:404:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:405:3
	reg [(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_MID_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_MID_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_MID_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_MID_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] mid_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:406:3
	reg [0:NUM_MID_REGS] mid_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:407:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:409:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:412:3
	wire [1:1] sv2v_tmp_56A72;
	assign sv2v_tmp_56A72 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_56A72;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:413:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_2D21E;
	assign sv2v_tmp_2D21E = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_2D21E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:414:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_00793;
	assign sv2v_tmp_00793 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_00793;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:415:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_B4C85;
	assign sv2v_tmp_B4C85 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_B4C85;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:416:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_83404;
	assign sv2v_tmp_83404 = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_83404;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:417:3
	wire [1:1] sv2v_tmp_6F5F7;
	assign sv2v_tmp_6F5F7 = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6F5F7;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:418:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_CEAB3;
	assign sv2v_tmp_CEAB3 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_CEAB3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:419:3
	wire [1:1] sv2v_tmp_D7BD0;
	assign sv2v_tmp_D7BD0 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_D7BD0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:420:3
	wire [3:1] sv2v_tmp_A74E2;
	assign sv2v_tmp_A74E2 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_A74E2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:421:3
	wire [1:1] sv2v_tmp_7DEC5;
	assign sv2v_tmp_7DEC5 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_7DEC5;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:422:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_4A83E;
	assign sv2v_tmp_4A83E = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_4A83E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:423:3
	wire [5:1] sv2v_tmp_EC01B;
	assign sv2v_tmp_EC01B = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_EC01B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:424:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_D3C2C;
	assign sv2v_tmp_D3C2C = inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	always @(*) mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_D3C2C;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:425:3
	wire [1:1] sv2v_tmp_CDA0E;
	assign sv2v_tmp_CDA0E = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) mid_pipe_aux_q[0] = sv2v_tmp_CDA0E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:426:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:428:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:431:3
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:433:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:437:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:439:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:439:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:439:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:439:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:441:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:443:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:443:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:443:189
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:443:297
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:444:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:444:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:444:189
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:444:297
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:445:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:445:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:445:189
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:445:297
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:446:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:446:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:446:189
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:446:297
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:447:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:447:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:447:189
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:447:297
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:448:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:448:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:448:189
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:448:297
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:449:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:449:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:449:189
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:449:297
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:450:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:450:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:450:189
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:450:297
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:451:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:451:145
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:451:201
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:451:309
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:452:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:452:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:452:189
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:452:297
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:453:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:453:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:453:189
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:453:297
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:454:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:454:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:454:189
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:454:297
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:455:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:455:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:455:199
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:455:307
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:456:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:456:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:456:199
					mid_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:456:307
					mid_pipe_aux_q[i + 1] <= (reg_ena ? mid_pipe_aux_q[i] : mid_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:459:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:460:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:461:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:462:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:463:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:464:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:465:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:466:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:467:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:468:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:469:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:470:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:475:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:476:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:477:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:478:3
	wire lzc_zeroes;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:480:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:481:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:483:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:484:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:485:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:486:3
	wire sticky_after_norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:488:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:490:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:493:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:502:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:505:3
	always @(*) begin : norm_shift_amount
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:507:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:509:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:511:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:512:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:516:9
					norm_shamt = $unsigned(($signed(PRECISION_BITS) + 2) + exponent_product_q);
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:517:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:521:7
			norm_shamt = addend_shamt_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:522:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:527:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:531:3
	always @(*) begin : small_norm
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:533:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:534:5
		final_exponent = normalized_exponent;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:537:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:538:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:539:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:545:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:546:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:549:7
			final_exponent = 1'sb0;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:554:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:559:3
	wire pre_round_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:560:3
	wire [EXP_BITS - 1:0] pre_round_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:561:3
	wire [MAN_BITS - 1:0] pre_round_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:562:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:563:3
	wire [1:0] round_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:565:3
	wire of_before_round;
	wire of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:566:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:567:3
	wire result_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:569:3
	wire rounded_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:570:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] rounded_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:573:3
	assign of_before_round = final_exponent >= ((2 ** EXP_BITS) - 1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:574:3
	assign uf_before_round = final_exponent == 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:577:3
	assign pre_round_sign = final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:578:3
	assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : $unsigned(final_exponent[EXP_BITS - 1:0]));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:579:3
	assign pre_round_mantissa = (of_before_round ? {MAN_BITS {1'sb1}} : final_mantissa[MAN_BITS:1]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:580:3
	assign pre_round_abs = {pre_round_exponent, pre_round_mantissa};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:583:3
	assign round_sticky_bits = (of_before_round ? 2'b11 : {final_mantissa[0], sticky_after_norm});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:586:3
	fpnew_rounding #(.AbsWidth(EXP_BITS + MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:600:3
	assign uf_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:601:3
	assign of_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:606:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:607:3
	wire [4:0] regular_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:610:3
	assign regular_result = {rounded_sign, rounded_abs};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:611:3
	assign regular_status[4] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:612:3
	assign regular_status[3] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:613:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:614:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:615:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:618:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:619:3
	wire [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:622:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:623:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:629:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:630:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:631:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:632:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:633:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:635:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:638:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_0252C;
	assign sv2v_tmp_0252C = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_0252C;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:639:3
	wire [5:1] sv2v_tmp_2A843;
	assign sv2v_tmp_2A843 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_2A843;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:640:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_0C03D;
	assign sv2v_tmp_0C03D = mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_0C03D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:641:3
	wire [1:1] sv2v_tmp_9E262;
	assign sv2v_tmp_9E262 = mid_pipe_aux_q[NUM_MID_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_9E262;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:642:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:644:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:646:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:648:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:652:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:654:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:654:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:654:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:654:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:656:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:658:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:658:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:658:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:658:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:659:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:659:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:659:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:659:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:660:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:660:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:660:189
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:660:297
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:661:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:661:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:661:189
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:661:297
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:664:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:666:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:667:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:668:3
	assign extension_bit_o = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:669:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:670:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:671:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma.sv:672:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_fma_multi_53FD4_8108B (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// removed localparam type TagType_TagType_TagType_TagType_TAGW_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:18:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:19:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:20:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:21:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:23:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:306:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:307:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:310:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:24:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:26:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:27:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:29:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:30:3
	input wire [14:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:31:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:32:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:33:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:34:3
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:35:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:36:3
	input wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:37:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:39:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:40:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:41:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:43:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:44:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:45:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:46:3
	output wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:47:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:49:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:50:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:52:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:59:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:338:49
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:339:5
		reg [63:0] res;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:340:5
			res = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:5
			begin : sv2v_autoblock_2
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:10
				reg [31:0] fmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:343:9
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt))));
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:344:9
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:61:3
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:62:3
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:65:3
	localparam [31:0] PRECISION_BITS = SUPER_MAN_BITS + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:67:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:68:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:72:3
	localparam [31:0] EXP_WIDTH = fpnew_pkg_maximum(SUPER_EXP_BITS + 2, LZC_RESULT_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:74:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 3);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:76:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:81:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:86:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:95:3
	// removed localparam type fp_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:105:3
	wire [(3 * WIDTH) - 1:0] operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:106:3
	wire [2:0] src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:107:3
	wire [2:0] dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:110:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:111:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)) + 1) * 3) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)) + 1) * 3) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3 : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3)] inp_pipe_is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:112:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:113:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:114:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:115:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:116:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:117:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:118:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:119:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:121:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:124:3
	wire [3 * WIDTH:1] sv2v_tmp_5DCC9;
	assign sv2v_tmp_5DCC9 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_5DCC9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:125:3
	wire [15:1] sv2v_tmp_7F60B;
	assign sv2v_tmp_7F60B = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] = sv2v_tmp_7F60B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:126:3
	wire [3:1] sv2v_tmp_700C1;
	assign sv2v_tmp_700C1 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_700C1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:127:3
	wire [4:1] sv2v_tmp_3923B;
	assign sv2v_tmp_3923B = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_3923B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:128:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:129:3
	wire [3:1] sv2v_tmp_6B115;
	assign sv2v_tmp_6B115 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_6B115;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:130:3
	wire [3:1] sv2v_tmp_B8677;
	assign sv2v_tmp_B8677 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_B8677;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:131:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_3F8BA;
	assign sv2v_tmp_3F8BA = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_3F8BA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:132:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_90EDD;
	assign sv2v_tmp_90EDD = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_90EDD;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:133:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:135:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:137:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] sv2v_cast_5B742;
		input reg [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] inp;
		sv2v_cast_5B742 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:139:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:143:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:145:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:145:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:145:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:145:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:147:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:149:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:149:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:149:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:149:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:150:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:150:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:150:183
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:150:291
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= (reg_ena ? inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] : inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:151:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:151:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:151:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:151:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:152:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:152:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:152:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:152:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:153:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:153:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:153:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:153:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:154:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:154:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:154:207
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:154:315
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:155:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:155:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:155:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:155:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:156:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:156:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:156:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:156:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:157:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:157:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:157:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:157:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:160:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:161:3
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:162:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:167:3
	wire [14:0] fmt_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:168:3
	wire signed [(15 * SUPER_EXP_BITS) - 1:0] fmt_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:169:3
	wire [(15 * SUPER_MAN_BITS) - 1:0] fmt_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:171:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [119:0] info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:174:3
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [SUPER_EXP_BITS - 1:0] sv2v_cast_A3BB6_signed;
		input reg signed [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_A3BB6_signed = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_52F63;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_52F63 = inp;
	endfunction
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : fmt_init_inputs
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:176:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:177:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:178:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:181:7
				wire [(3 * FP_WIDTH) - 1:0] trimmed_ops;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:184:7
				fpnew_classifier #(
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.NumOperands(3)
				) i_fpnew_classifier(
					.operands_i(trimmed_ops),
					.is_boxed_i(inp_pipe_is_boxed_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1))) * 3+:3]),
					.info_o(info_q[8 * (fmt * 3)+:24])
				);
				genvar op;
				for (op = 0; op < 3; op = op + 1) begin : gen_operands
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:193:9
					assign trimmed_ops[op * fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))+:fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH];
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:194:9
					assign fmt_sign[(fmt * 3) + op] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)];
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:195:9
					assign fmt_exponent[((fmt * 3) + op) * SUPER_EXP_BITS+:SUPER_EXP_BITS] = $signed({1'b0, operands_q[(op * WIDTH) + MAN_BITS+:EXP_BITS]});
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:196:9
					assign fmt_mantissa[((fmt * 3) + op) * SUPER_MAN_BITS+:SUPER_MAN_BITS] = {info_q[(((fmt * 3) + op) * 8) + 7], operands_q[(op * WIDTH) + (MAN_BITS - 1)-:MAN_BITS]} << (SUPER_MAN_BITS - MAN_BITS);
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:200:7
				assign info_q[8 * (fmt * 3)+:24] = {3 {sv2v_cast_8(fpnew_pkg_DONT_CARE)}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:201:7
				assign fmt_sign[fmt * 3+:3] = fpnew_pkg_DONT_CARE;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:202:7
				assign fmt_exponent[SUPER_EXP_BITS * (fmt * 3)+:SUPER_EXP_BITS * 3] = {3 {sv2v_cast_A3BB6_signed(fpnew_pkg_DONT_CARE)}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:203:7
				assign fmt_mantissa[SUPER_MAN_BITS * (fmt * 3)+:SUPER_MAN_BITS * 3] = {3 {sv2v_cast_52F63(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:207:3
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_a;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_b;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:208:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:222:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:334:40
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:335:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_A3BB6;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_A3BB6 = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_FC661;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_FC661 = inp;
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_705CC;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_705CC = inp;
	endfunction
	always @(*) begin : op_select
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:225:5
		operand_a = {fmt_sign[src_fmt_q * 3], fmt_exponent[(src_fmt_q * 3) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[(src_fmt_q * 3) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:226:5
		operand_b = {fmt_sign[(src_fmt_q * 3) + 1], fmt_exponent[((src_fmt_q * 3) + 1) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((src_fmt_q * 3) + 1) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:227:5
		operand_c = {fmt_sign[(dst_fmt_q * 3) + 2], fmt_exponent[((dst_fmt_q * 3) + 2) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((dst_fmt_q * 3) + 2) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:228:5
		info_a = info_q[(src_fmt_q * 3) * 8+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:229:5
		info_b = info_q[((src_fmt_q * 3) + 1) * 8+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:230:5
		info_c = info_q[((dst_fmt_q * 3) + 2) * 8+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:233:5
		operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:235:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(0):
				;
			sv2v_cast_A53F3(1):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:237:26
				operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = ~operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
			sv2v_cast_A53F3(2): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:239:9
				operand_a = {1'b0, sv2v_cast_A3BB6(fpnew_pkg_bias(src_fmt_q)), sv2v_cast_FC661(1'sb0)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:240:9
				info_a = 8'b10000001;
			end
			sv2v_cast_A53F3(3): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:243:9
				operand_c = {1'b1, sv2v_cast_705CC(1'sb0), sv2v_cast_FC661(1'sb0)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:244:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:247:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:248:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:249:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:250:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:251:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:252:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:260:3
	wire any_operand_inf;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:261:3
	wire any_operand_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:262:3
	wire signalling_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:263:3
	wire effective_subtraction;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:264:3
	wire tentative_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:267:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:268:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:269:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:271:3
	assign effective_subtraction = (operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))]) ^ operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:273:3
	assign tentative_sign = operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:278:3
	wire [WIDTH - 1:0] special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:279:3
	wire [4:0] special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:280:3
	wire result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:282:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:283:3
	reg [24:0] fmt_special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:284:3
	reg [4:0] fmt_result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:287:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_special_results
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:289:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:290:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:291:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:293:5
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:294:5
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:295:5
			localparam [MAN_BITS - 1:0] ZERO_MANTISSA = 1'sb0;
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:298:7
				always @(*) begin : special_results
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:299:9
					reg [FP_WIDTH - 1:0] special_res;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:302:9
					special_res = {1'b0, QNAN_EXPONENT, QNAN_MANTISSA};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:303:9
					fmt_special_status[fmt * 5+:5] = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:304:9
					fmt_result_is_special[fmt] = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:310:9
					if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:311:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:312:11
						fmt_special_status[(fmt * 5) + 4] = 1'b1;
					end
					else if (any_operand_nan) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:315:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:316:11
						fmt_special_status[(fmt * 5) + 4] = signalling_nan;
					end
					else if (any_operand_inf) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:319:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:321:11
						if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:322:13
							fmt_special_status[(fmt * 5) + 4] = 1'b1;
						else if (info_a[4] || info_b[4])
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:326:13
							special_res = {operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
						else if (info_c[4])
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:330:13
							special_res = {operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
					end
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:334:9
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:335:9
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:338:7
				wire [WIDTH * 1:1] sv2v_tmp_7740B;
				assign sv2v_tmp_7740B = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_7740B;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:339:7
				wire [5:1] sv2v_tmp_899F4;
				assign sv2v_tmp_899F4 = 1'sb0;
				always @(*) fmt_special_status[fmt * 5+:5] = sv2v_tmp_899F4;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:340:7
				wire [1:1] sv2v_tmp_77BE5;
				assign sv2v_tmp_77BE5 = 1'b0;
				always @(*) fmt_result_is_special[fmt] = sv2v_tmp_77BE5;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:345:3
	assign result_is_special = fmt_result_is_special[dst_fmt_q];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:347:3
	assign special_status = fmt_special_status[dst_fmt_q * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:349:3
	assign special_result = fmt_special_result[dst_fmt_q * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:354:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:355:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:356:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:359:3
	assign exponent_a = $signed({1'b0, operand_a[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:360:3
	assign exponent_b = $signed({1'b0, operand_b[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:361:3
	assign exponent_c = $signed({1'b0, operand_c[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:365:3
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:367:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(fpnew_pkg_bias(dst_fmt_q)) : $signed(((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - (2 * $signed(fpnew_pkg_bias(src_fmt_q)))) + $signed(fpnew_pkg_bias(dst_fmt_q))));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:374:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:376:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:379:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:381:3
	always @(*) begin : addend_shift_amount
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:383:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:384:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:387:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:390:7
			addend_shamt = 0;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:396:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:397:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:398:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:401:3
	assign mantissa_a = {info_a[7], operand_a[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:402:3
	assign mantissa_b = {info_b[7], operand_b[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:403:3
	assign mantissa_c = {info_c[7], operand_c[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:406:3
	assign product = mantissa_a * mantissa_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:411:3
	assign product_shifted = product << 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:416:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:417:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:418:3
	wire sticky_before_add;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:419:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:420:3
	wire inject_carry_in;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:430:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:433:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:436:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:437:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:442:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:443:3
	wire sum_carry;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:444:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:445:3
	wire final_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:448:3
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:449:3
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:452:3
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:455:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:463:3
	wire effective_subtraction_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:464:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:465:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:466:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:467:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:468:3
	wire sticky_before_add_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:469:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:470:3
	wire final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:471:3
	wire [2:0] dst_fmt_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:472:3
	wire [2:0] rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:473:3
	wire result_is_special_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:474:3
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] special_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:475:3
	wire [4:0] special_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:477:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:478:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:479:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:480:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:481:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:482:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:483:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:484:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:485:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:486:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:487:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:488:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) + ((NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:489:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:490:3
	reg [(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_MID_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_MID_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_MID_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_MID_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_MID_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_MID_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_MID_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] mid_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:491:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:492:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:494:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:497:3
	wire [1:1] sv2v_tmp_56A72;
	assign sv2v_tmp_56A72 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_56A72;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:498:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_8565A;
	assign sv2v_tmp_8565A = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_8565A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:499:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_F1167;
	assign sv2v_tmp_F1167 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_F1167;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:500:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_19629;
	assign sv2v_tmp_19629 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_19629;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:501:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_037F4;
	assign sv2v_tmp_037F4 = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_037F4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:502:3
	wire [1:1] sv2v_tmp_6F5F7;
	assign sv2v_tmp_6F5F7 = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6F5F7;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:503:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_74CB3;
	assign sv2v_tmp_74CB3 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_74CB3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:504:3
	wire [1:1] sv2v_tmp_D7BD0;
	assign sv2v_tmp_D7BD0 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_D7BD0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:505:3
	wire [3:1] sv2v_tmp_2170E;
	assign sv2v_tmp_2170E = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_2170E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:506:3
	wire [3:1] sv2v_tmp_8A4AE;
	assign sv2v_tmp_8A4AE = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_8A4AE;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:507:3
	wire [1:1] sv2v_tmp_7DEC5;
	assign sv2v_tmp_7DEC5 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_7DEC5;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:508:3
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) * 1:1] sv2v_tmp_1ADE6;
	assign sv2v_tmp_1ADE6 = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] = sv2v_tmp_1ADE6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:509:3
	wire [5:1] sv2v_tmp_1A1E3;
	assign sv2v_tmp_1A1E3 = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_1A1E3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:510:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_C91E0;
	assign sv2v_tmp_C91E0 = inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	always @(*) mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_C91E0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:511:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_E7982;
	assign sv2v_tmp_E7982 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_E7982;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:512:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:514:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:517:3
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:519:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:523:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:525:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:525:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:525:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:525:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:527:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:529:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:529:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:529:189
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:529:297
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:530:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:530:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:530:189
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:530:297
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:531:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:531:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:531:189
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:531:297
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:532:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:532:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:532:189
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:532:297
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:533:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:533:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:533:189
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:533:297
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:534:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:534:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:534:189
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:534:297
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:535:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:535:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:535:189
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:535:297
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:536:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:536:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:536:189
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:536:297
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:537:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:537:145
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:537:201
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:537:309
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:538:101
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:538:157
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:538:213
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:538:321
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:539:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:539:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:539:189
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:539:297
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:540:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:540:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:540:189
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:540:297
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:541:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:541:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:541:189
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:541:297
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:542:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:542:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:542:199
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:542:307
					mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:543:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:543:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:543:199
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:543:307
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:546:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:547:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:548:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:549:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:550:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:551:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:552:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:553:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:554:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:555:3
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:556:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:557:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:558:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:563:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:564:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:565:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:566:3
	wire lzc_zeroes;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:568:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:569:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:571:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:572:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:573:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:574:3
	wire sticky_after_norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:576:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:578:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:581:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:590:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:593:3
	always @(*) begin : norm_shift_amount
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:595:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:597:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:599:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:600:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:604:9
					norm_shamt = $unsigned($signed((PRECISION_BITS + 2) + exponent_product_q));
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:605:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:609:7
			norm_shamt = addend_shamt_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:610:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:615:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:619:3
	always @(*) begin : small_norm
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:621:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:622:5
		final_exponent = normalized_exponent;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:625:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:626:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:627:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:633:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:634:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:637:7
			final_exponent = 1'sb0;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:642:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:647:3
	wire pre_round_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:648:3
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:649:3
	wire [1:0] round_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:651:3
	wire of_before_round;
	wire of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:652:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:654:3
	wire [(NUM_FORMATS * (SUPER_EXP_BITS + SUPER_MAN_BITS)) - 1:0] fmt_pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:655:3
	wire [9:0] fmt_round_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:657:3
	reg [4:0] fmt_of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:658:3
	reg [4:0] fmt_uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:660:3
	wire rounded_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:661:3
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] rounded_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:662:3
	wire result_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:665:3
	assign of_before_round = final_exponent >= ((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:666:3
	assign uf_before_round = final_exponent == 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:669:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_res_assemble
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:671:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:672:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:674:5
			wire [EXP_BITS - 1:0] pre_round_exponent;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:675:5
			wire [MAN_BITS - 1:0] pre_round_mantissa;
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:679:7
				assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : final_exponent[EXP_BITS - 1:0]);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:680:7
				assign pre_round_mantissa = (of_before_round ? {fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt)) {1'sb1}} : final_mantissa[SUPER_MAN_BITS-:MAN_BITS]);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:682:7
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {pre_round_exponent, pre_round_mantissa};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:685:7
				assign fmt_round_sticky_bits[(fmt * 2) + 1] = final_mantissa[SUPER_MAN_BITS - MAN_BITS] | of_before_round;
				if (MAN_BITS < SUPER_MAN_BITS) begin : narrow_sticky
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:690:9
					assign fmt_round_sticky_bits[fmt * 2] = (|final_mantissa[(SUPER_MAN_BITS - MAN_BITS) - 1:0] | sticky_after_norm) | of_before_round;
				end
				else begin : normal_sticky
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:693:9
					assign fmt_round_sticky_bits[fmt * 2] = sticky_after_norm | of_before_round;
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:696:7
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {SUPER_EXP_BITS + SUPER_MAN_BITS {fpnew_pkg_DONT_CARE}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:697:7
				assign fmt_round_sticky_bits[fmt * 2+:2] = {2 {fpnew_pkg_DONT_CARE}};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:702:3
	assign pre_round_sign = final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:703:3
	assign pre_round_abs = fmt_pre_round_abs[dst_fmt_q2 * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:706:3
	assign round_sticky_bits = fmt_round_sticky_bits[dst_fmt_q2 * 2+:2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:709:3
	fpnew_rounding #(.AbsWidth(SUPER_EXP_BITS + SUPER_MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:722:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:724:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_sign_inject
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:726:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:727:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:728:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:731:7
				always @(*) begin : post_process
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:733:9
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:734:9
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:737:9
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:738:9
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]};
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:741:7
				wire [1:1] sv2v_tmp_4A747;
				assign sv2v_tmp_4A747 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4A747;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:742:7
				wire [1:1] sv2v_tmp_90681;
				assign sv2v_tmp_90681 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_90681;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:743:7
				wire [WIDTH * 1:1] sv2v_tmp_143A7;
				assign sv2v_tmp_143A7 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_143A7;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:748:3
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:749:3
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:755:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:756:3
	wire [4:0] regular_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:759:3
	assign regular_result = fmt_result[dst_fmt_q2 * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:760:3
	assign regular_status[4] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:761:3
	assign regular_status[3] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:762:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:763:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:764:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:767:3
	wire [WIDTH - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:768:3
	wire [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:771:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:772:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:778:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:779:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:780:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:781:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:782:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:784:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:787:3
	wire [WIDTH * 1:1] sv2v_tmp_1212D;
	assign sv2v_tmp_1212D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_1212D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:788:3
	wire [5:1] sv2v_tmp_F691B;
	assign sv2v_tmp_F691B = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_F691B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:789:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_95B09;
	assign sv2v_tmp_95B09 = mid_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_95B09;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:790:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_E2659;
	assign sv2v_tmp_E2659 = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_E2659;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:791:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:793:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:795:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:797:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:801:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:803:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:803:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:803:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:803:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:805:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:807:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:807:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:807:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:807:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:808:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:808:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:808:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:808:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:809:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:809:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:809:189
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:809:297
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:810:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:810:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:810:189
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:810:297
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:813:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:815:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:816:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:817:3
	assign extension_bit_o = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:818:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:819:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:820:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:821:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_fma_multi_7F4A8_72E9B (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type AuxType_AUX_BITS_type
	parameter [31:0] AuxType_AUX_BITS = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:18:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:19:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:20:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:21:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:23:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:306:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:307:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:310:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:24:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:26:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:27:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:29:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:30:3
	input wire [14:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:31:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:32:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:33:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:34:3
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:35:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:36:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:37:3
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:39:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:40:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:41:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:43:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:44:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:45:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:46:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:47:3
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:49:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:50:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:52:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:59:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:338:49
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:339:5
		reg [63:0] res;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:340:5
			res = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:5
			begin : sv2v_autoblock_2
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:10
				reg [31:0] fmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:341:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:343:9
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt))));
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:344:9
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:61:3
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:62:3
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:65:3
	localparam [31:0] PRECISION_BITS = SUPER_MAN_BITS + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:67:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:68:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:72:3
	localparam [31:0] EXP_WIDTH = fpnew_pkg_maximum(SUPER_EXP_BITS + 2, LZC_RESULT_WIDTH);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:74:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 3);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:76:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:81:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:86:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:95:3
	// removed localparam type fp_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:105:3
	wire [(3 * WIDTH) - 1:0] operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:106:3
	wire [2:0] src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:107:3
	wire [2:0] dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:110:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:111:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)) + 1) * 3) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)) + 1) * 3) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3 : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3)] inp_pipe_is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:112:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:113:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:114:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:115:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:116:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:117:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:118:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:119:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:121:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:124:3
	wire [3 * WIDTH:1] sv2v_tmp_5DCC9;
	assign sv2v_tmp_5DCC9 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_5DCC9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:125:3
	wire [15:1] sv2v_tmp_7F60B;
	assign sv2v_tmp_7F60B = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] = sv2v_tmp_7F60B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:126:3
	wire [3:1] sv2v_tmp_700C1;
	assign sv2v_tmp_700C1 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_700C1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:127:3
	wire [4:1] sv2v_tmp_3923B;
	assign sv2v_tmp_3923B = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_3923B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:128:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:129:3
	wire [3:1] sv2v_tmp_6B115;
	assign sv2v_tmp_6B115 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_6B115;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:130:3
	wire [3:1] sv2v_tmp_B8677;
	assign sv2v_tmp_B8677 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_B8677;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:131:3
	wire [1:1] sv2v_tmp_76699;
	assign sv2v_tmp_76699 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_76699;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:132:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_61815;
	assign sv2v_tmp_61815 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_61815;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:133:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:135:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:137:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:139:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:143:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:145:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:145:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:145:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:145:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:147:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:149:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:149:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:149:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:149:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:150:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:150:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:150:183
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:150:291
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= (reg_ena ? inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] : inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:151:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:151:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:151:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:151:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:152:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:152:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:152:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:152:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:153:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:153:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:153:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:153:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:154:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:154:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:154:207
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:154:315
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:155:95
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:155:151
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:155:207
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:155:315
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:156:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:156:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:156:193
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:156:301
					inp_pipe_tag_q[i + 1] <= (reg_ena ? inp_pipe_tag_q[i] : inp_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:157:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:157:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:157:193
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:157:301
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:160:3
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:161:3
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:162:3
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:167:3
	wire [14:0] fmt_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:168:3
	wire signed [(15 * SUPER_EXP_BITS) - 1:0] fmt_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:169:3
	wire [(15 * SUPER_MAN_BITS) - 1:0] fmt_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:171:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [119:0] info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:174:3
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [SUPER_EXP_BITS - 1:0] sv2v_cast_A3BB6_signed;
		input reg signed [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_A3BB6_signed = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_52F63;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_52F63 = inp;
	endfunction
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : fmt_init_inputs
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:176:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:177:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:178:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:181:7
				wire [(3 * FP_WIDTH) - 1:0] trimmed_ops;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:184:7
				fpnew_classifier #(
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.NumOperands(3)
				) i_fpnew_classifier(
					.operands_i(trimmed_ops),
					.is_boxed_i(inp_pipe_is_boxed_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1))) * 3+:3]),
					.info_o(info_q[8 * (fmt * 3)+:24])
				);
				genvar op;
				for (op = 0; op < 3; op = op + 1) begin : gen_operands
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:193:9
					assign trimmed_ops[op * fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))+:fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH];
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:194:9
					assign fmt_sign[(fmt * 3) + op] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)];
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:195:9
					assign fmt_exponent[((fmt * 3) + op) * SUPER_EXP_BITS+:SUPER_EXP_BITS] = $signed({1'b0, operands_q[(op * WIDTH) + MAN_BITS+:EXP_BITS]});
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:196:9
					assign fmt_mantissa[((fmt * 3) + op) * SUPER_MAN_BITS+:SUPER_MAN_BITS] = {info_q[(((fmt * 3) + op) * 8) + 7], operands_q[(op * WIDTH) + (MAN_BITS - 1)-:MAN_BITS]} << (SUPER_MAN_BITS - MAN_BITS);
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:200:7
				assign info_q[8 * (fmt * 3)+:24] = {3 {sv2v_cast_8(fpnew_pkg_DONT_CARE)}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:201:7
				assign fmt_sign[fmt * 3+:3] = fpnew_pkg_DONT_CARE;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:202:7
				assign fmt_exponent[SUPER_EXP_BITS * (fmt * 3)+:SUPER_EXP_BITS * 3] = {3 {sv2v_cast_A3BB6_signed(fpnew_pkg_DONT_CARE)}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:203:7
				assign fmt_mantissa[SUPER_MAN_BITS * (fmt * 3)+:SUPER_MAN_BITS * 3] = {3 {sv2v_cast_52F63(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:207:3
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_a;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_b;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:208:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:222:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:334:40
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:335:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_A3BB6;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_A3BB6 = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_FC661;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_FC661 = inp;
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_705CC;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_705CC = inp;
	endfunction
	always @(*) begin : op_select
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:225:5
		operand_a = {fmt_sign[src_fmt_q * 3], fmt_exponent[(src_fmt_q * 3) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[(src_fmt_q * 3) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:226:5
		operand_b = {fmt_sign[(src_fmt_q * 3) + 1], fmt_exponent[((src_fmt_q * 3) + 1) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((src_fmt_q * 3) + 1) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:227:5
		operand_c = {fmt_sign[(dst_fmt_q * 3) + 2], fmt_exponent[((dst_fmt_q * 3) + 2) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((dst_fmt_q * 3) + 2) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:228:5
		info_a = info_q[(src_fmt_q * 3) * 8+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:229:5
		info_b = info_q[((src_fmt_q * 3) + 1) * 8+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:230:5
		info_c = info_q[((dst_fmt_q * 3) + 2) * 8+:8];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:233:5
		operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:235:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(0):
				;
			sv2v_cast_A53F3(1):
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:237:26
				operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = ~operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
			sv2v_cast_A53F3(2): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:239:9
				operand_a = {1'b0, sv2v_cast_A3BB6(fpnew_pkg_bias(src_fmt_q)), sv2v_cast_FC661(1'sb0)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:240:9
				info_a = 8'b10000001;
			end
			sv2v_cast_A53F3(3): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:243:9
				operand_c = {1'b1, sv2v_cast_705CC(1'sb0), sv2v_cast_FC661(1'sb0)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:244:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:247:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:248:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:249:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:250:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:251:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:252:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:260:3
	wire any_operand_inf;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:261:3
	wire any_operand_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:262:3
	wire signalling_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:263:3
	wire effective_subtraction;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:264:3
	wire tentative_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:267:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:268:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:269:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:271:3
	assign effective_subtraction = (operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))]) ^ operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:273:3
	assign tentative_sign = operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:278:3
	wire [WIDTH - 1:0] special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:279:3
	wire [4:0] special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:280:3
	wire result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:282:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:283:3
	reg [24:0] fmt_special_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:284:3
	reg [4:0] fmt_result_is_special;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:287:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_special_results
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:289:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:290:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:291:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:293:5
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:294:5
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:295:5
			localparam [MAN_BITS - 1:0] ZERO_MANTISSA = 1'sb0;
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:298:7
				always @(*) begin : special_results
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:299:9
					reg [FP_WIDTH - 1:0] special_res;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:302:9
					special_res = {1'b0, QNAN_EXPONENT, QNAN_MANTISSA};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:303:9
					fmt_special_status[fmt * 5+:5] = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:304:9
					fmt_result_is_special[fmt] = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:310:9
					if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:311:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:312:11
						fmt_special_status[(fmt * 5) + 4] = 1'b1;
					end
					else if (any_operand_nan) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:315:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:316:11
						fmt_special_status[(fmt * 5) + 4] = signalling_nan;
					end
					else if (any_operand_inf) begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:319:11
						fmt_result_is_special[fmt] = 1'b1;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:321:11
						if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:322:13
							fmt_special_status[(fmt * 5) + 4] = 1'b1;
						else if (info_a[4] || info_b[4])
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:326:13
							special_res = {operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
						else if (info_c[4])
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:330:13
							special_res = {operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
					end
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:334:9
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:335:9
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:338:7
				wire [WIDTH * 1:1] sv2v_tmp_7740B;
				assign sv2v_tmp_7740B = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_7740B;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:339:7
				wire [5:1] sv2v_tmp_899F4;
				assign sv2v_tmp_899F4 = 1'sb0;
				always @(*) fmt_special_status[fmt * 5+:5] = sv2v_tmp_899F4;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:340:7
				wire [1:1] sv2v_tmp_77BE5;
				assign sv2v_tmp_77BE5 = 1'b0;
				always @(*) fmt_result_is_special[fmt] = sv2v_tmp_77BE5;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:345:3
	assign result_is_special = fmt_result_is_special[dst_fmt_q];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:347:3
	assign special_status = fmt_special_status[dst_fmt_q * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:349:3
	assign special_result = fmt_special_result[dst_fmt_q * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:354:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:355:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:356:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:359:3
	assign exponent_a = $signed({1'b0, operand_a[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:360:3
	assign exponent_b = $signed({1'b0, operand_b[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:361:3
	assign exponent_c = $signed({1'b0, operand_c[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:365:3
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:367:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(fpnew_pkg_bias(dst_fmt_q)) : $signed(((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - (2 * $signed(fpnew_pkg_bias(src_fmt_q)))) + $signed(fpnew_pkg_bias(dst_fmt_q))));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:374:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:376:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:379:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:381:3
	always @(*) begin : addend_shift_amount
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:383:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:384:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:387:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:390:7
			addend_shamt = 0;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:396:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:397:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:398:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:401:3
	assign mantissa_a = {info_a[7], operand_a[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:402:3
	assign mantissa_b = {info_b[7], operand_b[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:403:3
	assign mantissa_c = {info_c[7], operand_c[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:406:3
	assign product = mantissa_a * mantissa_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:411:3
	assign product_shifted = product << 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:416:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:417:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:418:3
	wire sticky_before_add;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:419:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:420:3
	wire inject_carry_in;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:430:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:433:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:436:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:437:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:442:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:443:3
	wire sum_carry;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:444:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:445:3
	wire final_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:448:3
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:449:3
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:452:3
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:455:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:463:3
	wire effective_subtraction_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:464:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:465:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:466:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:467:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:468:3
	wire sticky_before_add_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:469:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:470:3
	wire final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:471:3
	wire [2:0] dst_fmt_q2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:472:3
	wire [2:0] rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:473:3
	wire result_is_special_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:474:3
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] special_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:475:3
	wire [4:0] special_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:477:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:478:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:479:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:480:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:481:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:482:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:483:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:484:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:485:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:486:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:487:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:488:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) + ((NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:489:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:490:3
	reg [0:NUM_MID_REGS] mid_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:491:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:492:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:494:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:497:3
	wire [1:1] sv2v_tmp_56A72;
	assign sv2v_tmp_56A72 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_56A72;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:498:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_8565A;
	assign sv2v_tmp_8565A = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_8565A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:499:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_F1167;
	assign sv2v_tmp_F1167 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_F1167;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:500:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_19629;
	assign sv2v_tmp_19629 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_19629;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:501:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_037F4;
	assign sv2v_tmp_037F4 = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_037F4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:502:3
	wire [1:1] sv2v_tmp_6F5F7;
	assign sv2v_tmp_6F5F7 = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6F5F7;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:503:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_74CB3;
	assign sv2v_tmp_74CB3 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_74CB3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:504:3
	wire [1:1] sv2v_tmp_D7BD0;
	assign sv2v_tmp_D7BD0 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_D7BD0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:505:3
	wire [3:1] sv2v_tmp_2170E;
	assign sv2v_tmp_2170E = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_2170E;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:506:3
	wire [3:1] sv2v_tmp_8A4AE;
	assign sv2v_tmp_8A4AE = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_8A4AE;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:507:3
	wire [1:1] sv2v_tmp_7DEC5;
	assign sv2v_tmp_7DEC5 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_7DEC5;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:508:3
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) * 1:1] sv2v_tmp_1ADE6;
	assign sv2v_tmp_1ADE6 = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] = sv2v_tmp_1ADE6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:509:3
	wire [5:1] sv2v_tmp_1A1E3;
	assign sv2v_tmp_1A1E3 = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_1A1E3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:510:3
	wire [1:1] sv2v_tmp_44BCE;
	assign sv2v_tmp_44BCE = inp_pipe_tag_q[NUM_INP_REGS];
	always @(*) mid_pipe_tag_q[0] = sv2v_tmp_44BCE;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:511:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_723C6;
	assign sv2v_tmp_723C6 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_723C6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:512:3
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:514:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:517:3
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:519:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:523:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:525:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:525:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:525:408
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:525:560
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:527:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:529:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:529:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:529:189
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:529:297
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:530:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:530:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:530:189
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:530:297
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:531:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:531:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:531:189
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:531:297
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:532:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:532:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:532:189
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:532:297
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:533:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:533:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:533:189
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:533:297
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:534:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:534:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:534:189
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:534:297
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:535:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:535:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:535:189
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:535:297
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:536:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:536:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:536:189
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:536:297
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:537:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:537:145
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:537:201
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:537:309
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:538:101
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:538:157
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:538:213
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:538:321
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:539:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:539:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:539:189
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:539:297
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:540:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:540:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:540:189
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:540:297
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:541:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:541:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:541:189
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:541:297
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:542:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:542:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:542:199
					mid_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:542:307
					mid_pipe_tag_q[i + 1] <= (reg_ena ? mid_pipe_tag_q[i] : mid_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:543:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:543:143
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:543:199
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:543:307
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:546:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:547:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:548:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:549:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:550:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:551:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:552:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:553:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:554:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:555:3
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:556:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:557:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:558:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:563:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:564:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:565:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:566:3
	wire lzc_zeroes;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:568:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:569:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:571:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:572:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:573:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:574:3
	wire sticky_after_norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:576:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:578:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:581:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:590:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:593:3
	always @(*) begin : norm_shift_amount
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:595:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:597:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:599:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:600:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:604:9
					norm_shamt = $unsigned($signed((PRECISION_BITS + 2) + exponent_product_q));
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:605:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:609:7
			norm_shamt = addend_shamt_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:610:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:615:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:619:3
	always @(*) begin : small_norm
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:621:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:622:5
		final_exponent = normalized_exponent;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:625:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:626:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:627:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:633:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:634:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:637:7
			final_exponent = 1'sb0;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:642:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:647:3
	wire pre_round_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:648:3
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:649:3
	wire [1:0] round_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:651:3
	wire of_before_round;
	wire of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:652:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:654:3
	wire [(NUM_FORMATS * (SUPER_EXP_BITS + SUPER_MAN_BITS)) - 1:0] fmt_pre_round_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:655:3
	wire [9:0] fmt_round_sticky_bits;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:657:3
	reg [4:0] fmt_of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:658:3
	reg [4:0] fmt_uf_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:660:3
	wire rounded_sign;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:661:3
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] rounded_abs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:662:3
	wire result_zero;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:665:3
	assign of_before_round = final_exponent >= ((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:666:3
	assign uf_before_round = final_exponent == 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:669:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_res_assemble
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:671:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:672:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:674:5
			wire [EXP_BITS - 1:0] pre_round_exponent;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:675:5
			wire [MAN_BITS - 1:0] pre_round_mantissa;
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:679:7
				assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : final_exponent[EXP_BITS - 1:0]);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:680:7
				assign pre_round_mantissa = (of_before_round ? {fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt)) {1'sb1}} : final_mantissa[SUPER_MAN_BITS-:MAN_BITS]);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:682:7
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {pre_round_exponent, pre_round_mantissa};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:685:7
				assign fmt_round_sticky_bits[(fmt * 2) + 1] = final_mantissa[SUPER_MAN_BITS - MAN_BITS] | of_before_round;
				if (MAN_BITS < SUPER_MAN_BITS) begin : narrow_sticky
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:690:9
					assign fmt_round_sticky_bits[fmt * 2] = (|final_mantissa[(SUPER_MAN_BITS - MAN_BITS) - 1:0] | sticky_after_norm) | of_before_round;
				end
				else begin : normal_sticky
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:693:9
					assign fmt_round_sticky_bits[fmt * 2] = sticky_after_norm | of_before_round;
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:696:7
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {SUPER_EXP_BITS + SUPER_MAN_BITS {fpnew_pkg_DONT_CARE}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:697:7
				assign fmt_round_sticky_bits[fmt * 2+:2] = {2 {fpnew_pkg_DONT_CARE}};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:702:3
	assign pre_round_sign = final_sign_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:703:3
	assign pre_round_abs = fmt_pre_round_abs[dst_fmt_q2 * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:706:3
	assign round_sticky_bits = fmt_round_sticky_bits[dst_fmt_q2 * 2+:2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:709:3
	fpnew_rounding #(.AbsWidth(SUPER_EXP_BITS + SUPER_MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:722:3
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:724:3
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_sign_inject
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:726:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:727:5
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:728:5
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:731:7
				always @(*) begin : post_process
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:733:9
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:734:9
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:737:9
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:738:9
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]};
				end
			end
			else begin : inactive_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:741:7
				wire [1:1] sv2v_tmp_4A747;
				assign sv2v_tmp_4A747 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4A747;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:742:7
				wire [1:1] sv2v_tmp_90681;
				assign sv2v_tmp_90681 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_90681;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:743:7
				wire [WIDTH * 1:1] sv2v_tmp_143A7;
				assign sv2v_tmp_143A7 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_143A7;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:748:3
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:749:3
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:755:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:756:3
	wire [4:0] regular_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:759:3
	assign regular_result = fmt_result[dst_fmt_q2 * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:760:3
	assign regular_status[4] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:761:3
	assign regular_status[3] = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:762:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:763:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:764:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:767:3
	wire [WIDTH - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:768:3
	wire [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:771:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:772:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:778:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:779:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:780:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:781:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:782:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:784:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:787:3
	wire [WIDTH * 1:1] sv2v_tmp_1212D;
	assign sv2v_tmp_1212D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_1212D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:788:3
	wire [5:1] sv2v_tmp_F691B;
	assign sv2v_tmp_F691B = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_F691B;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:789:3
	wire [1:1] sv2v_tmp_DF7DA;
	assign sv2v_tmp_DF7DA = mid_pipe_tag_q[NUM_MID_REGS];
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_DF7DA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:790:3
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_F2485;
	assign sv2v_tmp_F2485 = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_F2485;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:791:3
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:793:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:795:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:797:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:801:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:803:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:803:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:803:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:803:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:805:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:807:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:807:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:807:179
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:807:287
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:808:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:808:123
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:808:179
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:808:287
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:809:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:809:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:809:189
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:809:297
					out_pipe_tag_q[i + 1] <= (reg_ena ? out_pipe_tag_q[i] : out_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:810:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:810:133
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:810:189
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:810:297
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:813:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:815:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:816:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:817:3
	assign extension_bit_o = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:818:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:819:3
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:820:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_fma_multi.sv:821:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_noncomp_1F07E (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	class_mask_o,
	is_class_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:18:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:19:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:20:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:21:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:23:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:25:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:26:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:28:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:29:3
	input wire [1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:30:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:31:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:32:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:33:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:34:3
	input wire aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:36:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:37:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:38:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:40:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:41:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:42:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:43:3
	// removed localparam type fpnew_pkg_classmask_e
	output wire [9:0] class_mask_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:44:3
	output wire is_class_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:45:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:46:3
	output wire aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:48:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:49:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:51:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:57:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:58:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:60:3
	localparam NUM_INP_REGS = ((PipeConfig == 2'd0) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:65:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:74:3
	// removed localparam type fp_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:84:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:85:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)] inp_pipe_is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:86:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:87:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:88:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:89:3
	reg [0:NUM_INP_REGS] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:90:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:91:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:93:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:96:3
	wire [2 * WIDTH:1] sv2v_tmp_D1067;
	assign sv2v_tmp_D1067 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_D1067;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:97:3
	wire [2:1] sv2v_tmp_86D63;
	assign sv2v_tmp_86D63 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2+:2] = sv2v_tmp_86D63;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:98:3
	wire [3:1] sv2v_tmp_62109;
	assign sv2v_tmp_62109 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_62109;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:99:3
	wire [4:1] sv2v_tmp_0B797;
	assign sv2v_tmp_0B797 = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_0B797;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:100:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:101:3
	wire [1:1] sv2v_tmp_76699;
	assign sv2v_tmp_76699 = tag_i;
	always @(*) inp_pipe_tag_q[0] = sv2v_tmp_76699;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:102:3
	wire [1:1] sv2v_tmp_8D189;
	assign sv2v_tmp_8D189 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_8D189;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:103:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:105:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:107:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:109:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:113:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:115:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:115:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:115:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:115:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:117:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:119:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:119:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:119:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:119:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:120:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:120:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:120:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:120:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2+:2] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:121:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:121:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:121:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:121:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:122:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:122:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:122:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:122:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:123:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:123:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:123:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:123:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:124:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:124:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:124:193
					inp_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:124:301
					inp_pipe_tag_q[i + 1] <= (reg_ena ? inp_pipe_tag_q[i] : inp_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:125:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:125:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:125:193
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:125:301
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:131:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [15:0] info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:134:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(2)
	) i_class_a(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2+:2]),
		.info_o(info_q)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:143:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:144:3
	wire [7:0] info_a;
	wire [7:0] info_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:147:3
	assign operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:148:3
	assign operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:149:3
	assign info_a = info_q[0+:8];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:150:3
	assign info_b = info_q[8+:8];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:152:3
	wire any_operand_inf;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:153:3
	wire any_operand_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:154:3
	wire signalling_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:157:3
	assign any_operand_inf = |{info_a[4], info_b[4]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:158:3
	assign any_operand_nan = |{info_a[3], info_b[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:159:3
	assign signalling_nan = |{info_a[2], info_b[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:161:3
	wire operands_equal;
	wire operand_a_smaller;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:164:3
	assign operands_equal = (operand_a == operand_b) || (info_a[5] && info_b[5]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:166:3
	assign operand_a_smaller = (operand_a < operand_b) ^ (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] || operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:171:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] sgnj_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:172:3
	wire [4:0] sgnj_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:173:3
	wire sgnj_extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:177:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_F2D56;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_F2D56 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_14681;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_14681 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_91364;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_91364 = inp;
	endfunction
	always @(*) begin : sign_injections
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:178:5
		reg sign_a;
		reg sign_b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:180:5
		sgnj_result = operand_a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:183:5
		if (!info_a[0])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:183:27
			sgnj_result = {1'b0, sv2v_cast_F2D56(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:186:5
		sign_a = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] & info_a[0];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:187:5
		sign_b = operand_b[1 + (EXP_BITS + (MAN_BITS - 1))] & info_b[0];
		case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
			3'b000:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:191:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_b;
			3'b001:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:192:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = ~sign_b;
			3'b010:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:193:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_a ^ sign_b;
			3'b011:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:194:23
				sgnj_result = operand_a;
			default:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:195:16
				sgnj_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:199:3
	assign sgnj_status = 1'sb0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:202:3
	assign sgnj_extension_bit = (inp_pipe_op_mod_q[NUM_INP_REGS] ? sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] : 1'b1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:207:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] minmax_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:208:3
	reg [4:0] minmax_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:209:3
	wire minmax_extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:213:3
	always @(*) begin : min_max
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:215:5
		minmax_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:218:5
		minmax_status[4] = signalling_nan;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:221:5
		if (info_a[3] && info_b[3])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:222:7
			minmax_result = {1'b0, sv2v_cast_F2D56(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		else if (info_a[3])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:224:29
			minmax_result = operand_b;
		else if (info_b[3])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:225:29
			minmax_result = operand_a;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:228:7
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:229:25
					minmax_result = (operand_a_smaller ? operand_a : operand_b);
				3'b001:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:230:25
					minmax_result = (operand_a_smaller ? operand_b : operand_a);
				default:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:231:18
					minmax_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
			endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:236:3
	assign minmax_extension_bit = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:241:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] cmp_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:242:3
	reg [4:0] cmp_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:243:3
	wire cmp_extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:248:3
	always @(*) begin : comparisons
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:250:5
		cmp_result = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:251:5
		cmp_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:254:5
		if (signalling_nan)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:254:25
			cmp_status[4] = 1'b1;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:257:7
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:259:11
					if (any_operand_nan)
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:259:32
						cmp_status[4] = 1'b1;
					else
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:260:16
						cmp_result = (operand_a_smaller | operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b001:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:263:11
					if (any_operand_nan)
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:263:32
						cmp_status[4] = 1'b1;
					else
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:264:16
						cmp_result = (operand_a_smaller & ~operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b010:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:267:11
					if (any_operand_nan)
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:267:32
						cmp_result = inp_pipe_op_mod_q[NUM_INP_REGS];
					else
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:268:16
						cmp_result = operands_equal ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				default:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:270:18
					cmp_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
			endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:275:3
	assign cmp_extension_bit = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:280:3
	wire [4:0] class_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:281:3
	wire class_extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:282:3
	reg [9:0] class_mask_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:285:3
	always @(*) begin : classify
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:286:5
		if (info_a[7])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:287:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000010 : 10'b0001000000);
		else if (info_a[6])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:289:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000100 : 10'b0000100000);
		else if (info_a[5])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:291:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000001000 : 10'b0000010000);
		else if (info_a[4])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:293:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000001 : 10'b0010000000);
		else if (info_a[3])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:295:7
			class_mask_d = (info_a[2] ? 10'b0100000000 : 10'b1000000000);
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:297:7
			class_mask_d = 10'b1000000000;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:301:3
	assign class_status = 1'sb0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:302:3
	assign class_extension_bit = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:307:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:308:3
	reg [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:309:3
	reg extension_bit_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:310:3
	wire is_class_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:313:3
	always @(*) begin : select_result
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:314:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(6): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:316:9
				result_d = sgnj_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:317:9
				status_d = sgnj_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:318:9
				extension_bit_d = sgnj_extension_bit;
			end
			sv2v_cast_A53F3(7): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:321:9
				result_d = minmax_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:322:9
				status_d = minmax_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:323:9
				extension_bit_d = minmax_extension_bit;
			end
			sv2v_cast_A53F3(8): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:326:9
				result_d = cmp_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:327:9
				status_d = cmp_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:328:9
				extension_bit_d = cmp_extension_bit;
			end
			sv2v_cast_A53F3(9): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:331:9
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:332:9
				status_d = class_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:333:9
				extension_bit_d = class_extension_bit;
			end
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:336:9
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:337:9
				status_d = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:338:9
				extension_bit_d = fpnew_pkg_DONT_CARE;
			end
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:343:3
	assign is_class_d = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(9);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:349:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:350:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:351:3
	reg [0:NUM_OUT_REGS] out_pipe_extension_bit_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:352:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 10) + ((NUM_OUT_REGS * 10) - 1) : ((NUM_OUT_REGS + 1) * 10) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 10 : 0)] out_pipe_class_mask_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:353:3
	reg [0:NUM_OUT_REGS] out_pipe_is_class_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:354:3
	reg [0:NUM_OUT_REGS] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:355:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:356:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:358:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:361:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_07494;
	assign sv2v_tmp_07494 = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_07494;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:362:3
	wire [5:1] sv2v_tmp_CCE43;
	assign sv2v_tmp_CCE43 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_CCE43;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:363:3
	wire [1:1] sv2v_tmp_8E9A9;
	assign sv2v_tmp_8E9A9 = extension_bit_d;
	always @(*) out_pipe_extension_bit_q[0] = sv2v_tmp_8E9A9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:364:3
	wire [10:1] sv2v_tmp_94259;
	assign sv2v_tmp_94259 = class_mask_d;
	always @(*) out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 10+:10] = sv2v_tmp_94259;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:365:3
	wire [1:1] sv2v_tmp_7DF01;
	assign sv2v_tmp_7DF01 = is_class_d;
	always @(*) out_pipe_is_class_q[0] = sv2v_tmp_7DF01;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:366:3
	wire [1:1] sv2v_tmp_35518;
	assign sv2v_tmp_35518 = inp_pipe_tag_q[NUM_INP_REGS];
	always @(*) out_pipe_tag_q[0] = sv2v_tmp_35518;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:367:3
	wire [1:1] sv2v_tmp_FA930;
	assign sv2v_tmp_FA930 = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_FA930;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:368:3
	wire [1:1] sv2v_tmp_2CB8C;
	assign sv2v_tmp_2CB8C = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_2CB8C;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:370:3
	assign inp_pipe_ready[NUM_INP_REGS] = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:372:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:374:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:378:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:380:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:380:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:380:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:380:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:382:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:384:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:384:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:384:193
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:384:301
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:385:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:385:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:385:193
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:385:301
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:386:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:386:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:386:193
					out_pipe_extension_bit_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:386:301
					out_pipe_extension_bit_q[i + 1] <= (reg_ena ? out_pipe_extension_bit_q[i] : out_pipe_extension_bit_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:387:94
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:387:150
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:387:206
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= 10'b1000000000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:387:314
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= (reg_ena ? out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 10+:10] : out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:388:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:388:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:388:193
					out_pipe_is_class_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:388:301
					out_pipe_is_class_q[i + 1] <= (reg_ena ? out_pipe_is_class_q[i] : out_pipe_is_class_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:389:91
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:389:147
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:389:203
					out_pipe_tag_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:389:311
					out_pipe_tag_q[i + 1] <= (reg_ena ? out_pipe_tag_q[i] : out_pipe_tag_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:390:91
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:390:147
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:390:203
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:390:311
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:393:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:395:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:396:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:397:3
	assign extension_bit_o = out_pipe_extension_bit_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:398:3
	assign class_mask_o = out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 10+:10];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:399:3
	assign is_class_o = out_pipe_is_class_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:400:3
	assign tag_o = out_pipe_tag_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:401:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:402:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:403:3
	assign busy_o = |{inp_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_noncomp_546BA_F0963 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	class_mask_o,
	is_class_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TagType_TagType_TagType_TAGW_type
	parameter signed [31:0] TagType_TagType_TagType_TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:17:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:18:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:19:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:20:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:21:38
	// removed localparam type AuxType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:23:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:25:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:26:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:28:3
	input wire [(2 * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:29:3
	input wire [1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:30:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:31:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:32:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:33:3
	input wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:34:3
	input wire aux_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:36:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:37:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:38:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:40:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:41:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:42:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:43:3
	// removed localparam type fpnew_pkg_classmask_e
	output wire [9:0] class_mask_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:44:3
	output wire is_class_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:45:3
	output wire [TagType_TagType_TagType_TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:46:3
	output wire aux_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:48:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:49:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:51:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:57:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:324:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:325:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:58:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:329:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:330:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:60:3
	localparam NUM_INP_REGS = ((PipeConfig == 2'd0) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:65:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:74:3
	// removed localparam type fp_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:84:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:85:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)] inp_pipe_is_boxed_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:86:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:87:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:88:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:89:3
	reg [(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_INP_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_INP_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_INP_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_INP_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_INP_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_INP_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_INP_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] inp_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:90:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:91:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:93:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:96:3
	wire [2 * WIDTH:1] sv2v_tmp_D1067;
	assign sv2v_tmp_D1067 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_D1067;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:97:3
	wire [2:1] sv2v_tmp_86D63;
	assign sv2v_tmp_86D63 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2+:2] = sv2v_tmp_86D63;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:98:3
	wire [3:1] sv2v_tmp_62109;
	assign sv2v_tmp_62109 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_62109;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:99:3
	wire [4:1] sv2v_tmp_0B797;
	assign sv2v_tmp_0B797 = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_0B797;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:100:3
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:101:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_2696A;
	assign sv2v_tmp_2696A = tag_i;
	always @(*) inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_2696A;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:102:3
	wire [1:1] sv2v_tmp_8D189;
	assign sv2v_tmp_8D189 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_8D189;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:103:3
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:105:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:107:3
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] sv2v_cast_5B742;
		input reg [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) - 1:0] inp;
		sv2v_cast_5B742 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:109:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:113:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:115:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:115:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:115:408
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:115:560
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:117:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:119:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:119:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:119:183
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:119:291
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:120:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:120:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:120:183
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:120:291
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2+:2] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:121:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:121:139
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:121:195
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:121:303
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:122:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:122:141
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:122:197
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:122:305
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:123:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:123:127
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:123:183
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:123:291
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:124:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:124:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:124:193
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:124:301
					inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:125:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:125:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:125:193
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:125:301
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:131:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [15:0] info_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:134:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(2)
	) i_class_a(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2+:2]),
		.info_o(info_q)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:143:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:144:3
	wire [7:0] info_a;
	wire [7:0] info_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:147:3
	assign operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:148:3
	assign operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:149:3
	assign info_a = info_q[0+:8];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:150:3
	assign info_b = info_q[8+:8];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:152:3
	wire any_operand_inf;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:153:3
	wire any_operand_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:154:3
	wire signalling_nan;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:157:3
	assign any_operand_inf = |{info_a[4], info_b[4]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:158:3
	assign any_operand_nan = |{info_a[3], info_b[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:159:3
	assign signalling_nan = |{info_a[2], info_b[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:161:3
	wire operands_equal;
	wire operand_a_smaller;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:164:3
	assign operands_equal = (operand_a == operand_b) || (info_a[5] && info_b[5]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:166:3
	assign operand_a_smaller = (operand_a < operand_b) ^ (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] || operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:171:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] sgnj_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:172:3
	wire [4:0] sgnj_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:173:3
	wire sgnj_extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:177:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_F2D56;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_F2D56 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_14681;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_14681 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_91364;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_91364 = inp;
	endfunction
	always @(*) begin : sign_injections
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:178:5
		reg sign_a;
		reg sign_b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:180:5
		sgnj_result = operand_a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:183:5
		if (!info_a[0])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:183:27
			sgnj_result = {1'b0, sv2v_cast_F2D56(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:186:5
		sign_a = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] & info_a[0];
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:187:5
		sign_b = operand_b[1 + (EXP_BITS + (MAN_BITS - 1))] & info_b[0];
		case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
			3'b000:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:191:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_b;
			3'b001:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:192:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = ~sign_b;
			3'b010:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:193:23
				sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_a ^ sign_b;
			3'b011:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:194:23
				sgnj_result = operand_a;
			default:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:195:16
				sgnj_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:199:3
	assign sgnj_status = 1'sb0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:202:3
	assign sgnj_extension_bit = (inp_pipe_op_mod_q[NUM_INP_REGS] ? sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] : 1'b1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:207:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] minmax_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:208:3
	reg [4:0] minmax_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:209:3
	wire minmax_extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:213:3
	always @(*) begin : min_max
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:215:5
		minmax_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:218:5
		minmax_status[4] = signalling_nan;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:221:5
		if (info_a[3] && info_b[3])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:222:7
			minmax_result = {1'b0, sv2v_cast_F2D56(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		else if (info_a[3])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:224:29
			minmax_result = operand_b;
		else if (info_b[3])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:225:29
			minmax_result = operand_a;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:228:7
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:229:25
					minmax_result = (operand_a_smaller ? operand_a : operand_b);
				3'b001:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:230:25
					minmax_result = (operand_a_smaller ? operand_b : operand_a);
				default:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:231:18
					minmax_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
			endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:236:3
	assign minmax_extension_bit = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:241:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] cmp_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:242:3
	reg [4:0] cmp_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:243:3
	wire cmp_extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:248:3
	always @(*) begin : comparisons
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:250:5
		cmp_result = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:251:5
		cmp_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:254:5
		if (signalling_nan)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:254:25
			cmp_status[4] = 1'b1;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:257:7
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:259:11
					if (any_operand_nan)
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:259:32
						cmp_status[4] = 1'b1;
					else
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:260:16
						cmp_result = (operand_a_smaller | operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b001:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:263:11
					if (any_operand_nan)
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:263:32
						cmp_status[4] = 1'b1;
					else
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:264:16
						cmp_result = (operand_a_smaller & ~operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b010:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:267:11
					if (any_operand_nan)
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:267:32
						cmp_result = inp_pipe_op_mod_q[NUM_INP_REGS];
					else
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:268:16
						cmp_result = operands_equal ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				default:
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:270:18
					cmp_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
			endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:275:3
	assign cmp_extension_bit = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:280:3
	wire [4:0] class_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:281:3
	wire class_extension_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:282:3
	reg [9:0] class_mask_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:285:3
	always @(*) begin : classify
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:286:5
		if (info_a[7])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:287:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000010 : 10'b0001000000);
		else if (info_a[6])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:289:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000100 : 10'b0000100000);
		else if (info_a[5])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:291:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000001000 : 10'b0000010000);
		else if (info_a[4])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:293:7
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000001 : 10'b0010000000);
		else if (info_a[3])
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:295:7
			class_mask_d = (info_a[2] ? 10'b0100000000 : 10'b1000000000);
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:297:7
			class_mask_d = 10'b1000000000;
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:301:3
	assign class_status = 1'sb0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:302:3
	assign class_extension_bit = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:307:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:308:3
	reg [4:0] status_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:309:3
	reg extension_bit_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:310:3
	wire is_class_d;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:313:3
	always @(*) begin : select_result
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:314:5
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(6): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:316:9
				result_d = sgnj_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:317:9
				status_d = sgnj_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:318:9
				extension_bit_d = sgnj_extension_bit;
			end
			sv2v_cast_A53F3(7): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:321:9
				result_d = minmax_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:322:9
				status_d = minmax_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:323:9
				extension_bit_d = minmax_extension_bit;
			end
			sv2v_cast_A53F3(8): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:326:9
				result_d = cmp_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:327:9
				status_d = cmp_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:328:9
				extension_bit_d = cmp_extension_bit;
			end
			sv2v_cast_A53F3(9): begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:331:9
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:332:9
				status_d = class_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:333:9
				extension_bit_d = class_extension_bit;
			end
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:336:9
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:337:9
				status_d = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:338:9
				extension_bit_d = fpnew_pkg_DONT_CARE;
			end
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:343:3
	assign is_class_d = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(9);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:349:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:350:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:351:3
	reg [0:NUM_OUT_REGS] out_pipe_extension_bit_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:352:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 10) + ((NUM_OUT_REGS * 10) - 1) : ((NUM_OUT_REGS + 1) * 10) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 10 : 0)] out_pipe_class_mask_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:353:3
	reg [0:NUM_OUT_REGS] out_pipe_is_class_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:354:3
	reg [(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((1 - NUM_OUT_REGS) * (TagType_TagType_TagType_TagType_TAGW + 2)) + ((NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1) : ((1 - NUM_OUT_REGS) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (((TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) - 1)) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? ((NUM_OUT_REGS + 1) * (TagType_TagType_TagType_TagType_TAGW + 2)) - 1 : ((NUM_OUT_REGS + 1) * (1 - (TagType_TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TagType_TAGW + 0))):(0 >= NUM_OUT_REGS ? ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? NUM_OUT_REGS * (TagType_TagType_TagType_TagType_TAGW + 2) : (TagType_TagType_TagType_TagType_TAGW + 1) + (NUM_OUT_REGS * (1 - (TagType_TagType_TagType_TagType_TAGW + 1)))) : ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1))] out_pipe_tag_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:355:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:356:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:358:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:361:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_07494;
	assign sv2v_tmp_07494 = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_07494;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:362:3
	wire [5:1] sv2v_tmp_CCE43;
	assign sv2v_tmp_CCE43 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_CCE43;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:363:3
	wire [1:1] sv2v_tmp_8E9A9;
	assign sv2v_tmp_8E9A9 = extension_bit_d;
	always @(*) out_pipe_extension_bit_q[0] = sv2v_tmp_8E9A9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:364:3
	wire [10:1] sv2v_tmp_94259;
	assign sv2v_tmp_94259 = class_mask_d;
	always @(*) out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 10+:10] = sv2v_tmp_94259;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:365:3
	wire [1:1] sv2v_tmp_7DF01;
	assign sv2v_tmp_7DF01 = is_class_d;
	always @(*) out_pipe_is_class_q[0] = sv2v_tmp_7DF01;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:366:3
	wire [((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)) * 1:1] sv2v_tmp_3B808;
	assign sv2v_tmp_3B808 = inp_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	always @(*) out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] = sv2v_tmp_3B808;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:367:3
	wire [1:1] sv2v_tmp_FA930;
	assign sv2v_tmp_FA930 = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_FA930;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:368:3
	wire [1:1] sv2v_tmp_2CB8C;
	assign sv2v_tmp_2CB8C = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_2CB8C;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:370:3
	assign inp_pipe_ready[NUM_INP_REGS] = out_pipe_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:372:3
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:374:5
			wire reg_ena;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:378:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:380:252
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:380:330
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:380:408
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:380:560
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:382:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:384:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:384:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:384:193
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:384:301
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:385:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:385:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:385:193
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:385:301
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:386:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:386:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:386:193
					out_pipe_extension_bit_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:386:301
					out_pipe_extension_bit_q[i + 1] <= (reg_ena ? out_pipe_extension_bit_q[i] : out_pipe_extension_bit_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:387:94
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:387:150
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:387:206
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= 10'b1000000000;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:387:314
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= (reg_ena ? out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 10+:10] : out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:388:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:388:137
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:388:193
					out_pipe_is_class_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:388:301
					out_pipe_is_class_q[i + 1] <= (reg_ena ? out_pipe_is_class_q[i] : out_pipe_is_class_q[i + 1]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:389:91
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:389:147
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:389:203
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= sv2v_cast_5B742(1'sb0);
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:389:311
					out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] <= (reg_ena ? out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))] : out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))]);
			// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:390:91
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:390:147
				if (!rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:390:203
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:390:311
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:393:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:395:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:396:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:397:3
	assign extension_bit_o = out_pipe_extension_bit_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:398:3
	assign class_mask_o = out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 10+:10];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:399:3
	assign is_class_o = out_pipe_is_class_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:400:3
	assign tag_o = out_pipe_tag_q[((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TagType_TAGW + 1) + ((0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:401:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:402:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_noncomp.sv:403:3
	assign busy_o = |{inp_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_opgroup_block_398FA_A5D02 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TagType_TAGW_type
	parameter signed [31:0] TagType_TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:15:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:17:13
	parameter [31:0] Width = 32;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:18:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:19:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtMask = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:20:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtMask = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:21:13
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	parameter [159:0] FmtPipeRegs = {fpnew_pkg_NUM_FP_FORMATS {32'd0}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:22:13
	// removed localparam type fpnew_pkg_unit_type_t
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	parameter [9:0] FmtUnitTypes = {fpnew_pkg_NUM_FP_FORMATS {2'd1}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:23:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:24:41
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:26:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:27:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:376:48
		input reg [1:0] grp;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:377:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:29:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:30:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:32:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:33:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:34:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:35:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:36:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:37:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:38:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:39:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:40:3
	input wire vectorial_op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:41:3
	input wire [TagType_TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:43:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:44:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:45:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:47:3
	output wire [Width - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:48:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:49:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:50:3
	output wire [TagType_TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:52:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:53:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:55:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:61:3
	// removed localparam type output_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:69:3
	wire [4:0] fmt_in_ready;
	wire [4:0] fmt_out_valid;
	wire [4:0] fmt_out_ready;
	wire [4:0] fmt_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:70:3
	wire [(5 * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) - 1:0] fmt_outputs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:75:3
	assign in_ready_o = in_valid_i & fmt_in_ready[dst_fmt_i];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:80:3
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic fpnew_pkg_any_enabled_multi;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:456:46
		input reg [9:0] types;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:456:70
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:457:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:457:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:457:10
				begin : sv2v_autoblock_2
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_any_enabled_multi = 1'b1;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_any_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [2:0] fpnew_pkg_get_first_enabled_multi;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:474:58
		input reg [9:0] types;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:474:82
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:475:5
			begin : sv2v_autoblock_3
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:475:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:475:10
				begin : sv2v_autoblock_4
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_get_first_enabled_multi = sv2v_cast_0BC43(i);
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_get_first_enabled_multi = sv2v_cast_0BC43(0);
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic fpnew_pkg_is_first_enabled_multi;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:464:51
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:465:51
		input reg [9:0] types;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:466:51
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:467:5
			begin : sv2v_autoblock_5
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:467:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:467:10
				begin : sv2v_autoblock_6
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:468:7
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_is_first_enabled_multi = sv2v_cast_0BC43(i) == fmt;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_is_first_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic [((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) - 1:0] sv2v_cast_4D796;
		input reg [((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) - 1:0] inp;
		sv2v_cast_4D796 = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_parallel_slices
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:82:5
			localparam [0:0] ANY_MERGED = fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:83:5
			localparam [0:0] IS_FIRST_MERGED = fpnew_pkg_is_first_enabled_multi(sv2v_cast_0BC43(fmt), FmtUnitTypes, FpFmtMask);
			if (FpFmtMask[fmt] && (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd1)) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:89:7
				wire in_valid;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:91:7
				assign in_valid = in_valid_i & (dst_fmt_i == fmt);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:93:7
				fpnew_opgroup_fmt_slice_970CB_15734 #(
					.TagType_TagType_TagType_TAGW(TagType_TagType_TAGW),
					.OpGroup(OpGroup),
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.Width(Width),
					.EnableVectors(EnableVectors),
					.NumPipeRegs(FmtPipeRegs[(4 - fmt) * 32+:32]),
					.PipeConfig(PipeConfig)
				) i_fmt_slice(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.operands_i(operands_i),
					.is_boxed_i(is_boxed_i[fmt * NUM_OPERANDS+:NUM_OPERANDS]),
					.rnd_mode_i(rnd_mode_i),
					.op_i(op_i),
					.op_mod_i(op_mod_i),
					.vectorial_op_i(vectorial_op_i),
					.tag_i(tag_i),
					.in_valid_i(in_valid),
					.in_ready_o(fmt_in_ready[fmt]),
					.flush_i(flush_i),
					.result_o(fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))-:((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) >= (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) - (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))) + 1)]),
					.status_o(fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)-:((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) >= (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) - (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) + 1)]),
					.extension_bit_o(fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)]),
					.tag_o(fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) - 1)-:((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1))]),
					.out_valid_o(fmt_out_valid[fmt]),
					.out_ready_i(fmt_out_ready[fmt]),
					.busy_o(fmt_busy[fmt])
				);
			end
			else if ((FpFmtMask[fmt] && ANY_MERGED) && !IS_FIRST_MERGED) begin : merged_unused
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:125:7
				localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:127:7
				assign fmt_in_ready[fmt] = fmt_in_ready[sv2v_cast_32_signed(FMT)];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:129:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:130:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:132:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))-:((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) >= (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) - (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))) + 1)] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:133:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)-:((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) >= (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) - (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) + 1)] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:134:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)] = fpnew_pkg_DONT_CARE;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:135:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) - 1)-:((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1))] = sv2v_cast_4D796(fpnew_pkg_DONT_CARE);
			end
			else if (!FpFmtMask[fmt] || (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd0)) begin : disable_fmt
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:139:7
				assign fmt_in_ready[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:140:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:141:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:143:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))-:((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) >= (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) - (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))) + 1)] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:144:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)-:((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) >= (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) - (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) + 1)] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:145:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)] = fpnew_pkg_DONT_CARE;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:146:7
				assign fmt_outputs[(fmt * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) - 1)-:((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1))] = sv2v_cast_4D796(fpnew_pkg_DONT_CARE);
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:153:3
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_get_num_regs_multi;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:482:54
		input reg [159:0] regs;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:483:54
		input reg [9:0] types;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:484:54
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:485:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:486:5
			begin : sv2v_autoblock_7
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:486:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:486:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:487:7
						if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2))
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:487:41
							res = fpnew_pkg_maximum(res, regs[(4 - i) * 32+:32]);
					end
			end
			fpnew_pkg_get_num_regs_multi = res;
		end
	endfunction
	generate
		if (fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask)) begin : gen_merged_slice
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:155:5
			localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:156:5
			localparam REG = fpnew_pkg_get_num_regs_multi(FmtPipeRegs, FmtUnitTypes, FpFmtMask);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:158:5
			wire in_valid;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:160:5
			assign in_valid = in_valid_i & (FmtUnitTypes[(4 - dst_fmt_i) * 2+:2] == 2'd2);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:162:5
			fpnew_opgroup_multifmt_slice_F0F3F_DD878 #(
				.TagType_TagType_TagType_TAGW(TagType_TagType_TAGW),
				.OpGroup(OpGroup),
				.Width(Width),
				.FpFmtConfig(FpFmtMask),
				.IntFmtConfig(IntFmtMask),
				.EnableVectors(EnableVectors),
				.NumPipeRegs(REG),
				.PipeConfig(PipeConfig)
			) i_multifmt_slice(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i),
				.is_boxed_i(is_boxed_i),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.in_valid_i(in_valid),
				.in_ready_o(fmt_in_ready[FMT]),
				.flush_i(flush_i),
				.result_o(fmt_outputs[(FMT * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))-:((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) >= (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) - (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))) + 1)]),
				.status_o(fmt_outputs[(FMT * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)-:((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) >= (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) - (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) + 1)]),
				.extension_bit_o(fmt_outputs[(FMT * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)]),
				.tag_o(fmt_outputs[(FMT * ((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)))) + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) - 1)-:((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1))]),
				.out_valid_o(fmt_out_valid[FMT]),
				.out_ready_i(fmt_out_ready[FMT]),
				.busy_o(fmt_busy[FMT])
			);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:201:3
	wire [((Width + 6) + ((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1))) - 1:0] arbiter_output;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:204:3
	rr_arb_tree_4FDAD_74659 #(
		.DataType_TagType_TagType_TAGW(TagType_TagType_TAGW),
		.DataType_Width(Width),
		.NumIn(NUM_FORMATS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(1'sb0),
		.req_i(fmt_out_valid),
		.gnt_o(fmt_out_ready),
		.data_i(fmt_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:223:3
	assign result_o = arbiter_output[Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)-:((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) >= (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) - (6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((6 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (Width + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5))) + 1)];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:224:3
	assign status_o = arbiter_output[((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5-:((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) >= (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) ? ((((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5) - (1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0))) + 1 : ((1 + (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0)) - (((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 5)) + 1)];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:225:3
	assign extension_bit_o = arbiter_output[((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) + 0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:226:3
	assign tag_o = arbiter_output[((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1)) - 1-:((TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:228:3
	assign busy_o = |fmt_busy;
endmodule
module fpnew_opgroup_block_E7A9E (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:15:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:17:13
	parameter [31:0] Width = 32;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:18:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:19:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtMask = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:20:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtMask = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:21:13
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	parameter [159:0] FmtPipeRegs = {fpnew_pkg_NUM_FP_FORMATS {32'd0}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:22:13
	// removed localparam type fpnew_pkg_unit_type_t
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	parameter [9:0] FmtUnitTypes = {fpnew_pkg_NUM_FP_FORMATS {2'd1}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:23:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:24:41
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:26:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:27:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:376:48
		input reg [1:0] grp;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:377:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:29:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:30:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:32:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:33:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:34:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:35:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:36:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:37:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:38:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:39:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:40:3
	input wire vectorial_op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:41:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:43:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:44:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:45:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:47:3
	output wire [Width - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:48:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:49:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:50:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:52:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:53:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:55:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:61:3
	// removed localparam type output_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:69:3
	wire [4:0] fmt_in_ready;
	wire [4:0] fmt_out_valid;
	wire [4:0] fmt_out_ready;
	wire [4:0] fmt_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:70:3
	wire [((Width + 6) >= 0 ? (5 * (Width + 7)) - 1 : (5 * (1 - (Width + 6))) + (Width + 5)):((Width + 6) >= 0 ? 0 : Width + 6)] fmt_outputs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:75:3
	assign in_ready_o = in_valid_i & fmt_in_ready[dst_fmt_i];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:80:3
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic fpnew_pkg_any_enabled_multi;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:456:46
		input reg [9:0] types;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:456:70
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:457:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:457:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:457:10
				begin : sv2v_autoblock_2
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_any_enabled_multi = 1'b1;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_any_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [2:0] fpnew_pkg_get_first_enabled_multi;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:474:58
		input reg [9:0] types;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:474:82
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:475:5
			begin : sv2v_autoblock_3
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:475:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:475:10
				begin : sv2v_autoblock_4
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_get_first_enabled_multi = sv2v_cast_0BC43(i);
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_get_first_enabled_multi = sv2v_cast_0BC43(0);
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic fpnew_pkg_is_first_enabled_multi;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:464:51
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:465:51
		input reg [9:0] types;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:466:51
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:467:5
			begin : sv2v_autoblock_5
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:467:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:467:10
				begin : sv2v_autoblock_6
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:468:7
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_is_first_enabled_multi = sv2v_cast_0BC43(i) == fmt;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_is_first_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_parallel_slices
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:82:5
			localparam [0:0] ANY_MERGED = fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:83:5
			localparam [0:0] IS_FIRST_MERGED = fpnew_pkg_is_first_enabled_multi(sv2v_cast_0BC43(fmt), FmtUnitTypes, FpFmtMask);
			if (FpFmtMask[fmt] && (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd1)) begin : active_format
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:89:7
				wire in_valid;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:91:7
				assign in_valid = in_valid_i & (dst_fmt_i == fmt);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:93:7
				fpnew_opgroup_fmt_slice_09303 #(
					.OpGroup(OpGroup),
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.Width(Width),
					.EnableVectors(EnableVectors),
					.NumPipeRegs(FmtPipeRegs[(4 - fmt) * 32+:32]),
					.PipeConfig(PipeConfig)
				) i_fmt_slice(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.operands_i(operands_i),
					.is_boxed_i(is_boxed_i[fmt * NUM_OPERANDS+:NUM_OPERANDS]),
					.rnd_mode_i(rnd_mode_i),
					.op_i(op_i),
					.op_mod_i(op_mod_i),
					.vectorial_op_i(vectorial_op_i),
					.tag_i(tag_i),
					.in_valid_i(in_valid),
					.in_ready_o(fmt_in_ready[fmt]),
					.flush_i(flush_i),
					.result_o(fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6)) : (((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6))) + ((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))) - 1)-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))]),
					.status_o(fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0) : ((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0)) + 4)-:5]),
					.extension_bit_o(fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 1 : Width + 5)]),
					.tag_o(fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 0 : Width + 6)]),
					.out_valid_o(fmt_out_valid[fmt]),
					.out_ready_i(fmt_out_ready[fmt]),
					.busy_o(fmt_busy[fmt])
				);
			end
			else if ((FpFmtMask[fmt] && ANY_MERGED) && !IS_FIRST_MERGED) begin : merged_unused
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:125:7
				localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:127:7
				assign fmt_in_ready[fmt] = fmt_in_ready[sv2v_cast_32_signed(FMT)];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:129:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:130:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:132:7
				assign fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6)) : (((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6))) + ((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))) - 1)-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:133:7
				assign fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0) : ((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0)) + 4)-:5] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:134:7
				assign fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 1 : Width + 5)] = fpnew_pkg_DONT_CARE;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:135:7
				assign fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 0 : Width + 6)] = fpnew_pkg_DONT_CARE;
			end
			else if (!FpFmtMask[fmt] || (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd0)) begin : disable_fmt
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:139:7
				assign fmt_in_ready[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:140:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:141:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:143:7
				assign fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6)) : (((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6))) + ((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))) - 1)-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:144:7
				assign fmt_outputs[((Width + 6) >= 0 ? (fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0) : ((fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0)) + 4)-:5] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:145:7
				assign fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 1 : Width + 5)] = fpnew_pkg_DONT_CARE;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:146:7
				assign fmt_outputs[(fmt * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 0 : Width + 6)] = fpnew_pkg_DONT_CARE;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:153:3
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_get_num_regs_multi;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:482:54
		input reg [159:0] regs;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:483:54
		input reg [9:0] types;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:484:54
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:485:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:486:5
			begin : sv2v_autoblock_7
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:486:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:486:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:487:7
						if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2))
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:487:41
							res = fpnew_pkg_maximum(res, regs[(4 - i) * 32+:32]);
					end
			end
			fpnew_pkg_get_num_regs_multi = res;
		end
	endfunction
	generate
		if (fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask)) begin : gen_merged_slice
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:155:5
			localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:156:5
			localparam REG = fpnew_pkg_get_num_regs_multi(FmtPipeRegs, FmtUnitTypes, FpFmtMask);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:158:5
			wire in_valid;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:160:5
			assign in_valid = in_valid_i & (FmtUnitTypes[(4 - dst_fmt_i) * 2+:2] == 2'd2);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:162:5
			fpnew_opgroup_multifmt_slice_180FF #(
				.OpGroup(OpGroup),
				.Width(Width),
				.FpFmtConfig(FpFmtMask),
				.IntFmtConfig(IntFmtMask),
				.EnableVectors(EnableVectors),
				.NumPipeRegs(REG),
				.PipeConfig(PipeConfig)
			) i_multifmt_slice(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i),
				.is_boxed_i(is_boxed_i),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.in_valid_i(in_valid),
				.in_ready_o(fmt_in_ready[FMT]),
				.flush_i(flush_i),
				.result_o(fmt_outputs[((Width + 6) >= 0 ? (FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6)) : (((FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? Width + 6 : (Width + 6) - (Width + 6))) + ((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))) - 1)-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))]),
				.status_o(fmt_outputs[((Width + 6) >= 0 ? (FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0) : ((FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 6 : Width + 0)) + 4)-:5]),
				.extension_bit_o(fmt_outputs[(FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 1 : Width + 5)]),
				.tag_o(fmt_outputs[(FMT * ((Width + 6) >= 0 ? Width + 7 : 1 - (Width + 6))) + ((Width + 6) >= 0 ? 0 : Width + 6)]),
				.out_valid_o(fmt_out_valid[FMT]),
				.out_ready_i(fmt_out_ready[FMT]),
				.busy_o(fmt_busy[FMT])
			);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:201:3
	wire [Width + 6:0] arbiter_output;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:204:3
	rr_arb_tree_3B043_A8992 #(
		.DataType_Width(Width),
		.NumIn(NUM_FORMATS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(1'sb0),
		.req_i(fmt_out_valid),
		.gnt_o(fmt_out_ready),
		.data_i(fmt_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:223:3
	assign result_o = arbiter_output[Width + 6-:((Width + 6) >= 7 ? Width + 0 : 8 - (Width + 6))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:224:3
	assign status_o = arbiter_output[6-:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:225:3
	assign extension_bit_o = arbiter_output[1];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:226:3
	assign tag_o = arbiter_output[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_block.sv:228:3
	assign busy_o = |fmt_busy;
endmodule
module fpnew_opgroup_fmt_slice_09303 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:15:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:16:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:18:13
	parameter [31:0] Width = 32;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:19:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:20:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:21:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:22:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:24:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:376:48
		input reg [1:0] grp;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:377:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:26:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:27:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:29:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:30:3
	input wire [NUM_OPERANDS - 1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:31:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:32:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:33:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:34:3
	input wire vectorial_op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:35:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:37:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:38:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:39:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:41:3
	output wire [Width - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:42:3
	// removed localparam type fpnew_pkg_status_t
	output reg [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:43:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:44:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:46:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:47:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:49:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:52:3
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:53:3
	function automatic [31:0] fpnew_pkg_num_lanes;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:387:45
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:387:65
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:387:82
		input reg vec;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:388:5
		fpnew_pkg_num_lanes = (vec ? width / fpnew_pkg_fp_width(fmt) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_num_lanes(Width, FpFormat, EnableVectors);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:56:3
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:57:3
	wire vectorial_op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:59:3
	wire [(NUM_LANES * FP_WIDTH) - 1:0] slice_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:60:3
	wire [Width - 1:0] slice_regular_result;
	wire [Width - 1:0] slice_class_result;
	wire [Width - 1:0] slice_vec_class_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:62:3
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:63:3
	wire [NUM_LANES - 1:0] lane_ext_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:64:3
	// removed localparam type fpnew_pkg_classmask_e
	wire [(NUM_LANES * 10) - 1:0] lane_class_mask;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:65:3
	wire [NUM_LANES - 1:0] lane_tags;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:66:3
	wire [NUM_LANES - 1:0] lane_vectorial;
	wire [NUM_LANES - 1:0] lane_busy;
	wire [NUM_LANES - 1:0] lane_is_class;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:68:3
	wire result_is_vector;
	wire result_is_class;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:73:3
	assign in_ready_o = lane_in_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:74:3
	assign vectorial_op = vectorial_op_i & EnableVectors;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:79:3
	genvar lane;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (lane = 0; lane < sv2v_cast_32_signed(NUM_LANES); lane = lane + 1) begin : gen_num_lanes
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:80:5
			wire [FP_WIDTH - 1:0] local_result;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:81:5
			wire local_sign;
			if ((lane == 0) || EnableVectors) begin : active_lane
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:85:7
				wire in_valid;
				wire out_valid;
				wire out_ready;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:87:7
				reg [(NUM_OPERANDS * FP_WIDTH) - 1:0] local_operands;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:88:7
				wire [FP_WIDTH - 1:0] op_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:89:7
				wire [4:0] op_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:91:7
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:93:7
				always @(*) begin : prepare_input
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:94:9
					begin : sv2v_autoblock_1
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:94:14
						reg signed [31:0] i;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:94:14
						for (i = 0; i < sv2v_cast_32_signed(NUM_OPERANDS); i = i + 1)
							begin
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:95:11
								local_operands[i * FP_WIDTH+:FP_WIDTH] = operands_i[(i * Width) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (($unsigned(lane) + 1) * FP_WIDTH) - 1 : (((($unsigned(lane) + 1) * FP_WIDTH) - 1) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:(((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)];
							end
					end
				end
				if (OpGroup == 2'd0) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:101:9
					fpnew_fma_141C6 #(
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fma(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:129:9
					assign lane_is_class[lane] = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:130:9
					assign lane_class_mask[lane * 10+:10] = 10'b0000000001;
				end
				
				else if (OpGroup == 2'd2) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:162:9
					fpnew_noncomp_1F07E #(
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_noncomp(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.class_mask_o(lane_class_mask[lane * 10+:10]),
						.is_class_o(lane_is_class[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:195:7
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:196:7
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:199:7
				assign local_result = (lane_out_valid[lane] ? op_result : {FP_WIDTH {lane_ext_bit[0]}});
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:200:7
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] ? op_status : {5 {1'sb0}});
			end
			else begin : genblk1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:204:7
				assign lane_out_valid[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:205:7
				assign lane_in_ready[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:206:7
				assign local_result = {FP_WIDTH {lane_ext_bit[0]}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:207:7
				assign lane_status[lane * 5+:5] = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:208:7
				assign lane_busy[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:209:7
				assign lane_is_class[lane] = 1'b0;
			end
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:213:5
			assign slice_result[(($unsigned(lane) + 1) * FP_WIDTH) - 1:$unsigned(lane) * FP_WIDTH] = local_result;
			if (((lane + 1) * 8) <= Width) begin : vectorial_class
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:217:7
				assign local_sign = (((lane_class_mask[lane * 10+:10] == 10'b0000000001) || (lane_class_mask[lane * 10+:10] == 10'b0000000010)) || (lane_class_mask[lane * 10+:10] == 10'b0000000100)) || (lane_class_mask[lane * 10+:10] == 10'b0000001000);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:222:7
				assign slice_vec_class_result[((lane + 1) * 8) - 1:lane * 8] = {local_sign, ~local_sign, lane_class_mask[lane * 10+:10] == 10'b1000000000, lane_class_mask[lane * 10+:10] == 10'b0100000000, (lane_class_mask[lane * 10+:10] == 10'b0000010000) || (lane_class_mask[lane * 10+:10] == 10'b0000001000), (lane_class_mask[lane * 10+:10] == 10'b0000100000) || (lane_class_mask[lane * 10+:10] == 10'b0000000100), (lane_class_mask[lane * 10+:10] == 10'b0001000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000010), (lane_class_mask[lane * 10+:10] == 10'b0010000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000001)};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:242:3
	assign result_is_vector = lane_vectorial[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:243:3
	assign result_is_class = lane_is_class[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:245:3
	assign slice_regular_result = $signed({extension_bit_o, slice_result});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:247:3
	localparam [31:0] CLASS_VEC_BITS = ((NUM_LANES * 8) > Width ? 8 * (Width / 8) : NUM_LANES * 8);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:250:3
	generate
		if (CLASS_VEC_BITS < Width) begin : pad_vectorial_class
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:251:5
			assign slice_vec_class_result[Width - 1:CLASS_VEC_BITS] = 1'sb0;
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:256:3
	assign slice_class_result = (result_is_vector ? slice_vec_class_result : lane_class_mask[0+:10]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:259:3
	assign result_o = (result_is_class ? slice_class_result : slice_regular_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:261:3
	assign extension_bit_o = lane_ext_bit[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:262:3
	assign tag_o = lane_tags[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:263:3
	assign busy_o = |lane_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:264:3
	assign out_valid_o = lane_out_valid[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:268:3
	always @(*) begin : output_processing
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:270:5
		reg [4:0] temp_status;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:271:5
		temp_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:272:5
		begin : sv2v_autoblock_2
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:272:10
			reg signed [31:0] i;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:272:10
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:273:7
					temp_status = temp_status | lane_status[i * 5+:5];
				end
		end
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:274:5
		status_o = temp_status;
	end
endmodule
module fpnew_opgroup_fmt_slice_970CB_15734 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TagType_TagType_TAGW_type
	parameter signed [31:0] TagType_TagType_TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:15:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:16:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:18:13
	parameter [31:0] Width = 32;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:19:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:20:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:21:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:22:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:24:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:376:48
		input reg [1:0] grp;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:377:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:26:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:27:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:29:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:30:3
	input wire [NUM_OPERANDS - 1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:31:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:32:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:33:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:34:3
	input wire vectorial_op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:35:3
	input wire [TagType_TagType_TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:37:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:38:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:39:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:41:3
	output wire [Width - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:42:3
	// removed localparam type fpnew_pkg_status_t
	output reg [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:43:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:44:3
	output wire [TagType_TagType_TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:46:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:47:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:49:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:52:3
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:53:3
	function automatic [31:0] fpnew_pkg_num_lanes;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:387:45
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:387:65
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:387:82
		input reg vec;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:388:5
		fpnew_pkg_num_lanes = (vec ? width / fpnew_pkg_fp_width(fmt) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_num_lanes(Width, FpFormat, EnableVectors);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:56:3
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:57:3
	wire vectorial_op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:59:3
	wire [(NUM_LANES * FP_WIDTH) - 1:0] slice_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:60:3
	wire [Width - 1:0] slice_regular_result;
	wire [Width - 1:0] slice_class_result;
	wire [Width - 1:0] slice_vec_class_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:62:3
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:63:3
	wire [NUM_LANES - 1:0] lane_ext_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:64:3
	// removed localparam type fpnew_pkg_classmask_e
	wire [(NUM_LANES * 10) - 1:0] lane_class_mask;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:65:3
	wire [((TagType_TagType_TagType_TAGW + 1) >= 0 ? (NUM_LANES * (TagType_TagType_TagType_TAGW + 2)) - 1 : (NUM_LANES * (1 - (TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TAGW + 0)):((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1)] lane_tags;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:66:3
	wire [NUM_LANES - 1:0] lane_vectorial;
	wire [NUM_LANES - 1:0] lane_busy;
	wire [NUM_LANES - 1:0] lane_is_class;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:68:3
	wire result_is_vector;
	wire result_is_class;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:73:3
	assign in_ready_o = lane_in_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:74:3
	assign vectorial_op = vectorial_op_i & EnableVectors;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:79:3
	genvar lane;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (lane = 0; lane < sv2v_cast_32_signed(NUM_LANES); lane = lane + 1) begin : gen_num_lanes
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:80:5
			wire [FP_WIDTH - 1:0] local_result;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:81:5
			wire local_sign;
			if ((lane == 0) || EnableVectors) begin : active_lane
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:85:7
				wire in_valid;
				wire out_valid;
				wire out_ready;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:87:7
				reg [(NUM_OPERANDS * FP_WIDTH) - 1:0] local_operands;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:88:7
				wire [FP_WIDTH - 1:0] op_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:89:7
				wire [4:0] op_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:91:7
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:93:7
				always @(*) begin : prepare_input
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:94:9
					begin : sv2v_autoblock_1
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:94:14
						reg signed [31:0] i;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:94:14
						for (i = 0; i < sv2v_cast_32_signed(NUM_OPERANDS); i = i + 1)
							begin
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:95:11
								local_operands[i * FP_WIDTH+:FP_WIDTH] = operands_i[(i * Width) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (($unsigned(lane) + 1) * FP_WIDTH) - 1 : (((($unsigned(lane) + 1) * FP_WIDTH) - 1) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:(((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)];
							end
					end
				end
				if (OpGroup == 2'd0) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:101:9
					fpnew_fma_1D182_0A4E9 #(
						.TagType_TagType_TagType_TagType_TAGW(TagType_TagType_TagType_TAGW),
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fma(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1) + (lane * ((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1))]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:129:9
					assign lane_is_class[lane] = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:130:9
					assign lane_class_mask[lane * 10+:10] = 10'b0000000001;
				end
				
				else if (OpGroup == 2'd2) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:162:9
					fpnew_noncomp_546BA_F0963 #(
						.TagType_TagType_TagType_TagType_TAGW(TagType_TagType_TagType_TAGW),
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_noncomp(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.class_mask_o(lane_class_mask[lane * 10+:10]),
						.is_class_o(lane_is_class[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1) + (lane * ((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1))]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:195:7
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:196:7
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:199:7
				assign local_result = (lane_out_valid[lane] ? op_result : {FP_WIDTH {lane_ext_bit[0]}});
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:200:7
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] ? op_status : {5 {1'sb0}});
			end
			else begin : genblk1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:204:7
				assign lane_out_valid[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:205:7
				assign lane_in_ready[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:206:7
				assign local_result = {FP_WIDTH {lane_ext_bit[0]}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:207:7
				assign lane_status[lane * 5+:5] = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:208:7
				assign lane_busy[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:209:7
				assign lane_is_class[lane] = 1'b0;
			end
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:213:5
			assign slice_result[(($unsigned(lane) + 1) * FP_WIDTH) - 1:$unsigned(lane) * FP_WIDTH] = local_result;
			if (((lane + 1) * 8) <= Width) begin : vectorial_class
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:217:7
				assign local_sign = (((lane_class_mask[lane * 10+:10] == 10'b0000000001) || (lane_class_mask[lane * 10+:10] == 10'b0000000010)) || (lane_class_mask[lane * 10+:10] == 10'b0000000100)) || (lane_class_mask[lane * 10+:10] == 10'b0000001000);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:222:7
				assign slice_vec_class_result[((lane + 1) * 8) - 1:lane * 8] = {local_sign, ~local_sign, lane_class_mask[lane * 10+:10] == 10'b1000000000, lane_class_mask[lane * 10+:10] == 10'b0100000000, (lane_class_mask[lane * 10+:10] == 10'b0000010000) || (lane_class_mask[lane * 10+:10] == 10'b0000001000), (lane_class_mask[lane * 10+:10] == 10'b0000100000) || (lane_class_mask[lane * 10+:10] == 10'b0000000100), (lane_class_mask[lane * 10+:10] == 10'b0001000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000010), (lane_class_mask[lane * 10+:10] == 10'b0010000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000001)};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:242:3
	assign result_is_vector = lane_vectorial[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:243:3
	assign result_is_class = lane_is_class[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:245:3
	assign slice_regular_result = $signed({extension_bit_o, slice_result});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:247:3
	localparam [31:0] CLASS_VEC_BITS = ((NUM_LANES * 8) > Width ? 8 * (Width / 8) : NUM_LANES * 8);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:250:3
	generate
		if (CLASS_VEC_BITS < Width) begin : pad_vectorial_class
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:251:5
			assign slice_vec_class_result[Width - 1:CLASS_VEC_BITS] = 1'sb0;
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:256:3
	assign slice_class_result = (result_is_vector ? slice_vec_class_result : lane_class_mask[0+:10]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:259:3
	assign result_o = (result_is_class ? slice_class_result : slice_regular_result);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:261:3
	assign extension_bit_o = lane_ext_bit[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:262:3
	assign tag_o = lane_tags[((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1) + 0+:((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:263:3
	assign busy_o = |lane_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:264:3
	assign out_valid_o = lane_out_valid[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:268:3
	always @(*) begin : output_processing
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:270:5
		reg [4:0] temp_status;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:271:5
		temp_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:272:5
		begin : sv2v_autoblock_2
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:272:10
			reg signed [31:0] i;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:272:10
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:273:7
					temp_status = temp_status | lane_status[i * 5+:5];
				end
		end
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_fmt_slice.sv:274:5
		status_o = temp_status;
	end
endmodule
module fpnew_opgroup_multifmt_slice_180FF (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:17:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:18:13
	parameter [31:0] Width = 64;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:20:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:21:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:22:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:23:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:24:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:25:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:27:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:376:48
		input reg [1:0] grp;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:377:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:28:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:30:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:31:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:33:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:34:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:35:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:36:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:37:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:38:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:39:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:40:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:41:3
	input wire vectorial_op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:42:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:44:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:45:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:46:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:48:3
	output wire [Width - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:49:3
	// removed localparam type fpnew_pkg_status_t
	output reg [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:50:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:51:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:53:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:54:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:56:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:59:3
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:306:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:307:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:310:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] MAX_FP_WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:60:3
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:86:45
		input reg [1:0] ifmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:87:5
		case (ifmt)
			sv2v_cast_87CC5(0): fpnew_pkg_int_width = 8;
			sv2v_cast_87CC5(1): fpnew_pkg_int_width = 16;
			sv2v_cast_87CC5(2): fpnew_pkg_int_width = 32;
			sv2v_cast_87CC5(3): fpnew_pkg_int_width = 64;
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:94:9
				$fatal(1, "Invalid INT format supplied");
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:98:9
				fpnew_pkg_int_width = sv2v_cast_87CC5(0);
			end
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:353:49
		input reg [0:3] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:354:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:5
			begin : sv2v_autoblock_2
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:10
				reg signed [31:0] ifmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:356:7
						if (cfg[ifmt])
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:356:22
							res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)));
					end
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:61:3
	function automatic signed [31:0] fpnew_pkg_minimum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:289:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:289:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:290:5
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:315:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:316:5
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:317:5
			begin : sv2v_autoblock_3
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:317:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:317:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:319:9
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:392:49
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:392:69
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:392:86
		input reg vec;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:393:5
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_max_num_lanes(Width, FpFmtConfig, 1'b1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:62:3
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:64:3
	localparam [31:0] FMT_BITS = fpnew_pkg_maximum(3, 2);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:66:3
	localparam [31:0] AUX_BITS = FMT_BITS + 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:68:3
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:69:3
	wire vectorial_op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:70:3
	wire [FMT_BITS - 1:0] dst_fmt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:71:3
	wire [AUX_BITS - 1:0] aux_data;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:74:3
	wire dst_fmt_is_int;
	wire dst_is_cpk;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:75:3
	wire [1:0] dst_vec_op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:76:3
	wire [2:0] target_aux_d;
	wire [2:0] target_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:77:3
	wire is_up_cast;
	wire is_down_cast;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:79:3
	wire [(NUM_FORMATS * Width) - 1:0] fmt_slice_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:80:3
	wire [(NUM_INT_FORMATS * Width) - 1:0] ifmt_slice_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:81:3
	wire [Width - 1:0] conv_slice_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:84:3
	wire [Width - 1:0] conv_target_d;
	wire [Width - 1:0] conv_target_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:86:3
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:87:3
	wire [NUM_LANES - 1:0] lane_ext_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:88:3
	wire [NUM_LANES - 1:0] lane_tags;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:89:3
	wire [(NUM_LANES * AUX_BITS) - 1:0] lane_aux;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:90:3
	wire [NUM_LANES - 1:0] lane_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:92:3
	wire result_is_vector;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:93:3
	wire [FMT_BITS - 1:0] result_fmt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:94:3
	wire result_fmt_is_int;
	wire result_is_cpk;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:95:3
	wire [1:0] result_vec_op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:100:3
	assign in_ready_o = lane_in_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:101:3
	assign vectorial_op = vectorial_op_i & EnableVectors;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:104:3
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	assign dst_fmt_is_int = (OpGroup == 2'd3) & (op_i == sv2v_cast_A53F3(11));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:105:3
	assign dst_is_cpk = (OpGroup == 2'd3) & ((op_i == sv2v_cast_A53F3(13)) || (op_i == sv2v_cast_A53F3(14)));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:107:3
	assign dst_vec_op = (OpGroup == 2'd3) & {op_i == sv2v_cast_A53F3(14), op_mod_i};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:109:3
	assign is_up_cast = fpnew_pkg_fp_width(dst_fmt_i) > fpnew_pkg_fp_width(src_fmt_i);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:110:3
	assign is_down_cast = fpnew_pkg_fp_width(dst_fmt_i) < fpnew_pkg_fp_width(src_fmt_i);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:113:3
	assign dst_fmt = (dst_fmt_is_int ? int_fmt_i : dst_fmt_i);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:116:3
	assign aux_data = {dst_fmt_is_int, vectorial_op, dst_fmt};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:117:3
	assign target_aux_d = {dst_vec_op, dst_is_cpk};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:120:3
	generate
		if (OpGroup == 2'd3) begin : conv_target
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:121:5
			assign conv_target_d = (dst_is_cpk ? operands_i[2 * Width+:Width] : operands_i[Width+:Width]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:125:3
	reg [4:0] is_boxed_1op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:126:3
	reg [9:0] is_boxed_2op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:128:3
	always @(*) begin : boxed_2op
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:129:5
		begin : sv2v_autoblock_4
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:129:10
			reg signed [31:0] fmt;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:129:10
			for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
				begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:130:7
					is_boxed_1op[fmt] = is_boxed_i[fmt * NUM_OPERANDS];
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:131:7
					is_boxed_2op[fmt * 2+:2] = is_boxed_i[(fmt * NUM_OPERANDS) + 1-:2];
				end
		end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:138:3
	genvar lane;
	localparam [0:4] fpnew_pkg_CPK_FORMATS = 5'b11000;
	function automatic [0:4] fpnew_pkg_get_conv_lane_formats;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:426:56
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:427:56
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:428:56
		input reg [31:0] lane_no;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:429:5
		reg [0:4] res;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:430:5
			begin : sv2v_autoblock_5
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:430:10
				reg [31:0] fmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:430:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:432:7
						res[fmt] = cfg[fmt] && (((width / fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))) > lane_no) || (fpnew_pkg_CPK_FORMATS[fmt] && (lane_no < 2)));
					end
			end
			fpnew_pkg_get_conv_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_conv_lane_int_formats;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:438:61
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:439:61
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:440:61
		input reg [0:3] icfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:441:61
		input reg [31:0] lane_no;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:442:5
		reg [0:3] res;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:443:5
		reg [0:4] lanefmts;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:444:5
			res = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:445:5
			lanefmts = fpnew_pkg_get_conv_lane_formats(width, cfg, lane_no);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:447:5
			begin : sv2v_autoblock_6
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:447:10
				reg [31:0] ifmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:447:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_7
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:448:12
						reg [31:0] fmt;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:448:12
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							begin
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:450:9
								res[ifmt] = res[ifmt] | ((icfg[ifmt] && lanefmts[fmt]) && (fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt)) == fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt))));
							end
					end
			end
			fpnew_pkg_get_conv_lane_int_formats = res;
		end
	endfunction
	function automatic [0:4] fpnew_pkg_get_lane_formats;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:397:51
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:398:51
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:399:51
		input reg [31:0] lane_no;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:400:5
		reg [0:4] res;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:401:5
			begin : sv2v_autoblock_8
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:401:10
				reg [31:0] fmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:401:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:403:7
						res[fmt] = cfg[fmt] & ((width / fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))) > lane_no);
					end
			end
			fpnew_pkg_get_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_lane_int_formats;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:408:56
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:409:56
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:410:56
		input reg [0:3] icfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:411:56
		input reg [31:0] lane_no;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:412:5
		reg [0:3] res;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:413:5
		reg [0:4] lanefmts;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:414:5
			res = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:415:5
			lanefmts = fpnew_pkg_get_lane_formats(width, cfg, lane_no);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:417:5
			begin : sv2v_autoblock_9
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:417:10
				reg [31:0] ifmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:417:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_10
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:418:12
						reg [31:0] fmt;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:418:12
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							if (fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt)) == fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)))
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:421:11
								res[ifmt] = res[ifmt] | (icfg[ifmt] && lanefmts[fmt]);
					end
			end
			fpnew_pkg_get_lane_int_formats = res;
		end
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [4:0] sv2v_cast_F8FCA;
		input reg [4:0] inp;
		sv2v_cast_F8FCA = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (lane = 0; lane < sv2v_cast_32_signed(NUM_LANES); lane = lane + 1) begin : gen_num_lanes
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:139:5
			localparam [31:0] LANE = $unsigned(lane);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:141:5
			localparam [0:4] ACTIVE_FORMATS = fpnew_pkg_get_lane_formats(Width, FpFmtConfig, LANE);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:143:5
			localparam [0:3] ACTIVE_INT_FORMATS = fpnew_pkg_get_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:145:5
			localparam [31:0] MAX_WIDTH = fpnew_pkg_max_fp_width(ACTIVE_FORMATS);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:148:5
			localparam [0:4] CONV_FORMATS = fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, LANE);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:150:5
			localparam [0:3] CONV_INT_FORMATS = fpnew_pkg_get_conv_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:152:5
			localparam [31:0] CONV_WIDTH = fpnew_pkg_max_fp_width(CONV_FORMATS);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:155:5
			localparam [0:4] LANE_FORMATS = (OpGroup == 2'd3 ? CONV_FORMATS : ACTIVE_FORMATS);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:157:5
			localparam [31:0] LANE_WIDTH = (OpGroup == 2'd3 ? CONV_WIDTH : MAX_WIDTH);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:159:5
			wire [LANE_WIDTH - 1:0] local_result;
			if ((lane == 0) || EnableVectors) begin : active_lane
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:163:7
				wire in_valid;
				wire out_valid;
				wire out_ready;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:165:7
				reg [(NUM_OPERANDS * LANE_WIDTH) - 1:0] local_operands;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:166:7
				wire [LANE_WIDTH - 1:0] op_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:167:7
				wire [4:0] op_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:169:7
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:172:7
				always @(*) begin : prepare_input
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:173:9
					begin : sv2v_autoblock_11
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:173:14
						reg [31:0] i;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:173:14
						for (i = 0; i < NUM_OPERANDS; i = i + 1)
							begin
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:174:11
								local_operands[i * (OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[i * Width+:Width] >> (LANE * fpnew_pkg_fp_width(src_fmt_i));
							end
					end
					if (OpGroup == 2'd3)
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:180:11
						if (op_i == sv2v_cast_A53F3(12))
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:181:13
							local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[0+:Width] >> (LANE * fpnew_pkg_int_width(int_fmt_i));
						else if (op_i == sv2v_cast_A53F3(10)) begin
							begin
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:184:13
								if ((vectorial_op && op_mod_i) && is_up_cast)
									// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:185:15
									local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[0+:Width] >> ((LANE * fpnew_pkg_fp_width(src_fmt_i)) + (MAX_FP_WIDTH / 2));
							end
						end
						else if (dst_is_cpk)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:190:13
							if (lane == 1)
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:191:15
								local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[Width + (LANE_WIDTH - 1)-:LANE_WIDTH];
				end
				if (OpGroup == 2'd0) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:199:9
					fpnew_fma_multi_7F4A8_72E9B #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_fma_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				else if (OpGroup == 2'd1) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:231:9
					fpnew_divsqrt_multi_EA2AD_2C8BD #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_divsqrt_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) * 2]),
						.is_boxed_i(is_boxed_2op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				
				else if (OpGroup == 2'd3) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:262:9
					fpnew_cast_multi_7061A_0B31A #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.IntFmtConfig(CONV_INT_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_cast_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))]),
						.is_boxed_i(is_boxed_1op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.int_fmt_i(int_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:297:7
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:298:7
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:301:7
				assign local_result = (lane_out_valid[lane] ? op_result : {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) : fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))) {lane_ext_bit[0]}});
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:302:7
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] ? op_status : {5 {1'sb0}});
			end
			else begin : inactive_lane
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:306:7
				assign lane_out_valid[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:307:7
				assign lane_in_ready[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:308:7
				assign local_result = {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) : fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))) {lane_ext_bit[0]}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:309:7
				assign lane_status[lane * 5+:5] = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:310:7
				assign lane_busy[lane] = 1'b0;
			end
			genvar fmt;
			for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1) begin : pack_fp_result
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:316:7
				localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
				if (ACTIVE_FORMATS[fmt]) begin : genblk1
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:319:9
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = local_result[FP_WIDTH - 1:0];
				end
				else if (((LANE + 1) * FP_WIDTH) <= Width) begin : genblk1
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:322:9
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = {((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1) {lane_ext_bit[LANE]}};
				end
				else if ((LANE * FP_WIDTH) < Width) begin : genblk1
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:325:9
					assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (LANE * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[LANE]}};
				end
			end
			if (OpGroup == 2'd3) begin : int_results_enabled
				genvar ifmt;
				for (ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt = ifmt + 1) begin : pack_int_result
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:334:9
					localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
					if (ACTIVE_INT_FORMATS[ifmt]) begin : genblk1
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:336:11
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = local_result[INT_WIDTH - 1:0];
					end
					else if (((LANE + 1) * INT_WIDTH) <= Width) begin : genblk1
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:339:11
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = 1'sb0;
					end
					else if ((LANE * INT_WIDTH) < Width) begin : genblk1
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:341:11
						assign ifmt_slice_result[(ifmt * Width) + ((Width - 1) >= (LANE * INT_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (LANE * INT_WIDTH) ? ((Width - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (LANE * INT_WIDTH) ? ((Width - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (Width - 1)) + 1)] = 1'sb0;
					end
				end
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:348:3
	genvar fmt;
	generate
		for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1) begin : extend_fp_result
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:350:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			if ((NUM_LANES * FP_WIDTH) < Width) begin : genblk1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:352:7
				assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[0]}};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:356:3
	genvar ifmt;
	generate
		for (ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt = ifmt + 1) begin : int_results_disabled
			if (OpGroup != 2'd3) begin : mute_int_result
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:358:7
				assign ifmt_slice_result[ifmt * Width+:Width] = 1'sb0;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:363:3
	generate
		if (OpGroup == 2'd3) begin : target_regs
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:365:5
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * Width) + ((NumPipeRegs * Width) - 1) : ((NumPipeRegs + 1) * Width) - 1):(0 >= NumPipeRegs ? NumPipeRegs * Width : 0)] byp_pipe_target_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:366:5
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * 3) + ((NumPipeRegs * 3) - 1) : ((NumPipeRegs + 1) * 3) - 1):(0 >= NumPipeRegs ? NumPipeRegs * 3 : 0)] byp_pipe_aux_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:367:5
			reg [0:NumPipeRegs] byp_pipe_valid_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:369:5
			wire [0:NumPipeRegs] byp_pipe_ready;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:372:5
			wire [Width * 1:1] sv2v_tmp_FBD8C;
			assign sv2v_tmp_FBD8C = conv_target_d;
			always @(*) byp_pipe_target_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * Width+:Width] = sv2v_tmp_FBD8C;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:373:5
			wire [3:1] sv2v_tmp_A0A5D;
			assign sv2v_tmp_A0A5D = target_aux_d;
			always @(*) byp_pipe_aux_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * 3+:3] = sv2v_tmp_A0A5D;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:374:5
			wire [1:1] sv2v_tmp_49222;
			assign sv2v_tmp_49222 = in_valid_i & vectorial_op;
			always @(*) byp_pipe_valid_q[0] = sv2v_tmp_49222;
			genvar i;
			for (i = 0; i < NumPipeRegs; i = i + 1) begin : gen_bypass_pipeline
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:378:7
				wire reg_ena;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:382:7
				assign byp_pipe_ready[i] = byp_pipe_ready[i + 1] | ~byp_pipe_valid_q[i + 1];
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:384:254
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:384:332
					if (!rst_ni)
						// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:384:410
						byp_pipe_valid_q[i + 1] <= 1'b0;
					else
						// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:384:562
						byp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (byp_pipe_ready[i] ? byp_pipe_valid_q[i] : byp_pipe_valid_q[i + 1]));
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:386:7
				assign reg_ena = byp_pipe_ready[i] & byp_pipe_valid_q[i];
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:388:71
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:388:127
					if (!rst_ni)
						// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:388:183
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= 1'sb0;
					else
						// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:388:291
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= (reg_ena ? byp_pipe_target_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * Width+:Width] : byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width]);
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:389:71
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:389:127
					if (!rst_ni)
						// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:389:183
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= 1'sb0;
					else
						// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:389:291
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= (reg_ena ? byp_pipe_aux_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * 3+:3] : byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3]);
			end
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:392:5
			assign byp_pipe_ready[NumPipeRegs] = out_ready_i & result_is_vector;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:394:5
			assign conv_target_q = byp_pipe_target_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * Width+:Width];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:397:5
			assign {result_vec_op, result_is_cpk} = byp_pipe_aux_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * 3+:3];
		end
		else begin : no_conv
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:399:5
			assign {result_vec_op, result_is_cpk} = 1'sb0;
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:405:3
	assign {result_fmt_is_int, result_is_vector, result_fmt} = lane_aux[0+:AUX_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:407:3
	assign result_o = (result_fmt_is_int ? ifmt_slice_result[result_fmt * Width+:Width] : fmt_slice_result[result_fmt * Width+:Width]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:411:3
	assign extension_bit_o = lane_ext_bit[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:412:3
	assign tag_o = lane_tags[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:413:3
	assign busy_o = |lane_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:415:3
	assign out_valid_o = lane_out_valid[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:418:3
	always @(*) begin : output_processing
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:420:5
		reg [4:0] temp_status;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:421:5
		temp_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:422:5
		begin : sv2v_autoblock_12
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:422:10
			reg signed [31:0] i;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:422:10
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:423:7
					temp_status = temp_status | lane_status[i * 5+:5];
				end
		end
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:424:5
		status_o = temp_status;
	end
endmodule
module fpnew_opgroup_multifmt_slice_F0F3F_DD878 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TagType_TagType_TAGW_type
	parameter signed [31:0] TagType_TagType_TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:17:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:18:13
	parameter [31:0] Width = 64;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:20:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:21:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtConfig = 1'sb1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:22:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:23:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:24:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:25:38
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:27:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:376:48
		input reg [1:0] grp;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:377:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:28:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:30:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:31:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:33:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:34:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:35:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:36:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:37:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:38:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:39:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:40:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:41:3
	input wire vectorial_op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:42:3
	input wire [TagType_TagType_TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:44:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:45:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:46:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:48:3
	output wire [Width - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:49:3
	// removed localparam type fpnew_pkg_status_t
	output reg [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:50:3
	output wire extension_bit_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:51:3
	output wire [TagType_TagType_TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:53:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:54:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:56:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:59:3
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:293:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:294:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:306:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:307:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:5
			begin : sv2v_autoblock_1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:308:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:310:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] MAX_FP_WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:60:3
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:86:45
		input reg [1:0] ifmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:87:5
		case (ifmt)
			sv2v_cast_87CC5(0): fpnew_pkg_int_width = 8;
			sv2v_cast_87CC5(1): fpnew_pkg_int_width = 16;
			sv2v_cast_87CC5(2): fpnew_pkg_int_width = 32;
			sv2v_cast_87CC5(3): fpnew_pkg_int_width = 64;
			default: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:94:9
				$fatal(1, "Invalid INT format supplied");
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:98:9
				fpnew_pkg_int_width = sv2v_cast_87CC5(0);
			end
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:353:49
		input reg [0:3] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:354:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:5
			begin : sv2v_autoblock_2
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:10
				reg signed [31:0] ifmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:355:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:356:7
						if (cfg[ifmt])
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:356:22
							res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)));
					end
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:61:3
	function automatic signed [31:0] fpnew_pkg_minimum;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:289:34
		input reg signed [31:0] a;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:289:41
		input reg signed [31:0] b;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:290:5
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:315:48
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:316:5
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:317:5
			begin : sv2v_autoblock_3
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:317:10
				reg [31:0] i;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:317:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:319:9
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:392:49
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:392:69
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:392:86
		input reg vec;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:393:5
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_max_num_lanes(Width, FpFmtConfig, 1'b1);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:62:3
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:64:3
	localparam [31:0] FMT_BITS = fpnew_pkg_maximum(3, 2);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:66:3
	localparam [31:0] AUX_BITS = FMT_BITS + 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:68:3
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:69:3
	wire vectorial_op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:70:3
	wire [FMT_BITS - 1:0] dst_fmt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:71:3
	wire [AUX_BITS - 1:0] aux_data;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:74:3
	wire dst_fmt_is_int;
	wire dst_is_cpk;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:75:3
	wire [1:0] dst_vec_op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:76:3
	wire [2:0] target_aux_d;
	wire [2:0] target_aux_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:77:3
	wire is_up_cast;
	wire is_down_cast;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:79:3
	wire [(NUM_FORMATS * Width) - 1:0] fmt_slice_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:80:3
	wire [(NUM_INT_FORMATS * Width) - 1:0] ifmt_slice_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:81:3
	wire [Width - 1:0] conv_slice_result;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:84:3
	wire [Width - 1:0] conv_target_d;
	wire [Width - 1:0] conv_target_q;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:86:3
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:87:3
	wire [NUM_LANES - 1:0] lane_ext_bit;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:88:3
	wire [((TagType_TagType_TagType_TAGW + 1) >= 0 ? (NUM_LANES * (TagType_TagType_TagType_TAGW + 2)) - 1 : (NUM_LANES * (1 - (TagType_TagType_TagType_TAGW + 1))) + (TagType_TagType_TagType_TAGW + 0)):((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1)] lane_tags;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:89:3
	wire [(NUM_LANES * AUX_BITS) - 1:0] lane_aux;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:90:3
	wire [NUM_LANES - 1:0] lane_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:92:3
	wire result_is_vector;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:93:3
	wire [FMT_BITS - 1:0] result_fmt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:94:3
	wire result_fmt_is_int;
	wire result_is_cpk;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:95:3
	wire [1:0] result_vec_op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:100:3
	assign in_ready_o = lane_in_ready[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:101:3
	assign vectorial_op = vectorial_op_i & EnableVectors;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:104:3
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	assign dst_fmt_is_int = (OpGroup == 2'd3) & (op_i == sv2v_cast_A53F3(11));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:105:3
	assign dst_is_cpk = (OpGroup == 2'd3) & ((op_i == sv2v_cast_A53F3(13)) || (op_i == sv2v_cast_A53F3(14)));
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:107:3
	assign dst_vec_op = (OpGroup == 2'd3) & {op_i == sv2v_cast_A53F3(14), op_mod_i};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:109:3
	assign is_up_cast = fpnew_pkg_fp_width(dst_fmt_i) > fpnew_pkg_fp_width(src_fmt_i);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:110:3
	assign is_down_cast = fpnew_pkg_fp_width(dst_fmt_i) < fpnew_pkg_fp_width(src_fmt_i);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:113:3
	assign dst_fmt = (dst_fmt_is_int ? int_fmt_i : dst_fmt_i);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:116:3
	assign aux_data = {dst_fmt_is_int, vectorial_op, dst_fmt};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:117:3
	assign target_aux_d = {dst_vec_op, dst_is_cpk};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:120:3
	generate
		if (OpGroup == 2'd3) begin : conv_target
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:121:5
			assign conv_target_d = (dst_is_cpk ? operands_i[2 * Width+:Width] : operands_i[Width+:Width]);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:125:3
	reg [4:0] is_boxed_1op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:126:3
	reg [9:0] is_boxed_2op;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:128:3
	always @(*) begin : boxed_2op
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:129:5
		begin : sv2v_autoblock_4
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:129:10
			reg signed [31:0] fmt;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:129:10
			for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
				begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:130:7
					is_boxed_1op[fmt] = is_boxed_i[fmt * NUM_OPERANDS];
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:131:7
					is_boxed_2op[fmt * 2+:2] = is_boxed_i[(fmt * NUM_OPERANDS) + 1-:2];
				end
		end
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:138:3
	genvar lane;
	localparam [0:4] fpnew_pkg_CPK_FORMATS = 5'b11000;
	function automatic [0:4] fpnew_pkg_get_conv_lane_formats;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:426:56
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:427:56
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:428:56
		input reg [31:0] lane_no;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:429:5
		reg [0:4] res;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:430:5
			begin : sv2v_autoblock_5
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:430:10
				reg [31:0] fmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:430:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:432:7
						res[fmt] = cfg[fmt] && (((width / fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))) > lane_no) || (fpnew_pkg_CPK_FORMATS[fmt] && (lane_no < 2)));
					end
			end
			fpnew_pkg_get_conv_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_conv_lane_int_formats;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:438:61
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:439:61
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:440:61
		input reg [0:3] icfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:441:61
		input reg [31:0] lane_no;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:442:5
		reg [0:3] res;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:443:5
		reg [0:4] lanefmts;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:444:5
			res = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:445:5
			lanefmts = fpnew_pkg_get_conv_lane_formats(width, cfg, lane_no);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:447:5
			begin : sv2v_autoblock_6
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:447:10
				reg [31:0] ifmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:447:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_7
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:448:12
						reg [31:0] fmt;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:448:12
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							begin
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:450:9
								res[ifmt] = res[ifmt] | ((icfg[ifmt] && lanefmts[fmt]) && (fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt)) == fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt))));
							end
					end
			end
			fpnew_pkg_get_conv_lane_int_formats = res;
		end
	endfunction
	function automatic [0:4] fpnew_pkg_get_lane_formats;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:397:51
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:398:51
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:399:51
		input reg [31:0] lane_no;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:400:5
		reg [0:4] res;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:401:5
			begin : sv2v_autoblock_8
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:401:10
				reg [31:0] fmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:401:10
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:403:7
						res[fmt] = cfg[fmt] & ((width / fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))) > lane_no);
					end
			end
			fpnew_pkg_get_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_lane_int_formats;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:408:56
		input reg [31:0] width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:409:56
		input reg [0:4] cfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:410:56
		input reg [0:3] icfg;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:411:56
		input reg [31:0] lane_no;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:412:5
		reg [0:3] res;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:413:5
		reg [0:4] lanefmts;
		begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:414:5
			res = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:415:5
			lanefmts = fpnew_pkg_get_lane_formats(width, cfg, lane_no);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:417:5
			begin : sv2v_autoblock_9
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:417:10
				reg [31:0] ifmt;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:417:10
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_10
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:418:12
						reg [31:0] fmt;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:418:12
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							if (fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt)) == fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)))
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:421:11
								res[ifmt] = res[ifmt] | (icfg[ifmt] && lanefmts[fmt]);
					end
			end
			fpnew_pkg_get_lane_int_formats = res;
		end
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [4:0] sv2v_cast_F8FCA;
		input reg [4:0] inp;
		sv2v_cast_F8FCA = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (lane = 0; lane < sv2v_cast_32_signed(NUM_LANES); lane = lane + 1) begin : gen_num_lanes
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:139:5
			localparam [31:0] LANE = $unsigned(lane);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:141:5
			localparam [0:4] ACTIVE_FORMATS = fpnew_pkg_get_lane_formats(Width, FpFmtConfig, LANE);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:143:5
			localparam [0:3] ACTIVE_INT_FORMATS = fpnew_pkg_get_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:145:5
			localparam [31:0] MAX_WIDTH = fpnew_pkg_max_fp_width(ACTIVE_FORMATS);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:148:5
			localparam [0:4] CONV_FORMATS = fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, LANE);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:150:5
			localparam [0:3] CONV_INT_FORMATS = fpnew_pkg_get_conv_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:152:5
			localparam [31:0] CONV_WIDTH = fpnew_pkg_max_fp_width(CONV_FORMATS);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:155:5
			localparam [0:4] LANE_FORMATS = (OpGroup == 2'd3 ? CONV_FORMATS : ACTIVE_FORMATS);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:157:5
			localparam [31:0] LANE_WIDTH = (OpGroup == 2'd3 ? CONV_WIDTH : MAX_WIDTH);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:159:5
			wire [LANE_WIDTH - 1:0] local_result;
			if ((lane == 0) || EnableVectors) begin : active_lane
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:163:7
				wire in_valid;
				wire out_valid;
				wire out_ready;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:165:7
				reg [(NUM_OPERANDS * LANE_WIDTH) - 1:0] local_operands;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:166:7
				wire [LANE_WIDTH - 1:0] op_result;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:167:7
				wire [4:0] op_status;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:169:7
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:172:7
				always @(*) begin : prepare_input
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:173:9
					begin : sv2v_autoblock_11
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:173:14
						reg [31:0] i;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:173:14
						for (i = 0; i < NUM_OPERANDS; i = i + 1)
							begin
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:174:11
								local_operands[i * (OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[i * Width+:Width] >> (LANE * fpnew_pkg_fp_width(src_fmt_i));
							end
					end
					if (OpGroup == 2'd3)
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:180:11
						if (op_i == sv2v_cast_A53F3(12))
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:181:13
							local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[0+:Width] >> (LANE * fpnew_pkg_int_width(int_fmt_i));
						else if (op_i == sv2v_cast_A53F3(10)) begin
							begin
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:184:13
								if ((vectorial_op && op_mod_i) && is_up_cast)
									// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:185:15
									local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[0+:Width] >> ((LANE * fpnew_pkg_fp_width(src_fmt_i)) + (MAX_FP_WIDTH / 2));
							end
						end
						else if (dst_is_cpk)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:190:13
							if (lane == 1)
								// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:191:15
								local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[Width + (LANE_WIDTH - 1)-:LANE_WIDTH];
				end
				if (OpGroup == 2'd0) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:199:9
					fpnew_fma_multi_53FD4_8108B #(
						.AuxType_AUX_BITS(AUX_BITS),
						.TagType_TagType_TagType_TagType_TAGW(TagType_TagType_TagType_TAGW),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_fma_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1) + (lane * ((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1))]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				else if (OpGroup == 2'd1) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:231:9
					fpnew_divsqrt_multi_CBA5B_DFE5F #(
						.AuxType_AUX_BITS(AUX_BITS),
						.TagType_TagType_TagType_TagType_TAGW(TagType_TagType_TagType_TAGW),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_divsqrt_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) * 2]),
						.is_boxed_i(is_boxed_2op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1) + (lane * ((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1))]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				
				else if (OpGroup == 2'd3) begin : lane_instance
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:262:9
					fpnew_cast_multi_35196_62023 #(
						.AuxType_AUX_BITS(AUX_BITS),
						.TagType_TagType_TagType_TagType_TAGW(TagType_TagType_TagType_TAGW),
						.FpFmtConfig(LANE_FORMATS),
						.IntFmtConfig(CONV_INT_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_cast_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))]),
						.is_boxed_i(is_boxed_1op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.int_fmt_i(int_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1) + (lane * ((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1)))+:((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1))]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:297:7
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:298:7
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:301:7
				assign local_result = (lane_out_valid[lane] ? op_result : {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) : fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))) {lane_ext_bit[0]}});
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:302:7
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] ? op_status : {5 {1'sb0}});
			end
			else begin : inactive_lane
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:306:7
				assign lane_out_valid[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:307:7
				assign lane_in_ready[lane] = 1'b0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:308:7
				assign local_result = {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) : fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))) {lane_ext_bit[0]}};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:309:7
				assign lane_status[lane * 5+:5] = 1'sb0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:310:7
				assign lane_busy[lane] = 1'b0;
			end
			genvar fmt;
			for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1) begin : pack_fp_result
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:316:7
				localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
				if (ACTIVE_FORMATS[fmt]) begin : genblk1
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:319:9
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = local_result[FP_WIDTH - 1:0];
				end
				else if (((LANE + 1) * FP_WIDTH) <= Width) begin : genblk1
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:322:9
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = {((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1) {lane_ext_bit[LANE]}};
				end
				else if ((LANE * FP_WIDTH) < Width) begin : genblk1
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:325:9
					assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (LANE * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (LANE * FP_WIDTH) ? ((Width - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[LANE]}};
				end
			end
			if (OpGroup == 2'd3) begin : int_results_enabled
				genvar ifmt;
				for (ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt = ifmt + 1) begin : pack_int_result
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:334:9
					localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
					if (ACTIVE_INT_FORMATS[ifmt]) begin : genblk1
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:336:11
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = local_result[INT_WIDTH - 1:0];
					end
					else if (((LANE + 1) * INT_WIDTH) <= Width) begin : genblk1
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:339:11
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = 1'sb0;
					end
					else if ((LANE * INT_WIDTH) < Width) begin : genblk1
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:341:11
						assign ifmt_slice_result[(ifmt * Width) + ((Width - 1) >= (LANE * INT_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (LANE * INT_WIDTH) ? ((Width - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (LANE * INT_WIDTH) ? ((Width - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (Width - 1)) + 1)] = 1'sb0;
					end
				end
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:348:3
	genvar fmt;
	generate
		for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1) begin : extend_fp_result
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:350:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			if ((NUM_LANES * FP_WIDTH) < Width) begin : genblk1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:352:7
				assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[0]}};
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:356:3
	genvar ifmt;
	generate
		for (ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt = ifmt + 1) begin : int_results_disabled
			if (OpGroup != 2'd3) begin : mute_int_result
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:358:7
				assign ifmt_slice_result[ifmt * Width+:Width] = 1'sb0;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:363:3
	generate
		if (OpGroup == 2'd3) begin : target_regs
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:365:5
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * Width) + ((NumPipeRegs * Width) - 1) : ((NumPipeRegs + 1) * Width) - 1):(0 >= NumPipeRegs ? NumPipeRegs * Width : 0)] byp_pipe_target_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:366:5
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * 3) + ((NumPipeRegs * 3) - 1) : ((NumPipeRegs + 1) * 3) - 1):(0 >= NumPipeRegs ? NumPipeRegs * 3 : 0)] byp_pipe_aux_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:367:5
			reg [0:NumPipeRegs] byp_pipe_valid_q;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:369:5
			wire [0:NumPipeRegs] byp_pipe_ready;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:372:5
			wire [Width * 1:1] sv2v_tmp_FBD8C;
			assign sv2v_tmp_FBD8C = conv_target_d;
			always @(*) byp_pipe_target_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * Width+:Width] = sv2v_tmp_FBD8C;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:373:5
			wire [3:1] sv2v_tmp_A0A5D;
			assign sv2v_tmp_A0A5D = target_aux_d;
			always @(*) byp_pipe_aux_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * 3+:3] = sv2v_tmp_A0A5D;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:374:5
			wire [1:1] sv2v_tmp_49222;
			assign sv2v_tmp_49222 = in_valid_i & vectorial_op;
			always @(*) byp_pipe_valid_q[0] = sv2v_tmp_49222;
			genvar i;
			for (i = 0; i < NumPipeRegs; i = i + 1) begin : gen_bypass_pipeline
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:378:7
				wire reg_ena;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:382:7
				assign byp_pipe_ready[i] = byp_pipe_ready[i + 1] | ~byp_pipe_valid_q[i + 1];
				// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:384:254
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:384:332
					if (!rst_ni)
						// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:384:410
						byp_pipe_valid_q[i + 1] <= 1'b0;
					else
						// Trace: macro expansion of FFLARNC at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:384:562
						byp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (byp_pipe_ready[i] ? byp_pipe_valid_q[i] : byp_pipe_valid_q[i + 1]));
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:386:7
				assign reg_ena = byp_pipe_ready[i] & byp_pipe_valid_q[i];
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:388:71
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:388:127
					if (!rst_ni)
						// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:388:183
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= 1'sb0;
					else
						// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:388:291
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= (reg_ena ? byp_pipe_target_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * Width+:Width] : byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width]);
				// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:389:71
				always @(posedge clk_i or negedge rst_ni)
					// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:389:127
					if (!rst_ni)
						// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:389:183
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= 1'sb0;
					else
						// Trace: macro expansion of FFL at ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:389:291
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= (reg_ena ? byp_pipe_aux_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * 3+:3] : byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3]);
			end
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:392:5
			assign byp_pipe_ready[NumPipeRegs] = out_ready_i & result_is_vector;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:394:5
			assign conv_target_q = byp_pipe_target_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * Width+:Width];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:397:5
			assign {result_vec_op, result_is_cpk} = byp_pipe_aux_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * 3+:3];
		end
		else begin : no_conv
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:399:5
			assign {result_vec_op, result_is_cpk} = 1'sb0;
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:405:3
	assign {result_fmt_is_int, result_is_vector, result_fmt} = lane_aux[0+:AUX_BITS];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:407:3
	assign result_o = (result_fmt_is_int ? ifmt_slice_result[result_fmt * Width+:Width] : fmt_slice_result[result_fmt * Width+:Width]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:411:3
	assign extension_bit_o = lane_ext_bit[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:412:3
	assign tag_o = lane_tags[((TagType_TagType_TagType_TAGW + 1) >= 0 ? 0 : TagType_TagType_TagType_TAGW + 1) + 0+:((TagType_TagType_TagType_TAGW + 1) >= 0 ? TagType_TagType_TagType_TAGW + 2 : 1 - (TagType_TagType_TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:413:3
	assign busy_o = |lane_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:415:3
	assign out_valid_o = lane_out_valid[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:418:3
	always @(*) begin : output_processing
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:420:5
		reg [4:0] temp_status;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:421:5
		temp_status = 1'sb0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:422:5
		begin : sv2v_autoblock_12
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:422:10
			reg signed [31:0] i;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:422:10
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:423:7
					temp_status = temp_status | lane_status[i * 5+:5];
				end
		end
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_opgroup_multifmt_slice.sv:424:5
		status_o = temp_status;
	end
endmodule
// removed package "fpnew_pkg"
module fpnew_rounding (
	abs_value_i,
	sign_i,
	round_sticky_bits_i,
	rnd_mode_i,
	effective_subtraction_i,
	abs_rounded_o,
	sign_o,
	exact_zero_o
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:15:13
	parameter [31:0] AbsWidth = 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:18:3
	input wire [AbsWidth - 1:0] abs_value_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:19:3
	input wire sign_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:21:3
	input wire [1:0] round_sticky_bits_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:22:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:23:3
	input wire effective_subtraction_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:25:3
	output wire [AbsWidth - 1:0] abs_rounded_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:26:3
	output wire sign_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:28:3
	output wire exact_zero_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:31:3
	reg round_up;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:42:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	always @(*) begin : rounding_decision
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:43:5
		case (rnd_mode_i)
			3'b000:
				case (round_sticky_bits_i)
					2'b00, 2'b01:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:47:18
						round_up = 1'b0;
					2'b10:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:48:18
						round_up = abs_value_i[0];
					2'b11:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:49:18
						round_up = 1'b1;
					default:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:50:20
						round_up = fpnew_pkg_DONT_CARE;
				endcase
			3'b001:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:52:23
				round_up = 1'b0;
			3'b010:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:53:23
				round_up = (|round_sticky_bits_i ? sign_i : 1'b0);
			3'b011:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:54:23
				round_up = (|round_sticky_bits_i ? ~sign_i : 1'b0);
			3'b100:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:55:23
				round_up = round_sticky_bits_i[1];
			default:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:56:16
				round_up = fpnew_pkg_DONT_CARE;
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:61:3
	assign abs_rounded_o = abs_value_i + round_up;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:64:3
	assign exact_zero_o = (abs_value_i == {AbsWidth {1'sb0}}) && (round_sticky_bits_i == {2 {1'sb0}});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_rounding.sv:68:3
	assign sign_o = (exact_zero_o && effective_subtraction_i ? rnd_mode_i == 3'b010 : sign_i);
endmodule
module fpnew_top_3ED0B_1EC5F (
	clk_i,
	rst_ni,
	operands_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TAGW_type
	parameter signed [31:0] TagType_TAGW = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:16:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	// removed localparam type fpnew_pkg_fpu_features_t
	localparam [42:0] fpnew_pkg_RV64D_Xsflt = 43'h000000207ff;
	parameter [42:0] Features = fpnew_pkg_RV64D_Xsflt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:17:13
	// removed localparam type fpnew_pkg_pipe_config_t
	// removed localparam type fpnew_pkg_unit_type_t
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unit_types_t
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unsigned_t
	// removed localparam type fpnew_pkg_fpu_implementation_t
	function automatic [159:0] sv2v_cast_B9240;
		input reg [159:0] inp;
		sv2v_cast_B9240 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_CDC93;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_CDC93 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_15FEF;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_15FEF = inp;
	endfunction
	localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] fpnew_pkg_DEFAULT_NOREGS = {sv2v_cast_CDC93({fpnew_pkg_NUM_OPGROUPS {sv2v_cast_B9240(0)}}), sv2v_cast_15FEF({{fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}, {fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}}), 2'd0};
	parameter [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] Implementation = fpnew_pkg_DEFAULT_NOREGS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:18:45
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:20:14
	localparam [31:0] WIDTH = Features[42-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:21:14
	localparam [31:0] NUM_OPERANDS = 3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:23:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:24:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:26:3
	input wire [(NUM_OPERANDS * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:27:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:28:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:29:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:30:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:31:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:32:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:33:3
	input wire vectorial_op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:34:3
	input wire [TagType_TAGW + 1:0] tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:36:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:37:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:38:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:40:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:41:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:42:3
	output wire [TagType_TAGW + 1:0] tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:44:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:45:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:47:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:50:3
	localparam [31:0] NUM_OPGROUPS = fpnew_pkg_NUM_OPGROUPS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:51:3
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:56:3
	// removed localparam type output_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:63:3
	wire [3:0] opgrp_in_ready;
	wire [3:0] opgrp_out_valid;
	wire [3:0] opgrp_out_ready;
	wire [3:0] opgrp_ext;
	wire [3:0] opgrp_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:64:3
	wire [(4 * ((WIDTH + 5) + (TagType_TAGW + 2))) - 1:0] opgrp_outputs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:66:3
	wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:71:3
	// removed localparam type fpnew_pkg_opgroup_e
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [1:0] fpnew_pkg_get_opgroup;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:365:44
		input reg [3:0] op;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:366:5
		case (op)
			sv2v_cast_A53F3(0), sv2v_cast_A53F3(1), sv2v_cast_A53F3(2), sv2v_cast_A53F3(3): fpnew_pkg_get_opgroup = 2'd0;
			sv2v_cast_A53F3(4), sv2v_cast_A53F3(5): fpnew_pkg_get_opgroup = 2'd1;
			sv2v_cast_A53F3(6), sv2v_cast_A53F3(7), sv2v_cast_A53F3(8), sv2v_cast_A53F3(9): fpnew_pkg_get_opgroup = 2'd2;
			sv2v_cast_A53F3(10), sv2v_cast_A53F3(11), sv2v_cast_A53F3(12), sv2v_cast_A53F3(13), sv2v_cast_A53F3(14): fpnew_pkg_get_opgroup = 2'd3;
			default: fpnew_pkg_get_opgroup = 2'd2;
		endcase
	endfunction
	assign in_ready_o = in_valid_i & opgrp_in_ready[fpnew_pkg_get_opgroup(op_i)];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:74:3
	genvar fmt;
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_nanbox_check
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:75:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			if (Features[9] && (FP_WIDTH < WIDTH)) begin : check
				genvar op;
				for (op = 0; op < sv2v_cast_32_signed(NUM_OPERANDS); op = op + 1) begin : operands
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:79:9
					assign is_boxed[(fmt * NUM_OPERANDS) + op] = (!vectorial_op_i ? operands_i[(op * WIDTH) + ((WIDTH - 1) >= FP_WIDTH ? WIDTH - 1 : ((WIDTH - 1) + ((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)) - 1)-:((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)] == {((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1) * 1 {1'sb1}} : 1'b1);
				end
			end
			else begin : no_check
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:84:7
				assign is_boxed[fmt * NUM_OPERANDS+:NUM_OPERANDS] = 1'sb1;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:91:3
	genvar opgrp;
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:376:48
		input reg [1:0] grp;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:377:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		for (opgrp = 0; opgrp < sv2v_cast_32_signed(NUM_OPGROUPS); opgrp = opgrp + 1) begin : gen_operation_groups
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:92:5
			localparam [31:0] NUM_OPS = fpnew_pkg_num_operands(sv2v_cast_2(opgrp));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:94:5
			wire in_valid;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:95:5
			reg [(NUM_FORMATS * NUM_OPS) - 1:0] input_boxed;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:97:5
			assign in_valid = in_valid_i & (fpnew_pkg_get_opgroup(op_i) == sv2v_cast_2(opgrp));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:100:5
			always @(*) begin : slice_inputs
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:101:7
				begin : sv2v_autoblock_1
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:101:12
					reg [31:0] fmt;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:101:12
					for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
						begin
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:102:9
							input_boxed[fmt * fpnew_pkg_num_operands(sv2v_cast_2(opgrp))+:fpnew_pkg_num_operands(sv2v_cast_2(opgrp))] = is_boxed[(fmt * NUM_OPERANDS) + (NUM_OPS - 1)-:NUM_OPS];
						end
				end
			end
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:105:5
			fpnew_opgroup_block_398FA_A5D02 #(
				.TagType_TagType_TAGW(TagType_TAGW),
				.OpGroup(sv2v_cast_2(opgrp)),
				.Width(WIDTH),
				.EnableVectors(Features[10]),
				.FpFmtMask(Features[8-:5]),
				.IntFmtMask(Features[3-:fpnew_pkg_NUM_INT_FORMATS]),
				.FmtPipeRegs(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + (((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1)) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) - 1) - (32 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:160]),
				.FmtUnitTypes(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) - 1) - (2 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:10]),
				.PipeConfig(Implementation[1-:2])
			) i_opgroup_block(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i[WIDTH * ((NUM_OPS - 1) - (NUM_OPS - 1))+:WIDTH * NUM_OPS]),
				.is_boxed_i(input_boxed),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.in_valid_i(in_valid),
				.in_ready_o(opgrp_in_ready[opgrp]),
				.flush_i(flush_i),
				.result_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + (TagType_TAGW + 2))) + (WIDTH + (5 + (TagType_TAGW + 1)))-:((WIDTH + (5 + (TagType_TAGW + 1))) >= (5 + (TagType_TAGW + 2)) ? ((WIDTH + (5 + (TagType_TAGW + 1))) - (5 + (TagType_TAGW + 2))) + 1 : ((5 + (TagType_TAGW + 2)) - (WIDTH + (5 + (TagType_TAGW + 1)))) + 1)]),
				.status_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + (TagType_TAGW + 2))) + (5 + (TagType_TAGW + 1))-:((5 + (TagType_TAGW + 1)) >= (TagType_TAGW + 2) ? ((5 + (TagType_TAGW + 1)) - (TagType_TAGW + 2)) + 1 : ((TagType_TAGW + 2) - (5 + (TagType_TAGW + 1))) + 1)]),
				.extension_bit_o(opgrp_ext[opgrp]),
				.tag_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + (TagType_TAGW + 2))) + (TagType_TAGW + 1)-:((TagType_TAGW + 1) >= 0 ? TagType_TAGW + 2 : 1 - (TagType_TAGW + 1))]),
				.out_valid_o(opgrp_out_valid[opgrp]),
				.out_ready_i(opgrp_out_ready[opgrp]),
				.busy_o(opgrp_busy[opgrp])
			);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:144:3
	wire [((WIDTH + 5) + (TagType_TAGW + 2)) - 1:0] arbiter_output;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:147:3
	rr_arb_tree_12F9A_F22A2 #(
		.DataType_TagType_TAGW(TagType_TAGW),
		.DataType_WIDTH(WIDTH),
		.NumIn(NUM_OPGROUPS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(1'sb0),
		.req_i(opgrp_out_valid),
		.gnt_o(opgrp_out_ready),
		.data_i(opgrp_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:166:3
	assign result_o = arbiter_output[WIDTH + (5 + (TagType_TAGW + 1))-:((WIDTH + (5 + (TagType_TAGW + 1))) >= (5 + (TagType_TAGW + 2)) ? ((WIDTH + (5 + (TagType_TAGW + 1))) - (5 + (TagType_TAGW + 2))) + 1 : ((5 + (TagType_TAGW + 2)) - (WIDTH + (5 + (TagType_TAGW + 1)))) + 1)];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:167:3
	assign status_o = arbiter_output[5 + (TagType_TAGW + 1)-:((5 + (TagType_TAGW + 1)) >= (TagType_TAGW + 2) ? ((5 + (TagType_TAGW + 1)) - (TagType_TAGW + 2)) + 1 : ((TagType_TAGW + 2) - (5 + (TagType_TAGW + 1))) + 1)];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:168:3
	assign tag_o = arbiter_output[TagType_TAGW + 1-:((TagType_TAGW + 1) >= 0 ? TagType_TAGW + 2 : 1 - (TagType_TAGW + 1))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:170:3
	assign busy_o = |opgrp_busy;
endmodule
module fpnew_top_FF541 (
	clk_i,
	rst_ni,
	operands_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:16:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	// removed localparam type fpnew_pkg_fpu_features_t
	localparam [42:0] fpnew_pkg_RV64D_Xsflt = 43'h000000207ff;
	parameter [42:0] Features = fpnew_pkg_RV64D_Xsflt;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:17:13
	// removed localparam type fpnew_pkg_pipe_config_t
	// removed localparam type fpnew_pkg_unit_type_t
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unit_types_t
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unsigned_t
	// removed localparam type fpnew_pkg_fpu_implementation_t
	function automatic [159:0] sv2v_cast_B9240;
		input reg [159:0] inp;
		sv2v_cast_B9240 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_CDC93;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_CDC93 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_15FEF;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_15FEF = inp;
	endfunction
	localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] fpnew_pkg_DEFAULT_NOREGS = {sv2v_cast_CDC93({fpnew_pkg_NUM_OPGROUPS {sv2v_cast_B9240(0)}}), sv2v_cast_15FEF({{fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}, {fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}}), 2'd0};
	parameter [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] Implementation = fpnew_pkg_DEFAULT_NOREGS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:18:45
	// removed localparam type TagType
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:20:14
	localparam [31:0] WIDTH = Features[42-:32];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:21:14
	localparam [31:0] NUM_OPERANDS = 3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:23:3
	input wire clk_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:24:3
	input wire rst_ni;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:26:3
	input wire [(NUM_OPERANDS * WIDTH) - 1:0] operands_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:27:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:28:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:29:3
	input wire op_mod_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:30:3
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	input wire [2:0] src_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:31:3
	input wire [2:0] dst_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:32:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:33:3
	input wire vectorial_op_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:34:3
	input wire tag_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:36:3
	input wire in_valid_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:37:3
	output wire in_ready_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:38:3
	input wire flush_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:40:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:41:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:42:3
	output wire tag_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:44:3
	output wire out_valid_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:45:3
	input wire out_ready_i;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:47:3
	output wire busy_o;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:50:3
	localparam [31:0] NUM_OPGROUPS = fpnew_pkg_NUM_OPGROUPS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:51:3
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:56:3
	// removed localparam type output_t
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:63:3
	wire [3:0] opgrp_in_ready;
	wire [3:0] opgrp_out_valid;
	wire [3:0] opgrp_out_ready;
	wire [3:0] opgrp_ext;
	wire [3:0] opgrp_busy;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:64:3
	wire [((WIDTH + 5) >= 0 ? (4 * (WIDTH + 6)) - 1 : (4 * (1 - (WIDTH + 5))) + (WIDTH + 4)):((WIDTH + 5) >= 0 ? 0 : WIDTH + 5)] opgrp_outputs;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:66:3
	wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:71:3
	// removed localparam type fpnew_pkg_opgroup_e
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [1:0] fpnew_pkg_get_opgroup;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:365:44
		input reg [3:0] op;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:366:5
		case (op)
			sv2v_cast_A53F3(0), sv2v_cast_A53F3(1), sv2v_cast_A53F3(2), sv2v_cast_A53F3(3): fpnew_pkg_get_opgroup = 2'd0;
			sv2v_cast_A53F3(4), sv2v_cast_A53F3(5): fpnew_pkg_get_opgroup = 2'd1;
			sv2v_cast_A53F3(6), sv2v_cast_A53F3(7), sv2v_cast_A53F3(8), sv2v_cast_A53F3(9): fpnew_pkg_get_opgroup = 2'd2;
			sv2v_cast_A53F3(10), sv2v_cast_A53F3(11), sv2v_cast_A53F3(12), sv2v_cast_A53F3(13), sv2v_cast_A53F3(14): fpnew_pkg_get_opgroup = 2'd3;
			default: fpnew_pkg_get_opgroup = 2'd2;
		endcase
	endfunction
	assign in_ready_o = in_valid_i & opgrp_in_ready[fpnew_pkg_get_opgroup(op_i)];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:74:3
	genvar fmt;
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:301:44
		input reg [2:0] fmt;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:302:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_nanbox_check
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:75:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			if (Features[9] && (FP_WIDTH < WIDTH)) begin : check
				genvar op;
				for (op = 0; op < sv2v_cast_32_signed(NUM_OPERANDS); op = op + 1) begin : operands
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:79:9
					assign is_boxed[(fmt * NUM_OPERANDS) + op] = (!vectorial_op_i ? operands_i[(op * WIDTH) + ((WIDTH - 1) >= FP_WIDTH ? WIDTH - 1 : ((WIDTH - 1) + ((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)) - 1)-:((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)] == {((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1) * 1 {1'sb1}} : 1'b1);
				end
			end
			else begin : no_check
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:84:7
				assign is_boxed[fmt * NUM_OPERANDS+:NUM_OPERANDS] = 1'sb1;
			end
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:91:3
	genvar opgrp;
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:376:48
		input reg [1:0] grp;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_pkg.sv:377:5
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		for (opgrp = 0; opgrp < sv2v_cast_32_signed(NUM_OPGROUPS); opgrp = opgrp + 1) begin : gen_operation_groups
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:92:5
			localparam [31:0] NUM_OPS = fpnew_pkg_num_operands(sv2v_cast_2(opgrp));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:94:5
			wire in_valid;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:95:5
			reg [(NUM_FORMATS * NUM_OPS) - 1:0] input_boxed;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:97:5
			assign in_valid = in_valid_i & (fpnew_pkg_get_opgroup(op_i) == sv2v_cast_2(opgrp));
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:100:5
			always @(*) begin : slice_inputs
				// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:101:7
				begin : sv2v_autoblock_1
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:101:12
					reg [31:0] fmt;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:101:12
					for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
						begin
							// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:102:9
							input_boxed[fmt * fpnew_pkg_num_operands(sv2v_cast_2(opgrp))+:fpnew_pkg_num_operands(sv2v_cast_2(opgrp))] = is_boxed[(fmt * NUM_OPERANDS) + (NUM_OPS - 1)-:NUM_OPS];
						end
				end
			end
			// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:105:5
			fpnew_opgroup_block_E7A9E #(
				.OpGroup(sv2v_cast_2(opgrp)),
				.Width(WIDTH),
				.EnableVectors(Features[10]),
				.FpFmtMask(Features[8-:5]),
				.IntFmtMask(Features[3-:fpnew_pkg_NUM_INT_FORMATS]),
				.FmtPipeRegs(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + (((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1)) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) - 1) - (32 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:160]),
				.FmtUnitTypes(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) - 1) - (2 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:10]),
				.PipeConfig(Implementation[1-:2])
			) i_opgroup_block(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i[WIDTH * ((NUM_OPS - 1) - (NUM_OPS - 1))+:WIDTH * NUM_OPS]),
				.is_boxed_i(input_boxed),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.in_valid_i(in_valid),
				.in_ready_o(opgrp_in_ready[opgrp]),
				.flush_i(flush_i),
				.result_o(opgrp_outputs[((WIDTH + 5) >= 0 ? (opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? WIDTH + 5 : (WIDTH + 5) - (WIDTH + 5)) : (((opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? WIDTH + 5 : (WIDTH + 5) - (WIDTH + 5))) + ((WIDTH + 5) >= 6 ? WIDTH + 0 : 7 - (WIDTH + 5))) - 1)-:((WIDTH + 5) >= 6 ? WIDTH + 0 : 7 - (WIDTH + 5))]),
				.status_o(opgrp_outputs[((WIDTH + 5) >= 0 ? (opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? 5 : WIDTH + 0) : ((opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? 5 : WIDTH + 0)) + 4)-:5]),
				.extension_bit_o(opgrp_ext[opgrp]),
				.tag_o(opgrp_outputs[(opgrp * ((WIDTH + 5) >= 0 ? WIDTH + 6 : 1 - (WIDTH + 5))) + ((WIDTH + 5) >= 0 ? 0 : WIDTH + 5)]),
				.out_valid_o(opgrp_out_valid[opgrp]),
				.out_ready_i(opgrp_out_ready[opgrp]),
				.busy_o(opgrp_busy[opgrp])
			);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:144:3
	wire [WIDTH + 5:0] arbiter_output;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:147:3
	rr_arb_tree_02E82_EBE23 #(
		.DataType_WIDTH(WIDTH),
		.NumIn(NUM_OPGROUPS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(1'sb0),
		.req_i(opgrp_out_valid),
		.gnt_o(opgrp_out_ready),
		.data_i(opgrp_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:166:3
	assign result_o = arbiter_output[WIDTH + 5-:((WIDTH + 5) >= 6 ? WIDTH + 0 : 7 - (WIDTH + 5))];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:167:3
	assign status_o = arbiter_output[5-:5];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:168:3
	assign tag_o = arbiter_output[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpnew_top.sv:170:3
	assign busy_o = |opgrp_busy;
endmodule
// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:41:1
// removed ["import defs_div_sqrt_mvp::*;"]
module control_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Start_SI,
	Kill_SI,
	Special_case_SBI,
	Special_case_dly_SBI,
	Precision_ctl_SI,
	Format_sel_SI,
	Numerator_DI,
	Exp_num_DI,
	Denominator_DI,
	Exp_den_DI,
	Div_start_dly_SO,
	Sqrt_start_dly_SO,
	Div_enable_SO,
	Sqrt_enable_SO,
	Full_precision_SO,
	FP32_SO,
	FP64_SO,
	FP16_SO,
	FP16ALT_SO,
	Ready_SO,
	Done_SO,
	Mant_result_prenorm_DO,
	Exp_result_prenorm_DO
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:46:4
	input wire Clk_CI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:47:4
	input wire Rst_RBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:48:4
	input wire Div_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:49:4
	input wire Sqrt_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:50:4
	input wire Start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:51:4
	input wire Kill_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:52:4
	input wire Special_case_SBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:53:4
	input wire Special_case_dly_SBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:54:4
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:55:4
	input wire [1:0] Format_sel_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:56:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Numerator_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:57:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_num_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:58:4
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Denominator_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:59:4
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_den_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:62:4
	output wire Div_start_dly_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:63:4
	output wire Sqrt_start_dly_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:64:4
	output reg Div_enable_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:65:4
	output reg Sqrt_enable_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:69:4
	output wire Full_precision_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:70:4
	output wire FP32_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:71:4
	output wire FP64_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:72:4
	output wire FP16_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:73:4
	output wire FP16ALT_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:75:4
	output reg Ready_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:76:4
	output reg Done_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:78:4
	output reg [56:0] Mant_result_prenorm_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:80:4
	output wire [12:0] Exp_result_prenorm_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:83:4
	reg [57:0] Partial_remainder_DN;
	reg [57:0] Partial_remainder_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:84:4
	reg [56:0] Quotient_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:88:4
	wire [53:0] Numerator_se_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:89:4
	wire [53:0] Denominator_se_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:90:4
	reg [53:0] Denominator_se_DB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:92:4
	assign Numerator_se_D = {1'b0, Numerator_DI};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:94:4
	assign Denominator_se_D = {1'b0, Denominator_DI};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:96:3
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:98:6
		if (FP32_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:100:10
			Denominator_se_DB = {~Denominator_se_D[53:29], {29 {1'b0}}};
		else if (FP64_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:103:10
			Denominator_se_DB = ~Denominator_se_D;
		else if (FP16_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:106:10
			Denominator_se_DB = {~Denominator_se_D[53:42], {42 {1'b0}}};
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:109:10
			Denominator_se_DB = {~Denominator_se_D[53:45], {45 {1'b0}}};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:114:4
	wire [53:0] Mant_D_sqrt_Norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:116:4
	assign Mant_D_sqrt_Norm = (Exp_num_DI[0] ? {1'b0, Numerator_DI} : {Numerator_DI, 1'b0});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:121:4
	reg [1:0] Format_sel_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:123:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:125:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:127:13
			Format_sel_S <= 'b0;
		else if (Start_SI && Ready_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:131:13
			Format_sel_S <= Format_sel_SI;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:135:13
			Format_sel_S <= Format_sel_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:139:4
	assign FP32_SO = Format_sel_S == 2'b00;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:140:4
	assign FP64_SO = Format_sel_S == 2'b01;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:141:4
	assign FP16_SO = Format_sel_S == 2'b10;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:142:4
	assign FP16ALT_SO = Format_sel_S == 2'b11;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:150:4
	reg [5:0] Precision_ctl_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:151:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:153:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:155:13
			Precision_ctl_S <= 'b0;
		else if (Start_SI && Ready_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:159:13
			Precision_ctl_S <= Precision_ctl_SI;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:163:13
			Precision_ctl_S <= Precision_ctl_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:166:3
	assign Full_precision_SO = Precision_ctl_S == 6'h00;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:170:6
	reg [5:0] State_ctl_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:171:6
	wire [5:0] State_Two_iteration_unit_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:172:6
	wire [5:0] State_Four_iteration_unit_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:174:5
	assign State_Two_iteration_unit_S = Precision_ctl_S[5:1];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:175:5
	assign State_Four_iteration_unit_S = Precision_ctl_S[5:2];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:176:6
	localparam defs_div_sqrt_mvp_Iteration_unit_num_S = 2'b10;
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:178:10
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:182:16
				case (Format_sel_S)
					2'b00:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:185:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:187:26
							State_ctl_S = 6'h1b;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:191:26
							State_ctl_S = Precision_ctl_S;
					2'b01:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:196:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:198:26
							State_ctl_S = 6'h38;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:202:26
							State_ctl_S = Precision_ctl_S;
					2'b10:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:207:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:209:26
							State_ctl_S = 6'h0e;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:213:26
							State_ctl_S = Precision_ctl_S;
					2'b11:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:218:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:220:26
							State_ctl_S = 6'h0b;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:224:26
							State_ctl_S = Precision_ctl_S;
				endcase
			2'b01:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:234:16
				case (Format_sel_S)
					2'b00:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:237:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:239:26
							State_ctl_S = 6'h0d;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:243:26
							State_ctl_S = State_Two_iteration_unit_S;
					2'b01:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:248:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:250:26
							State_ctl_S = 6'h1b;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:254:26
							State_ctl_S = State_Two_iteration_unit_S;
					2'b10:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:259:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:261:26
							State_ctl_S = 6'h06;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:265:26
							State_ctl_S = State_Two_iteration_unit_S;
					2'b11:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:270:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:272:26
							State_ctl_S = 6'h05;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:276:26
							State_ctl_S = State_Two_iteration_unit_S;
				endcase
			2'b10:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:286:16
				case (Format_sel_S)
					2'b00:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:289:22
						case (Precision_ctl_S)
							6'h00:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:292:28
								State_ctl_S = 6'h08;
							6'h06, 6'h07, 6'h08:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:296:28
								State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:300:28
								State_ctl_S = 6'h03;
							6'h0c, 6'h0d, 6'h0e:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:304:28
								State_ctl_S = 6'h04;
							6'h0f, 6'h10, 6'h11:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:308:28
								State_ctl_S = 6'h05;
							6'h12, 6'h13, 6'h14:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:312:28
								State_ctl_S = 6'h06;
							6'h15, 6'h16, 6'h17:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:316:28
								State_ctl_S = 6'h07;
							default:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:320:28
								State_ctl_S = 6'h08;
						endcase
					2'b01:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:326:22
						case (Precision_ctl_S)
							6'h00:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:329:28
								State_ctl_S = 6'h12;
							6'h06, 6'h07, 6'h08:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:333:28
								State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:337:28
								State_ctl_S = 6'h03;
							6'h0c, 6'h0d, 6'h0e:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:341:28
								State_ctl_S = 6'h04;
							6'h0f, 6'h10, 6'h11:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:345:28
								State_ctl_S = 6'h05;
							6'h12, 6'h13, 6'h14:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:349:28
								State_ctl_S = 6'h06;
							6'h15, 6'h16, 6'h17:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:353:28
								State_ctl_S = 6'h07;
							6'h18, 6'h19, 6'h1a:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:357:28
								State_ctl_S = 6'h08;
							6'h1b, 6'h1c, 6'h1d:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:361:28
								State_ctl_S = 6'h09;
							6'h1e, 6'h1f, 6'h20:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:365:28
								State_ctl_S = 6'h0a;
							6'h21, 6'h22, 6'h23:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:369:28
								State_ctl_S = 6'h0b;
							6'h24, 6'h25, 6'h26:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:373:28
								State_ctl_S = 6'h0c;
							6'h27, 6'h28, 6'h29:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:377:28
								State_ctl_S = 6'h0d;
							6'h2a, 6'h2b, 6'h2c:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:381:28
								State_ctl_S = 6'h0e;
							6'h2d, 6'h2e, 6'h2f:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:385:28
								State_ctl_S = 6'h0f;
							6'h30, 6'h31, 6'h32:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:389:28
								State_ctl_S = 6'h10;
							6'h33, 6'h34, 6'h35:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:393:28
								State_ctl_S = 6'h11;
							default:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:397:28
								State_ctl_S = 6'h12;
						endcase
					2'b10:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:403:22
						case (Precision_ctl_S)
							6'h00:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:406:28
								State_ctl_S = 6'h04;
							6'h06, 6'h07, 6'h08:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:410:28
								State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:414:28
								State_ctl_S = 6'h03;
							default:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:418:28
								State_ctl_S = 6'h04;
						endcase
					2'b11:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:424:22
						case (Precision_ctl_S)
							6'h00:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:427:28
								State_ctl_S = 6'h03;
							6'h06, 6'h07, 6'h08:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:431:28
								State_ctl_S = 6'h02;
							default:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:435:28
								State_ctl_S = 6'h03;
						endcase
				endcase
			2'b11:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:446:16
				case (Format_sel_S)
					2'b00:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:449:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:451:26
							State_ctl_S = 6'h06;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:455:26
							State_ctl_S = State_Four_iteration_unit_S;
					2'b01:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:460:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:462:26
							State_ctl_S = 6'h0d;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:466:26
							State_ctl_S = State_Four_iteration_unit_S;
					2'b10:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:471:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:473:26
							State_ctl_S = 6'h03;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:477:26
							State_ctl_S = State_Four_iteration_unit_S;
					2'b11:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:482:22
						if (Full_precision_SO)
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:484:26
							State_ctl_S = 6'h02;
						else
							// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:488:26
							State_ctl_S = State_Four_iteration_unit_S;
				endcase
		endcase
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:503:4
	reg Div_start_dly_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:505:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:507:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:509:13
			Div_start_dly_S <= 1'b0;
		else if (Div_start_SI && Ready_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:513:12
			Div_start_dly_S <= 1'b1;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:517:13
			Div_start_dly_S <= 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:521:4
	assign Div_start_dly_SO = Div_start_dly_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:523:3
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:524:5
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:525:7
			Div_enable_SO <= 1'b0;
		else if (Kill_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:528:7
			Div_enable_SO <= 1'b0;
		else if (Div_start_SI && Ready_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:530:7
			Div_enable_SO <= 1'b1;
		else if (Done_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:532:7
			Div_enable_SO <= 1'b0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:534:7
			Div_enable_SO <= Div_enable_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:537:4
	reg Sqrt_start_dly_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:539:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:541:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:543:13
			Sqrt_start_dly_S <= 1'b0;
		else if (Sqrt_start_SI && Ready_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:547:12
			Sqrt_start_dly_S <= 1'b1;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:551:13
			Sqrt_start_dly_S <= 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:554:5
	assign Sqrt_start_dly_SO = Sqrt_start_dly_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:556:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:557:5
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:558:7
			Sqrt_enable_SO <= 1'b0;
		else if (Kill_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:560:7
			Sqrt_enable_SO <= 1'b0;
		else if (Sqrt_start_SI && Ready_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:562:7
			Sqrt_enable_SO <= 1'b1;
		else if (Done_SO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:564:7
			Sqrt_enable_SO <= 1'b0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:566:7
			Sqrt_enable_SO <= Sqrt_enable_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:569:4
	reg [5:0] Crtl_cnt_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:570:4
	wire Start_dly_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:572:4
	assign Start_dly_S = Div_start_dly_S | Sqrt_start_dly_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:574:4
	wire Fsm_enable_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:575:4
	assign Fsm_enable_S = ((Start_dly_S | |Crtl_cnt_S) && ~Kill_SI) && Special_case_dly_SBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:577:4
	wire Final_state_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:578:4
	assign Final_state_S = Crtl_cnt_S == State_ctl_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:581:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:583:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:585:14
			Crtl_cnt_S <= 1'sb0;
		else if (Final_state_S | Kill_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:589:15
			Crtl_cnt_S <= 1'sb0;
		else if (Fsm_enable_S)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:593:15
			Crtl_cnt_S <= Crtl_cnt_S + 1;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:597:15
			Crtl_cnt_S <= 1'sb0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:603:5
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:605:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:607:13
			Done_SO <= 1'b0;
		else if (Start_SI && Ready_SO) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:611:13
				if (~Special_case_SBI)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:613:17
					Done_SO <= 1'b1;
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:617:17
					Done_SO <= 1'b0;
			end
		end
		else if (Final_state_S)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:622:13
			Done_SO <= 1'b1;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:626:13
			Done_SO <= 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:633:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:635:8
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:637:12
			Ready_SO <= 1'b1;
		else if (Start_SI && Ready_SO) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:642:13
				if (~Special_case_SBI)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:644:17
					Ready_SO <= 1'b1;
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:648:17
					Ready_SO <= 1'b0;
			end
		end
		else if (Final_state_S | Kill_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:653:12
			Ready_SO <= 1'b1;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:657:12
			Ready_SO <= Ready_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:666:3
	wire Qcnt_one_0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:667:3
	wire Qcnt_one_1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:668:3
	wire [1:0] Qcnt_one_2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:669:3
	wire [2:0] Qcnt_one_3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:670:3
	wire [3:0] Qcnt_one_4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:671:3
	wire [4:0] Qcnt_one_5;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:672:3
	wire [5:0] Qcnt_one_6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:673:3
	wire [6:0] Qcnt_one_7;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:674:3
	wire [7:0] Qcnt_one_8;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:675:3
	wire [8:0] Qcnt_one_9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:676:3
	wire [9:0] Qcnt_one_10;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:677:3
	wire [10:0] Qcnt_one_11;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:678:3
	wire [11:0] Qcnt_one_12;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:679:3
	wire [12:0] Qcnt_one_13;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:680:3
	wire [13:0] Qcnt_one_14;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:681:3
	wire [14:0] Qcnt_one_15;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:682:3
	wire [15:0] Qcnt_one_16;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:683:3
	wire [16:0] Qcnt_one_17;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:684:3
	wire [17:0] Qcnt_one_18;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:685:3
	wire [18:0] Qcnt_one_19;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:686:3
	wire [19:0] Qcnt_one_20;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:687:3
	wire [20:0] Qcnt_one_21;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:688:3
	wire [21:0] Qcnt_one_22;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:689:3
	wire [22:0] Qcnt_one_23;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:690:3
	wire [23:0] Qcnt_one_24;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:691:3
	wire [24:0] Qcnt_one_25;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:692:3
	wire [25:0] Qcnt_one_26;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:693:3
	wire [26:0] Qcnt_one_27;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:694:3
	wire [27:0] Qcnt_one_28;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:695:3
	wire [28:0] Qcnt_one_29;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:696:3
	wire [29:0] Qcnt_one_30;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:697:3
	wire [30:0] Qcnt_one_31;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:698:3
	wire [31:0] Qcnt_one_32;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:699:3
	wire [32:0] Qcnt_one_33;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:700:3
	wire [33:0] Qcnt_one_34;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:701:3
	wire [34:0] Qcnt_one_35;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:702:3
	wire [35:0] Qcnt_one_36;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:703:3
	wire [36:0] Qcnt_one_37;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:704:3
	wire [37:0] Qcnt_one_38;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:705:3
	wire [38:0] Qcnt_one_39;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:706:3
	wire [39:0] Qcnt_one_40;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:707:3
	wire [40:0] Qcnt_one_41;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:708:3
	wire [41:0] Qcnt_one_42;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:709:3
	wire [42:0] Qcnt_one_43;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:710:3
	wire [43:0] Qcnt_one_44;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:711:3
	wire [44:0] Qcnt_one_45;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:712:3
	wire [45:0] Qcnt_one_46;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:713:3
	wire [46:0] Qcnt_one_47;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:714:3
	wire [47:0] Qcnt_one_48;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:715:3
	wire [48:0] Qcnt_one_49;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:716:3
	wire [49:0] Qcnt_one_50;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:717:3
	wire [50:0] Qcnt_one_51;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:718:3
	wire [51:0] Qcnt_one_52;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:719:3
	wire [52:0] Qcnt_one_53;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:720:3
	wire [53:0] Qcnt_one_54;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:721:3
	wire [54:0] Qcnt_one_55;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:722:3
	wire [55:0] Qcnt_one_56;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:723:3
	wire [56:0] Qcnt_one_57;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:724:3
	wire [57:0] Qcnt_one_58;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:725:3
	wire [58:0] Qcnt_one_59;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:726:3
	wire [59:0] Qcnt_one_60;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:737:3
	wire [1:0] Qcnt_two_0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:738:3
	wire [2:0] Qcnt_two_1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:739:3
	wire [4:0] Qcnt_two_2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:740:3
	wire [6:0] Qcnt_two_3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:741:3
	wire [8:0] Qcnt_two_4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:742:3
	wire [10:0] Qcnt_two_5;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:743:3
	wire [12:0] Qcnt_two_6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:744:3
	wire [14:0] Qcnt_two_7;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:745:3
	wire [16:0] Qcnt_two_8;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:746:3
	wire [18:0] Qcnt_two_9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:747:3
	wire [20:0] Qcnt_two_10;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:748:3
	wire [22:0] Qcnt_two_11;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:749:3
	wire [24:0] Qcnt_two_12;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:750:3
	wire [26:0] Qcnt_two_13;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:751:3
	wire [28:0] Qcnt_two_14;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:752:3
	wire [30:0] Qcnt_two_15;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:753:3
	wire [32:0] Qcnt_two_16;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:754:3
	wire [34:0] Qcnt_two_17;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:755:3
	wire [36:0] Qcnt_two_18;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:756:3
	wire [38:0] Qcnt_two_19;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:757:3
	wire [40:0] Qcnt_two_20;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:758:3
	wire [42:0] Qcnt_two_21;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:759:3
	wire [44:0] Qcnt_two_22;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:760:3
	wire [46:0] Qcnt_two_23;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:761:3
	wire [48:0] Qcnt_two_24;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:762:3
	wire [50:0] Qcnt_two_25;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:763:3
	wire [52:0] Qcnt_two_26;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:764:3
	wire [54:0] Qcnt_two_27;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:765:3
	wire [56:0] Qcnt_two_28;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:774:3
	wire [2:0] Qcnt_three_0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:775:3
	wire [4:0] Qcnt_three_1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:776:3
	wire [7:0] Qcnt_three_2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:777:3
	wire [10:0] Qcnt_three_3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:778:3
	wire [13:0] Qcnt_three_4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:779:3
	wire [16:0] Qcnt_three_5;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:780:3
	wire [19:0] Qcnt_three_6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:781:3
	wire [22:0] Qcnt_three_7;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:782:3
	wire [25:0] Qcnt_three_8;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:783:3
	wire [28:0] Qcnt_three_9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:784:3
	wire [31:0] Qcnt_three_10;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:785:3
	wire [34:0] Qcnt_three_11;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:786:3
	wire [37:0] Qcnt_three_12;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:787:3
	wire [40:0] Qcnt_three_13;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:788:3
	wire [43:0] Qcnt_three_14;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:789:3
	wire [46:0] Qcnt_three_15;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:790:3
	wire [49:0] Qcnt_three_16;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:791:3
	wire [52:0] Qcnt_three_17;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:792:3
	wire [55:0] Qcnt_three_18;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:793:3
	wire [58:0] Qcnt_three_19;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:794:3
	wire [61:0] Qcnt_three_20;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:803:3
	wire [3:0] Qcnt_four_0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:804:3
	wire [6:0] Qcnt_four_1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:805:3
	wire [10:0] Qcnt_four_2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:806:3
	wire [14:0] Qcnt_four_3;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:807:3
	wire [18:0] Qcnt_four_4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:808:3
	wire [22:0] Qcnt_four_5;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:809:3
	wire [26:0] Qcnt_four_6;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:810:3
	wire [30:0] Qcnt_four_7;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:811:3
	wire [34:0] Qcnt_four_8;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:812:3
	wire [38:0] Qcnt_four_9;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:813:3
	wire [42:0] Qcnt_four_10;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:814:3
	wire [46:0] Qcnt_four_11;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:815:3
	wire [50:0] Qcnt_four_12;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:816:3
	wire [54:0] Qcnt_four_13;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:817:3
	wire [58:0] Qcnt_four_14;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:825:4
	wire [57:0] Sqrt_R0;
	reg [57:0] Sqrt_Q0;
	reg [57:0] Q_sqrt0;
	reg [57:0] Q_sqrt_com_0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:826:4
	wire [57:0] Sqrt_R1;
	reg [57:0] Sqrt_Q1;
	reg [57:0] Q_sqrt1;
	reg [57:0] Q_sqrt_com_1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:827:4
	wire [57:0] Sqrt_R2;
	reg [57:0] Sqrt_Q2;
	reg [57:0] Q_sqrt2;
	reg [57:0] Q_sqrt_com_2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:828:4
	wire [57:0] Sqrt_R3;
	reg [57:0] Sqrt_Q3;
	reg [57:0] Q_sqrt3;
	reg [57:0] Q_sqrt_com_3;
	wire [57:0] Sqrt_R4;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:831:4
	reg [1:0] Sqrt_DI [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:832:4
	wire [1:0] Sqrt_DO [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:833:4
	wire Sqrt_carry_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:836:3
	wire [57:0] Iteration_cell_a_D [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:837:3
	wire [57:0] Iteration_cell_b_D [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:838:3
	wire [57:0] Iteration_cell_a_BMASK_D [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:839:3
	wire [57:0] Iteration_cell_b_BMASK_D [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:840:3
	wire Iteration_cell_carry_D [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:841:3
	wire [57:0] Iteration_cell_sum_D [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:842:3
	wire [57:0] Iteration_cell_sum_AMASK_D [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:845:3
	reg [3:0] Sqrt_quotinent_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:848:4
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:850:7
		case (Format_sel_S)
			2'b00: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:853:13
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][28], ~Iteration_cell_sum_AMASK_D[1][28], ~Iteration_cell_sum_AMASK_D[2][28], ~Iteration_cell_sum_AMASK_D[3][28]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:854:13
				Q_sqrt_com_0 = {{29 {1'b0}}, ~Q_sqrt0[28:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:855:13
				Q_sqrt_com_1 = {{29 {1'b0}}, ~Q_sqrt1[28:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:856:13
				Q_sqrt_com_2 = {{29 {1'b0}}, ~Q_sqrt2[28:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:857:13
				Q_sqrt_com_3 = {{29 {1'b0}}, ~Q_sqrt3[28:0]};
			end
			2'b01: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:861:13
				Sqrt_quotinent_S = {Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2], Iteration_cell_carry_D[3]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:862:13
				Q_sqrt_com_0 = ~Q_sqrt0;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:863:13
				Q_sqrt_com_1 = ~Q_sqrt1;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:864:13
				Q_sqrt_com_2 = ~Q_sqrt2;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:865:13
				Q_sqrt_com_3 = ~Q_sqrt3;
			end
			2'b10: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:869:13
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][15], ~Iteration_cell_sum_AMASK_D[1][15], ~Iteration_cell_sum_AMASK_D[2][15], ~Iteration_cell_sum_AMASK_D[3][15]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:870:13
				Q_sqrt_com_0 = {{42 {1'b0}}, ~Q_sqrt0[15:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:871:13
				Q_sqrt_com_1 = {{42 {1'b0}}, ~Q_sqrt1[15:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:872:13
				Q_sqrt_com_2 = {{42 {1'b0}}, ~Q_sqrt2[15:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:873:13
				Q_sqrt_com_3 = {{42 {1'b0}}, ~Q_sqrt3[15:0]};
			end
			2'b11: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:877:13
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][12], ~Iteration_cell_sum_AMASK_D[1][12], ~Iteration_cell_sum_AMASK_D[2][12], ~Iteration_cell_sum_AMASK_D[3][12]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:878:13
				Q_sqrt_com_0 = {{45 {1'b0}}, ~Q_sqrt0[12:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:879:13
				Q_sqrt_com_1 = {{45 {1'b0}}, ~Q_sqrt1[12:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:880:13
				Q_sqrt_com_2 = {{45 {1'b0}}, ~Q_sqrt2[12:0]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:881:13
				Q_sqrt_com_3 = {{45 {1'b0}}, ~Q_sqrt3[12:0]};
			end
		endcase
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:888:3
	assign Qcnt_one_0 = 1'b0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:889:3
	assign Qcnt_one_1 = {Quotient_DP[0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:890:3
	assign Qcnt_one_2 = {Quotient_DP[1:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:891:3
	assign Qcnt_one_3 = {Quotient_DP[2:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:892:3
	assign Qcnt_one_4 = {Quotient_DP[3:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:893:3
	assign Qcnt_one_5 = {Quotient_DP[4:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:894:3
	assign Qcnt_one_6 = {Quotient_DP[5:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:895:3
	assign Qcnt_one_7 = {Quotient_DP[6:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:896:3
	assign Qcnt_one_8 = {Quotient_DP[7:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:897:3
	assign Qcnt_one_9 = {Quotient_DP[8:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:898:3
	assign Qcnt_one_10 = {Quotient_DP[9:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:899:3
	assign Qcnt_one_11 = {Quotient_DP[10:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:900:3
	assign Qcnt_one_12 = {Quotient_DP[11:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:901:3
	assign Qcnt_one_13 = {Quotient_DP[12:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:902:3
	assign Qcnt_one_14 = {Quotient_DP[13:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:903:3
	assign Qcnt_one_15 = {Quotient_DP[14:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:904:3
	assign Qcnt_one_16 = {Quotient_DP[15:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:905:3
	assign Qcnt_one_17 = {Quotient_DP[16:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:906:3
	assign Qcnt_one_18 = {Quotient_DP[17:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:907:3
	assign Qcnt_one_19 = {Quotient_DP[18:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:908:3
	assign Qcnt_one_20 = {Quotient_DP[19:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:909:3
	assign Qcnt_one_21 = {Quotient_DP[20:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:910:3
	assign Qcnt_one_22 = {Quotient_DP[21:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:911:3
	assign Qcnt_one_23 = {Quotient_DP[22:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:912:3
	assign Qcnt_one_24 = {Quotient_DP[23:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:913:3
	assign Qcnt_one_25 = {Quotient_DP[24:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:914:3
	assign Qcnt_one_26 = {Quotient_DP[25:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:915:3
	assign Qcnt_one_27 = {Quotient_DP[26:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:916:3
	assign Qcnt_one_28 = {Quotient_DP[27:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:917:3
	assign Qcnt_one_29 = {Quotient_DP[28:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:918:3
	assign Qcnt_one_30 = {Quotient_DP[29:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:919:3
	assign Qcnt_one_31 = {Quotient_DP[30:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:920:3
	assign Qcnt_one_32 = {Quotient_DP[31:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:921:3
	assign Qcnt_one_33 = {Quotient_DP[32:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:922:3
	assign Qcnt_one_34 = {Quotient_DP[33:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:923:3
	assign Qcnt_one_35 = {Quotient_DP[34:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:924:3
	assign Qcnt_one_36 = {Quotient_DP[35:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:925:3
	assign Qcnt_one_37 = {Quotient_DP[36:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:926:3
	assign Qcnt_one_38 = {Quotient_DP[37:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:927:3
	assign Qcnt_one_39 = {Quotient_DP[38:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:928:3
	assign Qcnt_one_40 = {Quotient_DP[39:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:929:3
	assign Qcnt_one_41 = {Quotient_DP[40:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:930:3
	assign Qcnt_one_42 = {Quotient_DP[41:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:931:3
	assign Qcnt_one_43 = {Quotient_DP[42:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:932:3
	assign Qcnt_one_44 = {Quotient_DP[43:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:933:3
	assign Qcnt_one_45 = {Quotient_DP[44:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:934:3
	assign Qcnt_one_46 = {Quotient_DP[45:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:935:3
	assign Qcnt_one_47 = {Quotient_DP[46:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:936:3
	assign Qcnt_one_48 = {Quotient_DP[47:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:937:3
	assign Qcnt_one_49 = {Quotient_DP[48:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:938:3
	assign Qcnt_one_50 = {Quotient_DP[49:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:939:3
	assign Qcnt_one_51 = {Quotient_DP[50:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:940:3
	assign Qcnt_one_52 = {Quotient_DP[51:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:941:3
	assign Qcnt_one_53 = {Quotient_DP[52:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:942:3
	assign Qcnt_one_54 = {Quotient_DP[53:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:943:3
	assign Qcnt_one_55 = {Quotient_DP[54:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:944:3
	assign Qcnt_one_56 = {Quotient_DP[55:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:945:3
	assign Qcnt_one_57 = {Quotient_DP[56:0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:948:3
	assign Qcnt_two_0 = {1'b0, Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:949:3
	assign Qcnt_two_1 = {Quotient_DP[1:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:950:3
	assign Qcnt_two_2 = {Quotient_DP[3:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:951:3
	assign Qcnt_two_3 = {Quotient_DP[5:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:952:3
	assign Qcnt_two_4 = {Quotient_DP[7:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:953:3
	assign Qcnt_two_5 = {Quotient_DP[9:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:954:3
	assign Qcnt_two_6 = {Quotient_DP[11:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:955:3
	assign Qcnt_two_7 = {Quotient_DP[13:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:956:3
	assign Qcnt_two_8 = {Quotient_DP[15:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:957:3
	assign Qcnt_two_9 = {Quotient_DP[17:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:958:3
	assign Qcnt_two_10 = {Quotient_DP[19:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:959:3
	assign Qcnt_two_11 = {Quotient_DP[21:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:960:3
	assign Qcnt_two_12 = {Quotient_DP[23:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:961:3
	assign Qcnt_two_13 = {Quotient_DP[25:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:962:3
	assign Qcnt_two_14 = {Quotient_DP[27:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:963:3
	assign Qcnt_two_15 = {Quotient_DP[29:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:964:3
	assign Qcnt_two_16 = {Quotient_DP[31:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:965:3
	assign Qcnt_two_17 = {Quotient_DP[33:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:966:3
	assign Qcnt_two_18 = {Quotient_DP[35:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:967:3
	assign Qcnt_two_19 = {Quotient_DP[37:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:968:3
	assign Qcnt_two_20 = {Quotient_DP[39:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:969:3
	assign Qcnt_two_21 = {Quotient_DP[41:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:970:3
	assign Qcnt_two_22 = {Quotient_DP[43:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:971:3
	assign Qcnt_two_23 = {Quotient_DP[45:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:972:3
	assign Qcnt_two_24 = {Quotient_DP[47:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:973:3
	assign Qcnt_two_25 = {Quotient_DP[49:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:974:3
	assign Qcnt_two_26 = {Quotient_DP[51:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:975:3
	assign Qcnt_two_27 = {Quotient_DP[53:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:976:3
	assign Qcnt_two_28 = {Quotient_DP[55:0], Sqrt_quotinent_S[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:979:3
	assign Qcnt_three_0 = {1'b0, Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:980:3
	assign Qcnt_three_1 = {Quotient_DP[2:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:981:3
	assign Qcnt_three_2 = {Quotient_DP[5:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:982:3
	assign Qcnt_three_3 = {Quotient_DP[8:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:983:3
	assign Qcnt_three_4 = {Quotient_DP[11:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:984:3
	assign Qcnt_three_5 = {Quotient_DP[14:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:985:3
	assign Qcnt_three_6 = {Quotient_DP[17:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:986:3
	assign Qcnt_three_7 = {Quotient_DP[20:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:987:3
	assign Qcnt_three_8 = {Quotient_DP[23:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:988:3
	assign Qcnt_three_9 = {Quotient_DP[26:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:989:3
	assign Qcnt_three_10 = {Quotient_DP[29:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:990:3
	assign Qcnt_three_11 = {Quotient_DP[32:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:991:3
	assign Qcnt_three_12 = {Quotient_DP[35:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:992:3
	assign Qcnt_three_13 = {Quotient_DP[38:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:993:3
	assign Qcnt_three_14 = {Quotient_DP[41:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:994:3
	assign Qcnt_three_15 = {Quotient_DP[44:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:995:3
	assign Qcnt_three_16 = {Quotient_DP[47:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:996:3
	assign Qcnt_three_17 = {Quotient_DP[50:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:997:3
	assign Qcnt_three_18 = {Quotient_DP[53:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:998:3
	assign Qcnt_three_19 = {Quotient_DP[56:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1001:3
	assign Qcnt_four_0 = {1'b0, Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1002:3
	assign Qcnt_four_1 = {Quotient_DP[3:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1003:3
	assign Qcnt_four_2 = {Quotient_DP[7:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1004:3
	assign Qcnt_four_3 = {Quotient_DP[11:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1005:3
	assign Qcnt_four_4 = {Quotient_DP[15:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1006:3
	assign Qcnt_four_5 = {Quotient_DP[19:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1007:3
	assign Qcnt_four_6 = {Quotient_DP[23:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1008:3
	assign Qcnt_four_7 = {Quotient_DP[27:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1009:3
	assign Qcnt_four_8 = {Quotient_DP[31:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1010:3
	assign Qcnt_four_9 = {Quotient_DP[35:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1011:3
	assign Qcnt_four_10 = {Quotient_DP[39:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1012:3
	assign Qcnt_four_11 = {Quotient_DP[43:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1013:3
	assign Qcnt_four_12 = {Quotient_DP[47:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1014:3
	assign Qcnt_four_13 = {Quotient_DP[51:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1015:3
	assign Qcnt_four_14 = {Quotient_DP[55:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1020:3
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1022:3
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1033:9
				case (Crtl_cnt_S)
					6'b000000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1037:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1038:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_one_0};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1039:15
						Sqrt_Q0 = Q_sqrt_com_0;
					end
					6'b000001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1043:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[51:50];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1044:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_one_1};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1045:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1049:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[49:48];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1050:15
						Q_sqrt0 = {{56 {1'b0}}, Qcnt_one_2};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1051:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1055:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[47:46];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1056:15
						Q_sqrt0 = {{55 {1'b0}}, Qcnt_one_3};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1057:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1061:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1062:15
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_one_4};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1063:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1067:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[43:42];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1068:15
						Q_sqrt0 = {{53 {1'b0}}, Qcnt_one_5};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1069:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1073:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1074:15
						Q_sqrt0 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_one_6};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1075:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1079:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[39:38];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1080:15
						Q_sqrt0 = {{51 {1'b0}}, Qcnt_one_7};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1081:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1085:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1086:15
						Q_sqrt0 = {{50 {1'b0}}, Qcnt_one_8};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1087:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1091:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[35:34];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1092:15
						Q_sqrt0 = {{49 {1'b0}}, Qcnt_one_9};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1093:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1097:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[33:32];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1098:15
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_one_10};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1099:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1103:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[31:30];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1104:15
						Q_sqrt0 = {{47 {1'b0}}, Qcnt_one_11};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1105:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1109:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1110:15
						Q_sqrt0 = {{46 {1'b0}}, Qcnt_one_12};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1111:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1115:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[27:26];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1116:15
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_one_13};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1117:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1121:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[25:24];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1122:15
						Q_sqrt0 = {{44 {1'b0}}, Qcnt_one_14};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1123:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1127:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[23:22];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1128:15
						Q_sqrt0 = {{43 {1'b0}}, Qcnt_one_15};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1129:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1133:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1134:15
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_one_16};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1135:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1139:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[19:18];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1140:15
						Q_sqrt0 = {{41 {1'b0}}, Qcnt_one_17};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1141:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1145:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1146:15
						Q_sqrt0 = {{40 {1'b0}}, Qcnt_one_18};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1147:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1151:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[15:14];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1152:15
						Q_sqrt0 = {{39 {1'b0}}, Qcnt_one_19};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1153:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1157:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1158:15
						Q_sqrt0 = {{38 {1'b0}}, Qcnt_one_20};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1159:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1163:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[11:10];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1164:15
						Q_sqrt0 = {{37 {1'b0}}, Qcnt_one_21};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1165:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1169:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[9:8];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1170:15
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_one_22};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1171:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1175:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[7:6];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1176:15
						Q_sqrt0 = {{35 {1'b0}}, Qcnt_one_23};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1177:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1181:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1182:15
						Q_sqrt0 = {{34 {1'b0}}, Qcnt_one_24};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1183:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1187:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[3:2];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1188:15
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_one_25};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1189:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1193:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[1:0];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1194:15
						Q_sqrt0 = {{32 {1'b0}}, Qcnt_one_26};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1195:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1199:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1200:15
						Q_sqrt0 = {{31 {1'b0}}, Qcnt_one_27};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1201:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1205:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1206:15
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_one_28};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1207:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1211:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1212:15
						Q_sqrt0 = {{29 {1'b0}}, Qcnt_one_29};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1213:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1217:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1218:15
						Q_sqrt0 = {{28 {1'b0}}, Qcnt_one_30};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1219:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1223:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1224:15
						Q_sqrt0 = {{27 {1'b0}}, Qcnt_one_31};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1225:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1229:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1230:15
						Q_sqrt0 = {{26 {1'b0}}, Qcnt_one_32};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1231:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1235:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1236:15
						Q_sqrt0 = {{25 {1'b0}}, Qcnt_one_33};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1237:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1241:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1242:15
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_one_34};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1243:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1247:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1248:15
						Q_sqrt0 = {{23 {1'b0}}, Qcnt_one_35};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1249:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1253:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1254:15
						Q_sqrt0 = {{22 {1'b0}}, Qcnt_one_36};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1255:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1259:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1260:15
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_one_37};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1261:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1265:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1266:15
						Q_sqrt0 = {{20 {1'b0}}, Qcnt_one_38};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1267:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1271:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1272:15
						Q_sqrt0 = {{19 {1'b0}}, Qcnt_one_39};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1273:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1277:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1278:15
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_one_40};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1279:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1283:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1284:15
						Q_sqrt0 = {{17 {1'b0}}, Qcnt_one_41};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1285:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1289:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1290:15
						Q_sqrt0 = {{16 {1'b0}}, Qcnt_one_42};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1291:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1295:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1296:15
						Q_sqrt0 = {{15 {1'b0}}, Qcnt_one_43};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1297:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1301:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1302:15
						Q_sqrt0 = {{14 {1'b0}}, Qcnt_one_44};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1303:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1307:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1308:15
						Q_sqrt0 = {{13 {1'b0}}, Qcnt_one_45};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1309:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1313:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1314:15
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_one_46};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1315:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1319:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1320:15
						Q_sqrt0 = {{11 {1'b0}}, Qcnt_one_47};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1321:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1325:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1326:15
						Q_sqrt0 = {{10 {1'b0}}, Qcnt_one_48};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1327:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1331:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1332:15
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_one_49};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1333:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1337:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1338:15
						Q_sqrt0 = {{8 {1'b0}}, Qcnt_one_50};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1339:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1343:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1344:15
						Q_sqrt0 = {{7 {1'b0}}, Qcnt_one_51};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1345:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1349:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1350:15
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_one_52};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1351:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1355:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1356:15
						Q_sqrt0 = {{5 {1'b0}}, Qcnt_one_53};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1357:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1361:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1362:15
						Q_sqrt0 = {{4 {1'b0}}, Qcnt_one_54};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1363:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1367:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1368:15
						Q_sqrt0 = {{3 {1'b0}}, Qcnt_one_55};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1369:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b111000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1373:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1374:15
						Q_sqrt0 = {{2 {1'b0}}, Qcnt_one_56};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1375:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					default: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1380:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1381:15
						Q_sqrt0 = 1'sb0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1382:15
						Sqrt_Q0 = 1'sb0;
					end
				endcase
			2'b01:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1398:9
				case (Crtl_cnt_S)
					6'b000000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1402:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1403:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_two_0[1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1404:15
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1405:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1406:15
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_two_0[1:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1407:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1412:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[49:48];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1413:15
						Q_sqrt0 = {{56 {1'b0}}, Qcnt_two_1[2:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1414:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1415:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[47:46];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1416:15
						Q_sqrt1 = {{55 {1'b0}}, Qcnt_two_1[2:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1417:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1422:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1423:15
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_two_2[4:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1424:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1425:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[43:42];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1426:15
						Q_sqrt1 = {{53 {1'b0}}, Qcnt_two_2[4:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1427:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1432:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1433:15
						Q_sqrt0 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_two_3[6:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1434:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1435:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[39:38];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1436:15
						Q_sqrt1 = {{51 {1'b0}}, Qcnt_two_3[6:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1437:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1442:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1443:15
						Q_sqrt0 = {{50 {1'b0}}, Qcnt_two_4[8:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1444:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1445:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[35:34];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1446:15
						Q_sqrt1 = {{49 {1'b0}}, Qcnt_two_4[8:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1447:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1452:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[33:32];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1453:15
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_two_5[10:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1454:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1455:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[31:30];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1456:15
						Q_sqrt1 = {{47 {1'b0}}, Qcnt_two_5[10:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1457:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1462:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1463:15
						Q_sqrt0 = {{46 {1'b0}}, Qcnt_two_6[12:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1464:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1465:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1466:15
						Q_sqrt1 = {{45 {1'b0}}, Qcnt_two_6[12:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1467:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1472:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[25:24];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1473:15
						Q_sqrt0 = {{44 {1'b0}}, Qcnt_two_7[14:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1474:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1475:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[23:22];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1476:15
						Q_sqrt1 = {{43 {1'b0}}, Qcnt_two_7[14:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1477:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1482:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1483:15
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_two_8[16:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1484:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1485:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[19:18];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1486:15
						Q_sqrt1 = {{41 {1'b0}}, Qcnt_two_8[16:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1487:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1492:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1493:15
						Q_sqrt0 = {{40 {1'b0}}, Qcnt_two_9[18:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1494:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1495:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[15:14];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1496:15
						Q_sqrt1 = {{39 {1'b0}}, Qcnt_two_9[18:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1497:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1502:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1503:15
						Q_sqrt0 = {{38 {1'b0}}, Qcnt_two_10[20:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1504:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1505:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[11:10];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1506:15
						Q_sqrt1 = {{37 {1'b0}}, Qcnt_two_10[20:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1507:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1512:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[9:8];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1513:15
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_two_11[22:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1514:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1515:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[7:6];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1516:15
						Q_sqrt1 = {{35 {1'b0}}, Qcnt_two_11[22:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1517:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1522:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1523:15
						Q_sqrt0 = {{34 {1'b0}}, Qcnt_two_12[24:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1524:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1525:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1526:15
						Q_sqrt1 = {{33 {1'b0}}, Qcnt_two_12[24:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1527:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1532:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[1:0];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1533:15
						Q_sqrt0 = {{32 {1'b0}}, Qcnt_two_13[26:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1534:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1535:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1536:15
						Q_sqrt1 = {{31 {1'b0}}, Qcnt_two_13[26:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1537:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1542:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1543:15
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_two_14[28:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1544:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1545:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1546:15
						Q_sqrt1 = {{29 {1'b0}}, Qcnt_two_14[28:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1547:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1552:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1553:15
						Q_sqrt0 = {{28 {1'b0}}, Qcnt_two_15[30:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1554:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1555:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1556:15
						Q_sqrt1 = {{27 {1'b0}}, Qcnt_two_15[30:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1557:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1562:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1563:15
						Q_sqrt0 = {{26 {1'b0}}, Qcnt_two_16[32:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1564:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1565:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1566:15
						Q_sqrt1 = {{25 {1'b0}}, Qcnt_two_16[32:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1567:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1572:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1573:15
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_two_17[34:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1574:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1575:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1576:15
						Q_sqrt1 = {{23 {1'b0}}, Qcnt_two_17[34:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1577:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1582:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1583:15
						Q_sqrt0 = {{22 {1'b0}}, Qcnt_two_18[36:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1584:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1585:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1586:15
						Q_sqrt1 = {{21 {1'b0}}, Qcnt_two_18[36:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1587:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1592:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1593:15
						Q_sqrt0 = {{20 {1'b0}}, Qcnt_two_19[38:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1594:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1595:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1596:15
						Q_sqrt1 = {{19 {1'b0}}, Qcnt_two_19[38:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1597:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1602:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1603:15
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_two_20[40:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1604:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1605:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1606:15
						Q_sqrt1 = {{17 {1'b0}}, Qcnt_two_20[40:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1607:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1612:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1613:15
						Q_sqrt0 = {{16 {1'b0}}, Qcnt_two_21[42:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1614:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1615:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1616:15
						Q_sqrt1 = {{15 {1'b0}}, Qcnt_two_21[42:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1617:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1622:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1623:15
						Q_sqrt0 = {{14 {1'b0}}, Qcnt_two_22[44:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1624:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1625:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1626:15
						Q_sqrt1 = {{13 {1'b0}}, Qcnt_two_22[44:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1627:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1632:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1633:15
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_two_23[46:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1634:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1635:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1636:15
						Q_sqrt1 = {{11 {1'b0}}, Qcnt_two_23[46:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1637:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1642:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1643:15
						Q_sqrt0 = {{10 {1'b0}}, Qcnt_two_24[48:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1644:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1645:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1646:15
						Q_sqrt1 = {{9 {1'b0}}, Qcnt_two_24[48:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1647:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1652:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1653:15
						Q_sqrt0 = {{8 {1'b0}}, Qcnt_two_25[50:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1654:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1655:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1656:15
						Q_sqrt1 = {{7 {1'b0}}, Qcnt_two_25[50:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1657:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1662:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1663:15
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_two_26[52:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1664:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1665:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1666:15
						Q_sqrt1 = {{5 {1'b0}}, Qcnt_two_26[52:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1667:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1672:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1673:15
						Q_sqrt0 = {{4 {1'b0}}, Qcnt_two_27[54:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1674:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1675:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1676:15
						Q_sqrt1 = {{3 {1'b0}}, Qcnt_two_27[54:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1677:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1682:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1683:15
						Q_sqrt0 = {{2 {1'b0}}, Qcnt_two_28[56:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1684:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1685:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1686:15
						Q_sqrt1 = {1'b0, Qcnt_two_28[56:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1687:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					default: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1692:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1693:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_two_0[1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1694:15
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1695:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1696:15
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_two_0[1:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1697:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
				endcase
			2'b10:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1714:9
				case (Crtl_cnt_S)
					6'b000000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1717:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1718:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_three_0[2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1719:15
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1720:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1721:15
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_three_0[2:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1722:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1723:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1724:15
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_three_0[2:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1725:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1730:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[47:46];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1731:15
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_three_1[4:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1732:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1733:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[45:44];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1734:15
						Q_sqrt1 = {{53 {1'b0}}, Qcnt_three_1[4:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1735:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1736:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[43:42];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1737:15
						Q_sqrt2 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_three_1[4:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1738:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1743:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1744:15
						Q_sqrt0 = {{51 {1'b0}}, Qcnt_three_2[7:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1745:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1746:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[39:38];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1747:15
						Q_sqrt1 = {{50 {1'b0}}, Qcnt_three_2[7:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1748:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1749:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[37:36];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1750:15
						Q_sqrt2 = {{49 {1'b0}}, Qcnt_three_2[7:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1751:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1756:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[35:34];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1757:15
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_three_3[10:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1758:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1759:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[33:32];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1760:15
						Q_sqrt1 = {{47 {1'b0}}, Qcnt_three_3[10:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1761:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1762:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[31:30];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1763:15
						Q_sqrt2 = {{46 {1'b0}}, Qcnt_three_3[10:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1764:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1769:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1770:15
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_three_4[13:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1771:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1772:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1773:15
						Q_sqrt1 = {{44 {1'b0}}, Qcnt_three_4[13:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1774:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1775:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[25:24];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1776:15
						Q_sqrt2 = {{43 {1'b0}}, Qcnt_three_4[13:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1777:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1782:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[23:22];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1783:15
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_three_5[16:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1784:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1785:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[21:20];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1786:15
						Q_sqrt1 = {{41 {1'b0}}, Qcnt_three_5[16:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1787:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1788:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[19:18];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1789:15
						Q_sqrt2 = {{40 {1'b0}}, Qcnt_three_5[16:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1790:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1795:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1796:15
						Q_sqrt0 = {{39 {1'b0}}, Qcnt_three_6[19:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1797:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1798:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[15:14];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1799:15
						Q_sqrt1 = {{38 {1'b0}}, Qcnt_three_6[19:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1800:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1801:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[13:12];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1802:15
						Q_sqrt2 = {{37 {1'b0}}, Qcnt_three_6[19:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1803:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1808:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[11:10];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1809:15
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_three_7[22:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1810:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1811:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[9:8];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1812:15
						Q_sqrt1 = {{35 {1'b0}}, Qcnt_three_7[22:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1813:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1814:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[7:6];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1815:15
						Q_sqrt2 = {{34 {1'b0}}, Qcnt_three_7[22:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1816:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1821:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1822:15
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_three_8[25:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1823:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1824:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1825:15
						Q_sqrt1 = {{32 {1'b0}}, Qcnt_three_8[25:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1826:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1827:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[1:0];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1828:15
						Q_sqrt2 = {{31 {1'b0}}, Qcnt_three_8[25:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1829:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1834:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1835:15
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_three_9[28:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1836:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1837:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1838:15
						Q_sqrt1 = {{29 {1'b0}}, Qcnt_three_9[28:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1839:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1840:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1841:15
						Q_sqrt2 = {{28 {1'b0}}, Qcnt_three_9[28:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1842:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1847:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1848:15
						Q_sqrt0 = {{27 {1'b0}}, Qcnt_three_10[31:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1849:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1850:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1851:15
						Q_sqrt1 = {{26 {1'b0}}, Qcnt_three_10[31:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1852:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1853:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1854:15
						Q_sqrt2 = {{25 {1'b0}}, Qcnt_three_10[31:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1855:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1860:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1861:15
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_three_11[34:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1862:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1863:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1864:15
						Q_sqrt1 = {{23 {1'b0}}, Qcnt_three_11[34:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1865:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1866:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1867:15
						Q_sqrt2 = {{22 {1'b0}}, Qcnt_three_11[34:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1868:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1873:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1874:15
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_three_12[37:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1875:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1876:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1877:15
						Q_sqrt1 = {{20 {1'b0}}, Qcnt_three_12[37:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1878:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1879:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1880:15
						Q_sqrt2 = {{19 {1'b0}}, Qcnt_three_12[37:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1881:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1886:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1887:15
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_three_13[40:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1888:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1889:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1890:15
						Q_sqrt1 = {{17 {1'b0}}, Qcnt_three_13[40:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1891:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1892:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1893:15
						Q_sqrt2 = {{16 {1'b0}}, Qcnt_three_13[40:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1894:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1899:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1900:15
						Q_sqrt0 = {{15 {1'b0}}, Qcnt_three_14[43:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1901:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1902:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1903:15
						Q_sqrt1 = {{14 {1'b0}}, Qcnt_three_14[43:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1904:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1905:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1906:15
						Q_sqrt2 = {{13 {1'b0}}, Qcnt_three_14[43:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1907:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1912:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1913:15
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_three_15[46:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1914:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1915:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1916:15
						Q_sqrt1 = {{11 {1'b0}}, Qcnt_three_15[46:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1917:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1918:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1919:15
						Q_sqrt2 = {{10 {1'b0}}, Qcnt_three_15[46:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1920:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1925:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1926:15
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_three_16[49:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1927:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1928:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1929:15
						Q_sqrt1 = {{8 {1'b0}}, Qcnt_three_16[49:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1930:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1931:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1932:15
						Q_sqrt2 = {{7 {1'b0}}, Qcnt_three_16[49:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1933:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1938:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1939:15
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_three_17[52:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1940:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1941:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1942:15
						Q_sqrt1 = {{5 {1'b0}}, Qcnt_three_17[52:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1943:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1944:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1945:15
						Q_sqrt2 = {{4 {1'b0}}, Qcnt_three_17[52:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1946:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1951:15
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1952:15
						Q_sqrt0 = {{3 {1'b0}}, Qcnt_three_18[55:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1953:15
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1954:15
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1955:15
						Q_sqrt1 = {{2 {1'b0}}, Qcnt_three_18[55:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1956:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1957:15
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1958:15
						Q_sqrt2 = {1'b0, Qcnt_three_18[55:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1959:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					default: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1964:15
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1965:15
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_three_0[2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1966:15
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1967:15
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1968:15
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_three_0[2:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1969:15
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1970:15
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1971:15
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_three_0[2:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1972:15
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
				endcase
			2'b11:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1988:15
				case (Crtl_cnt_S)
					6'b000000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1992:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1993:21
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_four_0[3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1994:21
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1995:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1996:21
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_four_0[3:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1997:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1998:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:1999:21
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_four_0[3:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2000:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2001:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[47:46];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2002:21
						Q_sqrt3 = {{54 {1'b0}}, Qcnt_four_0[3:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2003:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2008:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2009:21
						Q_sqrt0 = {{53 {1'b0}}, Qcnt_four_1[6:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2010:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2011:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[43:42];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2012:21
						Q_sqrt1 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_four_1[6:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2013:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2014:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[41:40];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2015:21
						Q_sqrt2 = {{51 {1'b0}}, Qcnt_four_1[6:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2016:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2017:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[39:38];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2018:21
						Q_sqrt3 = {{50 {1'b0}}, Qcnt_four_1[6:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2019:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2024:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2025:21
						Q_sqrt0 = {{49 {1'b0}}, Qcnt_four_2[10:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2026:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2027:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[35:34];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2028:21
						Q_sqrt1 = {{48 {1'b0}}, Qcnt_four_2[10:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2029:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2030:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[33:32];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2031:21
						Q_sqrt2 = {{47 {1'b0}}, Qcnt_four_2[10:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2032:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2033:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[31:30];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2034:21
						Q_sqrt3 = {{46 {1'b0}}, Qcnt_four_2[10:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2035:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2040:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2041:21
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_four_3[14:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2042:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2043:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2044:21
						Q_sqrt1 = {{44 {1'b0}}, Qcnt_four_3[14:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2045:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2046:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[25:24];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2047:21
						Q_sqrt2 = {{43 {1'b0}}, Qcnt_four_3[14:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2048:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2049:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[23:22];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2050:21
						Q_sqrt3 = {{42 {1'b0}}, Qcnt_four_3[14:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2051:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2056:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2057:21
						Q_sqrt0 = {{41 {1'b0}}, Qcnt_four_4[18:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2058:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2059:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[19:18];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2060:21
						Q_sqrt1 = {{40 {1'b0}}, Qcnt_four_4[18:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2061:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2062:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[17:16];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2063:21
						Q_sqrt2 = {{39 {1'b0}}, Qcnt_four_4[18:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2064:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2065:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[15:14];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2066:21
						Q_sqrt3 = {{38 {1'b0}}, Qcnt_four_4[18:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2067:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2072:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2073:21
						Q_sqrt0 = {{37 {1'b0}}, Qcnt_four_5[22:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2074:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2075:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[11:10];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2076:21
						Q_sqrt1 = {{36 {1'b0}}, Qcnt_four_5[22:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2077:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2078:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[9:8];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2079:21
						Q_sqrt2 = {{35 {1'b0}}, Qcnt_four_5[22:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2080:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2081:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[7:6];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2082:21
						Q_sqrt3 = {{34 {1'b0}}, Qcnt_four_5[22:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2083:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000110: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2088:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2089:21
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_four_6[26:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2090:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2091:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2092:21
						Q_sqrt1 = {{32 {1'b0}}, Qcnt_four_6[26:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2093:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2094:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[1:0];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2095:21
						Q_sqrt2 = {{31 {1'b0}}, Qcnt_four_6[26:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2096:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2097:21
						Sqrt_DI[3] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2098:21
						Q_sqrt3 = {{30 {1'b0}}, Qcnt_four_6[26:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2099:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000111: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2104:21
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2105:21
						Q_sqrt0 = {{29 {1'b0}}, Qcnt_four_7[30:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2106:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2107:21
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2108:21
						Q_sqrt1 = {{28 {1'b0}}, Qcnt_four_7[30:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2109:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2110:21
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2111:21
						Q_sqrt2 = {{27 {1'b0}}, Qcnt_four_7[30:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2112:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2113:21
						Sqrt_DI[3] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2114:21
						Q_sqrt3 = {{26 {1'b0}}, Qcnt_four_7[30:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2115:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001000: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2120:21
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2121:21
						Q_sqrt0 = {{25 {1'b0}}, Qcnt_four_8[34:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2122:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2123:21
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2124:21
						Q_sqrt1 = {{24 {1'b0}}, Qcnt_four_8[34:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2125:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2126:21
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2127:21
						Q_sqrt2 = {{23 {1'b0}}, Qcnt_four_8[34:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2128:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2129:21
						Sqrt_DI[3] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2130:21
						Q_sqrt3 = {{22 {1'b0}}, Qcnt_four_8[34:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2131:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001001: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2136:21
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2137:21
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_four_9[38:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2138:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2139:21
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2140:21
						Q_sqrt1 = {{20 {1'b0}}, Qcnt_four_9[38:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2141:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2142:21
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2143:21
						Q_sqrt2 = {{19 {1'b0}}, Qcnt_four_9[38:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2144:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2145:21
						Sqrt_DI[3] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2146:21
						Q_sqrt3 = {{18 {1'b0}}, Qcnt_four_9[38:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2147:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001010: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2152:21
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2153:21
						Q_sqrt0 = {{17 {1'b0}}, Qcnt_four_10[42:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2154:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2155:21
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2156:21
						Q_sqrt1 = {{16 {1'b0}}, Qcnt_four_10[42:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2157:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2158:21
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2159:21
						Q_sqrt2 = {{15 {1'b0}}, Qcnt_four_10[42:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2160:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2161:21
						Sqrt_DI[3] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2162:21
						Q_sqrt3 = {{14 {1'b0}}, Qcnt_four_10[42:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2163:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001011: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2168:21
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2169:21
						Q_sqrt0 = {{13 {1'b0}}, Qcnt_four_11[46:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2170:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2171:21
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2172:21
						Q_sqrt1 = {{12 {1'b0}}, Qcnt_four_11[46:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2173:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2174:21
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2175:21
						Q_sqrt2 = {{11 {1'b0}}, Qcnt_four_11[46:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2176:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2177:21
						Sqrt_DI[3] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2178:21
						Q_sqrt3 = {{10 {1'b0}}, Qcnt_four_11[46:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2179:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001100: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2184:21
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2185:21
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_four_12[50:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2186:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2187:21
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2188:21
						Q_sqrt1 = {{8 {1'b0}}, Qcnt_four_12[50:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2189:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2190:21
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2191:21
						Q_sqrt2 = {{7 {1'b0}}, Qcnt_four_12[50:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2192:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2193:21
						Sqrt_DI[3] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2194:21
						Q_sqrt3 = {{6 {1'b0}}, Qcnt_four_12[50:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2195:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001101: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2200:21
						Sqrt_DI[0] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2201:21
						Q_sqrt0 = {{5 {1'b0}}, Qcnt_four_13[54:3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2202:21
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2203:21
						Sqrt_DI[1] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2204:21
						Q_sqrt1 = {{4 {1'b0}}, Qcnt_four_13[54:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2205:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2206:21
						Sqrt_DI[2] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2207:21
						Q_sqrt2 = {{3 {1'b0}}, Qcnt_four_13[54:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2208:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2209:21
						Sqrt_DI[3] = 2'b00;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2210:21
						Q_sqrt3 = {{2 {1'b0}}, Qcnt_four_13[54:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2211:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					default: begin
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2216:21
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2217:21
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_four_0[3]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2218:21
						Sqrt_Q0 = Q_sqrt_com_0;
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2219:21
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2220:21
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_four_0[3:2]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2221:21
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2222:21
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2223:21
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_four_0[3:1]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2224:21
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2225:21
						Sqrt_DI[3] = Mant_D_sqrt_Norm[47:46];
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2226:21
						Q_sqrt3 = {{54 {1'b0}}, Qcnt_four_0[3:0]};
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2227:21
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
				endcase
		endcase
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2239:3
	assign Sqrt_R0 = (Sqrt_start_dly_S ? {58 {1'sb0}} : {Partial_remainder_DP[57:0]});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2240:3
	assign Sqrt_R1 = {Iteration_cell_sum_AMASK_D[0][57], Iteration_cell_sum_AMASK_D[0][54:0], Sqrt_DO[0]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2241:3
	assign Sqrt_R2 = {Iteration_cell_sum_AMASK_D[1][57], Iteration_cell_sum_AMASK_D[1][54:0], Sqrt_DO[1]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2242:3
	assign Sqrt_R3 = {Iteration_cell_sum_AMASK_D[2][57], Iteration_cell_sum_AMASK_D[2][54:0], Sqrt_DO[2]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2243:3
	assign Sqrt_R4 = {Iteration_cell_sum_AMASK_D[3][57], Iteration_cell_sum_AMASK_D[3][54:0], Sqrt_DO[3]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2245:3
	wire [57:0] Denominator_se_format_DB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2247:3
	assign Denominator_se_format_DB = {Denominator_se_DB[53:45], (FP16ALT_SO ? FP16ALT_SO : Denominator_se_DB[44]), Denominator_se_DB[43:42], (FP16_SO ? FP16_SO : Denominator_se_DB[41]), Denominator_se_DB[40:29], (FP32_SO ? FP32_SO : Denominator_se_DB[28]), Denominator_se_DB[27:0], FP64_SO, 3'b000};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2252:3
	wire [57:0] First_iteration_cell_div_a_D;
	wire [57:0] First_iteration_cell_div_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2253:3
	wire Sel_b_for_first_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2256:3
	assign First_iteration_cell_div_a_D = (Div_start_dly_S ? {Numerator_se_D[53:45], (FP16ALT_SO ? FP16ALT_SO : Numerator_se_D[44]), Numerator_se_D[43:42], (FP16_SO ? FP16_SO : Numerator_se_D[41]), Numerator_se_D[40:29], (FP32_SO ? FP32_SO : Numerator_se_D[28]), Numerator_se_D[27:0], FP64_SO, 3'b000} : {Partial_remainder_DP[56:48], (FP16ALT_SO ? Quotient_DP[0] : Partial_remainder_DP[47]), Partial_remainder_DP[46:45], (FP16_SO ? Quotient_DP[0] : Partial_remainder_DP[44]), Partial_remainder_DP[43:32], (FP32_SO ? Quotient_DP[0] : Partial_remainder_DP[31]), Partial_remainder_DP[30:3], FP64_SO && Quotient_DP[0], 3'b000});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2264:3
	assign Sel_b_for_first_S = (Div_start_dly_S ? 1 : Quotient_DP[0]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2265:3
	assign First_iteration_cell_div_b_D = (Sel_b_for_first_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2266:3
	assign Iteration_cell_a_BMASK_D[0] = (Sqrt_enable_SO ? Sqrt_R0 : {First_iteration_cell_div_a_D});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2267:3
	assign Iteration_cell_b_BMASK_D[0] = (Sqrt_enable_SO ? Sqrt_Q0 : {First_iteration_cell_div_b_D});
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2272:3
	wire [57:0] Sec_iteration_cell_div_a_D;
	wire [57:0] Sec_iteration_cell_div_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2273:3
	wire Sel_b_for_sec_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2274:3
	generate
		if (|defs_div_sqrt_mvp_Iteration_unit_num_S) begin : genblk1
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2277:9
			assign Sel_b_for_sec_S = ~Iteration_cell_sum_AMASK_D[0][57];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2278:9
			assign Sec_iteration_cell_div_a_D = {Iteration_cell_sum_AMASK_D[0][56:48], (FP16ALT_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][47]), Iteration_cell_sum_AMASK_D[0][46:45], (FP16_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][44]), Iteration_cell_sum_AMASK_D[0][43:32], (FP32_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][31]), Iteration_cell_sum_AMASK_D[0][30:3], FP64_SO && Sel_b_for_sec_S, 3'b000};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2282:9
			assign Sec_iteration_cell_div_b_D = (Sel_b_for_sec_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2283:9
			assign Iteration_cell_a_BMASK_D[1] = (Sqrt_enable_SO ? Sqrt_R1 : {Sec_iteration_cell_div_a_D});
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2284:9
			assign Iteration_cell_b_BMASK_D[1] = (Sqrt_enable_SO ? Sqrt_Q1 : {Sec_iteration_cell_div_b_D});
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2289:3
	wire [57:0] Thi_iteration_cell_div_a_D;
	wire [57:0] Thi_iteration_cell_div_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2290:3
	wire Sel_b_for_thi_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2291:3
	generate
		if (1'd1 | 1'd0) begin : genblk2
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2294:9
			assign Sel_b_for_thi_S = ~Iteration_cell_sum_AMASK_D[1][57];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2295:9
			assign Thi_iteration_cell_div_a_D = {Iteration_cell_sum_AMASK_D[1][56:48], (FP16ALT_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][47]), Iteration_cell_sum_AMASK_D[1][46:45], (FP16_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][44]), Iteration_cell_sum_AMASK_D[1][43:32], (FP32_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][31]), Iteration_cell_sum_AMASK_D[1][30:3], FP64_SO && Sel_b_for_thi_S, 3'b000};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2299:9
			assign Thi_iteration_cell_div_b_D = (Sel_b_for_thi_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2300:9
			assign Iteration_cell_a_BMASK_D[2] = (Sqrt_enable_SO ? Sqrt_R2 : {Thi_iteration_cell_div_a_D});
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2301:9
			assign Iteration_cell_b_BMASK_D[2] = (Sqrt_enable_SO ? Sqrt_Q2 : {Thi_iteration_cell_div_b_D});
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2306:3
	wire [57:0] Fou_iteration_cell_div_a_D;
	wire [57:0] Fou_iteration_cell_div_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2307:3
	wire Sel_b_for_fou_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2309:3
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2328:3
	wire [57:0] Mask_bits_ctl_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2330:3
	assign Mask_bits_ctl_S = 58'h3ffffffffffffff;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2337:3
	wire Div_enable_SI [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2338:3
	wire Div_start_dly_SI [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2339:3
	wire Sqrt_enable_SI [3:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2340:3
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2341:5
	genvar i;
	genvar j;
	generate
		for (i = 0; i <= defs_div_sqrt_mvp_Iteration_unit_num_S; i = i + 1) begin : genblk4
			for (j = 0; j <= 57; j = j + 1) begin : genblk1
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2345:15
				assign Iteration_cell_a_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_a_BMASK_D[i][j];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2346:15
				assign Iteration_cell_b_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_b_BMASK_D[i][j];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2347:15
				assign Iteration_cell_sum_AMASK_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_sum_D[i][j];
			end
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2350:11
			assign Div_enable_SI[i] = Div_enable_SO;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2351:11
			assign Div_start_dly_SI[i] = Div_start_dly_S;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2352:11
			assign Sqrt_enable_SI[i] = Sqrt_enable_SO;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2353:11
			iteration_div_sqrt_mvp #(.WIDTH(58)) iteration_div_sqrt(
				.A_DI(Iteration_cell_a_D[i]),
				.B_DI(Iteration_cell_b_D[i]),
				.Div_enable_SI(Div_enable_SI[i]),
				.Div_start_dly_SI(Div_start_dly_SI[i]),
				.Sqrt_enable_SI(Sqrt_enable_SI[i]),
				.D_DI(Sqrt_DI[i]),
				.D_DO(Sqrt_DO[i]),
				.Sum_DO(Iteration_cell_sum_D[i]),
				.Carry_out_DO(Iteration_cell_carry_D[i])
			);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2372:3
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2374:7
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2377:13
				if (Fsm_enable_S)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2378:16
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R1 : Iteration_cell_sum_AMASK_D[0]);
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2380:16
					Partial_remainder_DN = Partial_remainder_DP;
			2'b01:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2384:13
				if (Fsm_enable_S)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2385:16
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R2 : Iteration_cell_sum_AMASK_D[1]);
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2387:16
					Partial_remainder_DN = Partial_remainder_DP;
			2'b10:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2391:13
				if (Fsm_enable_S)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2392:16
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R3 : Iteration_cell_sum_AMASK_D[2]);
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2394:16
					Partial_remainder_DN = Partial_remainder_DP;
			2'b11:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2398:13
				if (Fsm_enable_S)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2399:16
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R4 : Iteration_cell_sum_AMASK_D[3]);
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2401:16
					Partial_remainder_DN = Partial_remainder_DP;
		endcase
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2408:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2410:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2412:14
			Partial_remainder_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2416:14
			Partial_remainder_DP <= Partial_remainder_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2420:4
	reg [56:0] Quotient_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2422:3
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2424:7
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2427:13
				if (Fsm_enable_S)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2428:16
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[55:0], Sqrt_quotinent_S[3]} : {Quotient_DP[55:0], Iteration_cell_carry_D[0]});
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2430:16
					Quotient_DN = Quotient_DP;
			2'b01:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2434:13
				if (Fsm_enable_S)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2435:16
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[54:0], Sqrt_quotinent_S[3:2]} : {Quotient_DP[54:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1]});
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2437:16
					Quotient_DN = Quotient_DP;
			2'b10:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2441:13
				if (Fsm_enable_S)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2442:16
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[53:0], Sqrt_quotinent_S[3:1]} : {Quotient_DP[53:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2]});
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2444:16
					Quotient_DN = Quotient_DP;
			2'b11:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2448:13
				if (Fsm_enable_S)
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2449:16
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP64:0], Sqrt_quotinent_S} : {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP64:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2], Iteration_cell_carry_D[3]});
				else
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2451:16
					Quotient_DN = Quotient_DP;
		endcase
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2456:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2458:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2460:11
			Quotient_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2463:11
			Quotient_DP <= Quotient_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2473:4
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:2814:4
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3030:4
	generate
		if (1) begin : genblk7
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3033:9
			always @(*)
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3035:13
				case (Format_sel_S)
					2'b00:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3038:19
						case (Precision_ctl_S)
							6'h00:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3041:25
								Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
							6'h17, 6'h16, 6'h15:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3045:25
								Mant_result_prenorm_DO = {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP32:0], {33 {1'b0}}};
							6'h14, 6'h13, 6'h12:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3049:25
								Mant_result_prenorm_DO = {Quotient_DP[20:0], {36 {1'b0}}};
							6'h11, 6'h10, 6'h0f:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3053:25
								Mant_result_prenorm_DO = {Quotient_DP[17:0], {39 {1'b0}}};
							6'h0e, 6'h0d, 6'h0c:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3057:25
								Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0b, 6'h0a, 6'h09:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3061:25
								Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h08, 6'h07, 6'h06:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3065:25
								Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3069:25
								Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
						endcase
					2'b01:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3076:19
						case (Precision_ctl_S)
							6'h00:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3079:25
								Mant_result_prenorm_DO = Quotient_DP[56:0];
							6'h34, 6'h33:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3083:25
								Mant_result_prenorm_DO = {Quotient_DP[53:1], {4 {1'b0}}};
							6'h32, 6'h31, 6'h30:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3087:25
								Mant_result_prenorm_DO = {Quotient_DP[50:0], {6 {1'b0}}};
							6'h2f, 6'h2e, 6'h2d:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3091:25
								Mant_result_prenorm_DO = {Quotient_DP[47:0], {9 {1'b0}}};
							6'h2c, 6'h2b, 6'h2a:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3095:25
								Mant_result_prenorm_DO = {Quotient_DP[44:0], {12 {1'b0}}};
							6'h29, 6'h28, 6'h27:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3099:25
								Mant_result_prenorm_DO = {Quotient_DP[41:0], {15 {1'b0}}};
							6'h26, 6'h25, 6'h24:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3103:25
								Mant_result_prenorm_DO = {Quotient_DP[38:0], {18 {1'b0}}};
							6'h23, 6'h22, 6'h21:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3107:25
								Mant_result_prenorm_DO = {Quotient_DP[35:0], {21 {1'b0}}};
							6'h20, 6'h1f, 6'h1e:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3111:25
								Mant_result_prenorm_DO = {Quotient_DP[32:0], {24 {1'b0}}};
							6'h1d, 6'h1c, 6'h1b:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3115:25
								Mant_result_prenorm_DO = {Quotient_DP[29:0], {27 {1'b0}}};
							6'h1a, 6'h19, 6'h18:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3119:25
								Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
							6'h17, 6'h16, 6'h15:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3123:25
								Mant_result_prenorm_DO = {Quotient_DP[23:0], {33 {1'b0}}};
							6'h14, 6'h13, 6'h12:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3127:25
								Mant_result_prenorm_DO = {Quotient_DP[20:0], {36 {1'b0}}};
							6'h11, 6'h10, 6'h0f:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3131:25
								Mant_result_prenorm_DO = {Quotient_DP[17:0], {39 {1'b0}}};
							6'h0e, 6'h0d, 6'h0c:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3135:25
								Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0b, 6'h0a, 6'h09:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3139:25
								Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h08, 6'h07, 6'h06:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3143:25
								Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3147:25
								Mant_result_prenorm_DO = Quotient_DP[56:0];
						endcase
					2'b10:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3154:19
						case (Precision_ctl_S)
							6'b000000:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3157:25
								Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0a, 6'h09:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3161:25
								Mant_result_prenorm_DO = {Quotient_DP[11:1], {46 {1'b0}}};
							6'h08, 6'h07, 6'h06:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3165:25
								Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3169:25
								Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
						endcase
					2'b11:
						// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3177:19
						case (Precision_ctl_S)
							6'b000000:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3180:25
								Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h07, 6'h06:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3184:25
								Mant_result_prenorm_DO = {Quotient_DP[8:1], {49 {1'b0}}};
							default:
								// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3188:25
								Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
						endcase
				endcase
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3199:4
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3356:4
	wire [12:0] Exp_result_prenorm_DN;
	reg [12:0] Exp_result_prenorm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3358:4
	wire [12:0] Exp_add_a_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3359:4
	wire [12:0] Exp_add_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3360:4
	wire [12:0] Exp_add_c_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3362:3
	integer C_BIAS_AONE;
	integer C_HALF_BIAS;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3363:3
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP16 = 5'h10;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP16ALT = 8'h80;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP32 = 8'h80;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP64 = 11'h400;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP16 = 7;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP16ALT = 63;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP32 = 63;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP64 = 511;
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3365:7
		case (Format_sel_S)
			2'b00: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3368:13
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP32;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3369:13
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP32;
			end
			2'b01: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3373:13
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP64;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3374:13
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP64;
			end
			2'b10: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3378:13
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP16;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3379:13
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP16;
			end
			2'b11: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3383:13
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP16ALT;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3384:13
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP16ALT;
			end
		endcase
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3393:3
	assign Exp_add_a_D = {(Sqrt_start_dly_S ? {Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64:1]} : {Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI})};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3394:3
	localparam defs_div_sqrt_mvp_C_EXP_ZERO_FP64 = 11'h000;
	assign Exp_add_b_D = {(Sqrt_start_dly_S ? {1'b0, defs_div_sqrt_mvp_C_EXP_ZERO_FP64, Exp_num_DI[0]} : {~Exp_den_DI[defs_div_sqrt_mvp_C_EXP_FP64], ~Exp_den_DI[defs_div_sqrt_mvp_C_EXP_FP64], ~Exp_den_DI})};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3395:3
	assign Exp_add_c_D = {(Div_start_dly_S ? {C_BIAS_AONE} : {C_HALF_BIAS})};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3396:3
	assign Exp_result_prenorm_DN = (Start_dly_S ? {(Exp_add_a_D + Exp_add_b_D) + Exp_add_c_D} : Exp_result_prenorm_DP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3399:3
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3401:7
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3403:11
			Exp_result_prenorm_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3407:11
			Exp_result_prenorm_DP <= Exp_result_prenorm_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/control_mvp.sv:3411:3
	assign Exp_result_prenorm_DO = Exp_result_prenorm_DP;
endmodule
// removed package "defs_div_sqrt_mvp"
// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:39:1
// removed ["import defs_div_sqrt_mvp::*;"]
module div_sqrt_mvp_wrapper (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Operand_a_DI,
	Operand_b_DI,
	RM_SI,
	Precision_ctl_SI,
	Format_sel_SI,
	Kill_SI,
	Result_DO,
	Fflags_SO,
	Ready_SO,
	Done_SO
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:43:16
	parameter PrePipeline_depth_S = 0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:44:16
	parameter PostPipeline_depth_S = 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:47:4
	input wire Clk_CI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:48:4
	input wire Rst_RBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:49:4
	input wire Div_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:50:4
	input wire Sqrt_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:53:4
	localparam defs_div_sqrt_mvp_C_OP_FP64 = 64;
	input wire [63:0] Operand_a_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:54:4
	input wire [63:0] Operand_b_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:57:4
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:58:4
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:59:4
	localparam defs_div_sqrt_mvp_C_FS = 2;
	input wire [1:0] Format_sel_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:60:4
	input wire Kill_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:63:4
	output wire [63:0] Result_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:66:4
	output wire [4:0] Fflags_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:67:4
	output wire Ready_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:68:4
	output wire Done_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:72:4
	reg Div_start_S_S;
	reg Sqrt_start_S_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:73:4
	reg [63:0] Operand_a_S_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:74:4
	reg [63:0] Operand_b_S_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:77:4
	reg [2:0] RM_S_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:78:4
	reg [5:0] Precision_ctl_S_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:79:4
	reg [1:0] Format_sel_S_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:80:4
	reg Kill_S_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:83:3
	wire [63:0] Result_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:84:3
	wire Ready_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:85:3
	wire Done_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:86:3
	wire [4:0] Fflags_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:89:3
	generate
		if (PrePipeline_depth_S == 1) begin : genblk1
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:93:10
			div_sqrt_top_mvp div_top_U0(
				.Clk_CI(Clk_CI),
				.Rst_RBI(Rst_RBI),
				.Div_start_SI(Div_start_S_S),
				.Sqrt_start_SI(Sqrt_start_S_S),
				.Operand_a_DI(Operand_a_S_D),
				.Operand_b_DI(Operand_b_S_D),
				.RM_SI(RM_S_S),
				.Precision_ctl_SI(Precision_ctl_S_S),
				.Format_sel_SI(Format_sel_S_S),
				.Kill_SI(Kill_S_S),
				.Result_DO(Result_D),
				.Fflags_SO(Fflags_S),
				.Ready_SO(Ready_S),
				.Done_SO(Done_S)
			);
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:113:12
			always @(posedge Clk_CI or negedge Rst_RBI)
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:115:17
				if (~Rst_RBI) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:117:21
					Div_start_S_S <= 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:118:21
					Sqrt_start_S_S <= 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:119:21
					Operand_a_S_D <= 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:120:21
					Operand_b_S_D <= 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:121:21
					RM_S_S <= 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:122:21
					Precision_ctl_S_S <= 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:123:21
					Format_sel_S_S <= 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:124:21
					Kill_S_S <= 1'sb0;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:128:21
					Div_start_S_S <= Div_start_SI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:129:21
					Sqrt_start_S_S <= Sqrt_start_SI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:130:21
					Operand_a_S_D <= Operand_a_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:131:21
					Operand_b_S_D <= Operand_b_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:132:21
					RM_S_S <= RM_SI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:133:21
					Precision_ctl_S_S <= Precision_ctl_SI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:134:21
					Format_sel_S_S <= Format_sel_SI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:135:21
					Kill_S_S <= Kill_SI;
				end
		end
		else begin : genblk1
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:142:11
			div_sqrt_top_mvp div_top_U0(
				.Clk_CI(Clk_CI),
				.Rst_RBI(Rst_RBI),
				.Div_start_SI(Div_start_SI),
				.Sqrt_start_SI(Sqrt_start_SI),
				.Operand_a_DI(Operand_a_DI),
				.Operand_b_DI(Operand_b_DI),
				.RM_SI(RM_SI),
				.Precision_ctl_SI(Precision_ctl_SI),
				.Format_sel_SI(Format_sel_SI),
				.Kill_SI(Kill_SI),
				.Result_DO(Result_D),
				.Fflags_SO(Fflags_S),
				.Ready_SO(Ready_S),
				.Done_SO(Done_S)
			);
		end
	endgenerate
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:166:3
	reg [63:0] Result_dly_S_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:167:3
	reg Ready_dly_S_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:168:3
	reg Done_dly_S_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:169:3
	reg [4:0] Fflags_dly_S_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:170:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:172:9
		if (~Rst_RBI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:174:13
			Result_dly_S_D <= 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:175:13
			Ready_dly_S_S <= 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:176:13
			Done_dly_S_S <= 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:177:13
			Fflags_dly_S_S <= 1'b0;
		end
		else begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:181:13
			Result_dly_S_D <= Result_D;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:182:13
			Ready_dly_S_S <= Ready_S;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:183:13
			Done_dly_S_S <= Done_S;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:184:13
			Fflags_dly_S_S <= Fflags_S;
		end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:192:3
	reg [63:0] Result_dly_D_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:193:3
	reg Ready_dly_D_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:194:3
	reg Done_dly_D_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:195:3
	reg [4:0] Fflags_dly_D_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:196:3
	generate
		if (PostPipeline_depth_S == 2) begin : genblk2
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:199:9
			always @(posedge Clk_CI or negedge Rst_RBI)
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:201:13
				if (~Rst_RBI) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:203:17
					Result_dly_D_D <= 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:204:17
					Ready_dly_D_S <= 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:205:17
					Done_dly_D_S <= 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:206:17
					Fflags_dly_D_S <= 1'b0;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:210:16
					Result_dly_D_D <= Result_dly_S_D;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:211:16
					Ready_dly_D_S <= Ready_dly_S_S;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:212:16
					Done_dly_D_S <= Done_dly_S_S;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:213:16
					Fflags_dly_D_S <= Fflags_dly_S_S;
				end
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:216:9
			assign Result_DO = Result_dly_D_D;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:217:9
			assign Ready_SO = Ready_dly_D_S;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:218:9
			assign Done_SO = Done_dly_D_S;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:219:9
			assign Fflags_SO = Fflags_dly_D_S;
		end
		else begin : genblk2
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:224:10
			assign Result_DO = Result_dly_S_D;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:225:10
			assign Ready_SO = Ready_dly_S_S;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:226:10
			assign Done_SO = Done_dly_S_S;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_mvp_wrapper.sv:227:10
			assign Fflags_SO = Fflags_dly_S_S;
		end
	endgenerate
endmodule
// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:35:1
// removed ["import defs_div_sqrt_mvp::*;"]
module div_sqrt_top_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Operand_a_DI,
	Operand_b_DI,
	RM_SI,
	Precision_ctl_SI,
	Format_sel_SI,
	Kill_SI,
	Result_DO,
	Fflags_SO,
	Ready_SO,
	Done_SO
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:40:4
	input wire Clk_CI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:41:4
	input wire Rst_RBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:42:4
	input wire Div_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:43:4
	input wire Sqrt_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:46:4
	localparam defs_div_sqrt_mvp_C_OP_FP64 = 64;
	input wire [63:0] Operand_a_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:47:4
	input wire [63:0] Operand_b_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:50:4
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:51:4
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:52:4
	localparam defs_div_sqrt_mvp_C_FS = 2;
	input wire [1:0] Format_sel_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:53:4
	input wire Kill_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:56:4
	output wire [63:0] Result_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:59:4
	output wire [4:0] Fflags_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:60:4
	output wire Ready_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:61:4
	output wire Done_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:69:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:70:4
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:71:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:72:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:74:4
	wire [12:0] Exp_z_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:75:4
	wire [56:0] Mant_z_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:76:4
	wire Sign_z_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:77:4
	wire Start_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:78:4
	wire [2:0] RM_dly_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:79:4
	wire Div_enable_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:80:4
	wire Sqrt_enable_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:81:4
	wire Inf_a_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:82:4
	wire Inf_b_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:83:4
	wire Zero_a_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:84:4
	wire Zero_b_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:85:4
	wire NaN_a_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:86:4
	wire NaN_b_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:87:4
	wire SNaN_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:88:4
	wire Special_case_SB;
	wire Special_case_dly_SB;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:90:4
	wire Full_precision_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:91:4
	wire FP32_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:92:4
	wire FP64_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:93:4
	wire FP16_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:94:4
	wire FP16ALT_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:97:2
	preprocess_mvp preprocess_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Ready_SI(Ready_SO),
		.Operand_a_DI(Operand_a_DI),
		.Operand_b_DI(Operand_b_DI),
		.RM_SI(RM_SI),
		.Format_sel_SI(Format_sel_SI),
		.Start_SO(Start_S),
		.Exp_a_DO_norm(Exp_a_D),
		.Exp_b_DO_norm(Exp_b_D),
		.Mant_a_DO_norm(Mant_a_D),
		.Mant_b_DO_norm(Mant_b_D),
		.RM_dly_SO(RM_dly_S),
		.Sign_z_DO(Sign_z_D),
		.Inf_a_SO(Inf_a_S),
		.Inf_b_SO(Inf_b_S),
		.Zero_a_SO(Zero_a_S),
		.Zero_b_SO(Zero_b_S),
		.NaN_a_SO(NaN_a_S),
		.NaN_b_SO(NaN_b_S),
		.SNaN_SO(SNaN_S),
		.Special_case_SBO(Special_case_SB),
		.Special_case_dly_SBO(Special_case_dly_SB)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:126:2
	nrbd_nrsc_mvp nrbd_nrsc_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Start_SI(Start_S),
		.Kill_SI(Kill_SI),
		.Special_case_SBI(Special_case_SB),
		.Special_case_dly_SBI(Special_case_dly_SB),
		.Div_enable_SO(Div_enable_S),
		.Sqrt_enable_SO(Sqrt_enable_S),
		.Precision_ctl_SI(Precision_ctl_SI),
		.Format_sel_SI(Format_sel_SI),
		.Exp_a_DI(Exp_a_D),
		.Exp_b_DI(Exp_b_D),
		.Mant_a_DI(Mant_a_D),
		.Mant_b_DI(Mant_b_D),
		.Full_precision_SO(Full_precision_S),
		.FP32_SO(FP32_S),
		.FP64_SO(FP64_S),
		.FP16_SO(FP16_S),
		.FP16ALT_SO(FP16ALT_S),
		.Ready_SO(Ready_SO),
		.Done_SO(Done_SO),
		.Exp_z_DO(Exp_z_D),
		.Mant_z_DO(Mant_z_D)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/div_sqrt_top_mvp.sv:156:2
	norm_div_sqrt_mvp fpu_norm_U0(
		.Mant_in_DI(Mant_z_D),
		.Exp_in_DI(Exp_z_D),
		.Sign_in_DI(Sign_z_D),
		.Div_enable_SI(Div_enable_S),
		.Sqrt_enable_SI(Sqrt_enable_S),
		.Inf_a_SI(Inf_a_S),
		.Inf_b_SI(Inf_b_S),
		.Zero_a_SI(Zero_a_S),
		.Zero_b_SI(Zero_b_S),
		.NaN_a_SI(NaN_a_S),
		.NaN_b_SI(NaN_b_S),
		.SNaN_SI(SNaN_S),
		.RM_SI(RM_dly_S),
		.Full_precision_SI(Full_precision_S),
		.FP32_SI(FP32_S),
		.FP64_SI(FP64_S),
		.FP16_SI(FP16_S),
		.FP16ALT_SI(FP16ALT_S),
		.Result_DO(Result_DO),
		.Fflags_SO(Fflags_SO)
	);
endmodule
module iteration_div_sqrt_mvp (
	A_DI,
	B_DI,
	Div_enable_SI,
	Div_start_dly_SI,
	Sqrt_enable_SI,
	D_DI,
	D_DO,
	Sum_DO,
	Carry_out_DO
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:34:16
	parameter WIDTH = 25;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:38:4
	input wire [WIDTH - 1:0] A_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:39:4
	input wire [WIDTH - 1:0] B_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:40:4
	input wire Div_enable_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:41:4
	input wire Div_start_dly_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:42:4
	input wire Sqrt_enable_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:43:4
	input wire [1:0] D_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:45:4
	output wire [1:0] D_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:46:4
	output wire [WIDTH - 1:0] Sum_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:47:4
	output wire Carry_out_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:50:4
	wire D_carry_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:51:4
	wire Sqrt_cin_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:52:4
	wire Cin_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:54:4
	assign D_DO[0] = ~D_DI[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:55:4
	assign D_DO[1] = ~(D_DI[1] ^ D_DI[0]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:56:4
	assign D_carry_D = D_DI[1] | D_DI[0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:57:4
	assign Sqrt_cin_D = Sqrt_enable_SI && D_carry_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:58:4
	assign Cin_D = (Div_enable_SI ? 1'b0 : Sqrt_cin_D);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/iteration_div_sqrt_mvp.sv:59:4
	assign {Carry_out_DO, Sum_DO} = (A_DI + B_DI) + Cin_D;
endmodule
// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:44:1
// removed ["import defs_div_sqrt_mvp::*;"]
module norm_div_sqrt_mvp (
	Mant_in_DI,
	Exp_in_DI,
	Sign_in_DI,
	Div_enable_SI,
	Sqrt_enable_SI,
	Inf_a_SI,
	Inf_b_SI,
	Zero_a_SI,
	Zero_b_SI,
	NaN_a_SI,
	NaN_b_SI,
	SNaN_SI,
	RM_SI,
	Full_precision_SI,
	FP32_SI,
	FP64_SI,
	FP16_SI,
	FP16ALT_SI,
	Result_DO,
	Fflags_SO
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:48:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [56:0] Mant_in_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:49:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire signed [12:0] Exp_in_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:50:4
	input wire Sign_in_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:51:4
	input wire Div_enable_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:52:4
	input wire Sqrt_enable_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:53:4
	input wire Inf_a_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:54:4
	input wire Inf_b_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:55:4
	input wire Zero_a_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:56:4
	input wire Zero_b_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:57:4
	input wire NaN_a_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:58:4
	input wire NaN_b_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:59:4
	input wire SNaN_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:60:4
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:61:4
	input wire Full_precision_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:62:4
	input wire FP32_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:63:4
	input wire FP64_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:64:4
	input wire FP16_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:65:4
	input wire FP16ALT_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:67:4
	output reg [63:0] Result_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:68:4
	output wire [4:0] Fflags_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:72:4
	reg Sign_res_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:74:4
	reg NV_OP_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:75:4
	reg Exp_OF_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:76:4
	reg Exp_UF_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:77:4
	reg Div_Zero_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:78:4
	wire In_Exact_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:83:4
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_res_norm_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:84:4
	reg [10:0] Exp_res_norm_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:90:3
	wire [12:0] Exp_Max_RS_FP64_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:91:3
	localparam defs_div_sqrt_mvp_C_EXP_FP32 = 8;
	wire [9:0] Exp_Max_RS_FP32_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:92:3
	localparam defs_div_sqrt_mvp_C_EXP_FP16 = 5;
	wire [6:0] Exp_Max_RS_FP16_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:93:3
	localparam defs_div_sqrt_mvp_C_EXP_FP16ALT = 8;
	wire [9:0] Exp_Max_RS_FP16ALT_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:95:3
	assign Exp_Max_RS_FP64_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] + defs_div_sqrt_mvp_C_MANT_FP64) + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:96:3
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	assign Exp_Max_RS_FP32_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP32:0] + defs_div_sqrt_mvp_C_MANT_FP32) + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:97:3
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	assign Exp_Max_RS_FP16_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16:0] + defs_div_sqrt_mvp_C_MANT_FP16) + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:98:3
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	assign Exp_Max_RS_FP16ALT_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16ALT:0] + defs_div_sqrt_mvp_C_MANT_FP16ALT) + 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:99:3
	wire [12:0] Num_RS_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:100:3
	assign Num_RS_D = ~Exp_in_DI + 2;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:101:3
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_RS_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:102:3
	wire [56:0] Mant_forsticky_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:103:3
	assign {Mant_RS_D, Mant_forsticky_D} = {Mant_in_DI, {53 {1'b0}}} >> Num_RS_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:105:3
	wire [12:0] Exp_subOne_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:106:3
	assign Exp_subOne_D = Exp_in_DI - 1;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:109:4
	reg [1:0] Mant_lower_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:110:4
	reg Mant_sticky_bit_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:111:4
	reg [56:0] Mant_forround_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:113:4
	localparam defs_div_sqrt_mvp_C_EXP_ONE_FP64 = 13'h0001;
	localparam defs_div_sqrt_mvp_C_MANT_NAN_FP64 = 52'h8000000000000;
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:116:8
		if (NaN_a_SI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:118:12
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:119:12
			Exp_OF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:120:12
			Exp_UF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:121:12
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:122:12
			Exp_res_norm_D = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:123:12
			Mant_forround_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:124:12
			Sign_res_D = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:125:12
			NV_OP_S = SNaN_SI;
		end
		else if (NaN_b_SI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:130:11
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:131:11
			Exp_OF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:132:11
			Exp_UF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:133:11
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:134:11
			Exp_res_norm_D = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:135:11
			Mant_forround_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:136:11
			Sign_res_D = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:137:11
			NV_OP_S = SNaN_SI;
		end
		else if (Inf_a_SI) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:142:11
				if (Div_enable_SI && Inf_b_SI) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:144:15
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:145:15
					Exp_OF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:146:15
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:147:15
					Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:148:15
					Exp_res_norm_D = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:149:15
					Mant_forround_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:150:15
					Sign_res_D = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:151:15
					NV_OP_S = 1'b1;
				end
				else if (Sqrt_enable_SI && Sign_in_DI) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:154:13
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:155:13
					Exp_OF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:156:13
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:157:13
					Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:158:13
					Exp_res_norm_D = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:159:13
					Mant_forround_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:160:13
					Sign_res_D = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:161:13
					NV_OP_S = 1'b1;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:163:13
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:164:13
					Exp_OF_S = 1'b1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:165:13
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:166:13
					Mant_res_norm_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:167:13
					Exp_res_norm_D = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:168:13
					Mant_forround_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:169:13
					Sign_res_D = Sign_in_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:170:13
					NV_OP_S = 1'b0;
				end
			end
		end
		else if (Div_enable_SI && Inf_b_SI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:176:11
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:177:11
			Exp_OF_S = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:178:11
			Exp_UF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:179:11
			Mant_res_norm_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:180:11
			Exp_res_norm_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:181:11
			Mant_forround_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:182:11
			Sign_res_D = Sign_in_DI;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:183:11
			NV_OP_S = 1'b0;
		end
		else if (Zero_a_SI) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:188:10
				if (Div_enable_SI && Zero_b_SI) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:190:15
					Div_Zero_S = 1'b1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:191:15
					Exp_OF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:192:15
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:193:15
					Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:194:15
					Exp_res_norm_D = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:195:15
					Mant_forround_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:196:15
					Sign_res_D = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:197:15
					NV_OP_S = 1'b1;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:201:14
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:202:14
					Exp_OF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:203:14
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:204:14
					Mant_res_norm_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:205:14
					Exp_res_norm_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:206:14
					Mant_forround_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:207:14
					Sign_res_D = Sign_in_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:208:14
					NV_OP_S = 1'b0;
				end
			end
		end
		else if (Div_enable_SI && Zero_b_SI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:214:10
			Div_Zero_S = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:215:10
			Exp_OF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:216:10
			Exp_UF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:217:10
			Mant_res_norm_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:218:10
			Exp_res_norm_D = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:219:10
			Mant_forround_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:220:10
			Sign_res_D = Sign_in_DI;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:221:10
			NV_OP_S = 1'b0;
		end
		else if (Sign_in_DI && Sqrt_enable_SI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:226:11
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:227:11
			Exp_OF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:228:11
			Exp_UF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:229:11
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:230:11
			Exp_res_norm_D = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:231:11
			Mant_forround_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:232:11
			Sign_res_D = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:233:11
			NV_OP_S = 1'b1;
		end
		else if (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] == {12 {1'sb0}}) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:238:10
				if (Mant_in_DI != {57 {1'sb0}}) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:240:14
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:241:14
					Exp_OF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:242:14
					Exp_UF_S = 1'b1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:243:14
					Mant_res_norm_D = {1'b0, Mant_in_DI[56:5]};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:244:14
					Exp_res_norm_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:245:14
					Mant_forround_D = {Mant_in_DI[4:0], {defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:246:14
					Sign_res_D = Sign_in_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:247:14
					NV_OP_S = 1'b0;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:251:14
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:252:14
					Exp_OF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:253:14
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:254:14
					Mant_res_norm_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:255:14
					Exp_res_norm_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:256:14
					Mant_forround_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:257:14
					Sign_res_D = Sign_in_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:258:14
					NV_OP_S = 1'b0;
				end
			end
		end
		else if ((Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] == defs_div_sqrt_mvp_C_EXP_ONE_FP64) && ~Mant_in_DI[56]) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:264:11
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:265:11
			Exp_OF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:266:11
			Exp_UF_S = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:267:11
			Mant_res_norm_D = Mant_in_DI[56:4];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:268:11
			Exp_res_norm_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:269:11
			Mant_forround_D = {Mant_in_DI[3:0], {53 {1'b0}}};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:270:11
			Sign_res_D = Sign_in_DI;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:271:11
			NV_OP_S = 1'b0;
		end
		else if (Exp_in_DI[12]) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:276:11
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:277:11
			Exp_OF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:278:11
			Exp_UF_S = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:279:11
			Mant_res_norm_D = {Mant_RS_D[defs_div_sqrt_mvp_C_MANT_FP64:0]};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:280:11
			Exp_res_norm_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:281:11
			Mant_forround_D = {Mant_forsticky_D[56:0]};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:282:11
			Sign_res_D = Sign_in_DI;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:283:11
			NV_OP_S = 1'b0;
		end
		else if ((((Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP32] && FP32_SI) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64] && FP64_SI)) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16] && FP16_SI)) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16ALT] && FP16ALT_SI)) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:288:11
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:289:11
			Exp_OF_S = 1'b1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:290:11
			Exp_UF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:291:11
			Mant_res_norm_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:292:11
			Exp_res_norm_D = 1'sb1;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:293:11
			Mant_forround_D = 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:294:11
			Sign_res_D = Sign_in_DI;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:295:11
			NV_OP_S = 1'b0;
		end
		else if (((((Exp_in_DI[7:0] == {8 {1'sb1}}) && FP32_SI) | ((Exp_in_DI[10:0] == {11 {1'sb1}}) && FP64_SI)) | ((Exp_in_DI[4:0] == {5 {1'sb1}}) && FP16_SI)) | ((Exp_in_DI[7:0] == {8 {1'sb1}}) && FP16ALT_SI)) begin
			begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:300:11
				if (~Mant_in_DI[56]) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:302:15
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:303:15
					Exp_OF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:304:15
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:305:15
					Mant_res_norm_D = Mant_in_DI[55:3];
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:306:15
					Exp_res_norm_D = Exp_subOne_D;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:307:15
					Mant_forround_D = {Mant_in_DI[2:0], {54 {1'b0}}};
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:308:15
					Sign_res_D = Sign_in_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:309:15
					NV_OP_S = 1'b0;
				end
				else if (Mant_in_DI != {57 {1'sb0}}) begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:313:15
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:314:15
					Exp_OF_S = 1'b1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:315:15
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:316:15
					Mant_res_norm_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:317:15
					Exp_res_norm_D = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:318:15
					Mant_forround_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:319:15
					Sign_res_D = Sign_in_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:320:15
					NV_OP_S = 1'b0;
				end
				else begin
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:324:15
					Div_Zero_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:325:15
					Exp_OF_S = 1'b1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:326:15
					Exp_UF_S = 1'b0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:327:15
					Mant_res_norm_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:328:15
					Exp_res_norm_D = 1'sb1;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:329:15
					Mant_forround_D = 1'sb0;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:330:15
					Sign_res_D = Sign_in_DI;
					// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:331:15
					NV_OP_S = 1'b0;
				end
			end
		end
		else if (Mant_in_DI[56]) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:337:12
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:338:12
			Exp_OF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:339:12
			Exp_UF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:340:12
			Mant_res_norm_D = Mant_in_DI[56:4];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:341:12
			Exp_res_norm_D = Exp_in_DI[10:0];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:342:12
			Mant_forround_D = {Mant_in_DI[3:0], {53 {1'b0}}};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:343:12
			Sign_res_D = Sign_in_DI;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:344:12
			NV_OP_S = 1'b0;
		end
		else begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:349:12
			Div_Zero_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:350:12
			Exp_OF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:351:12
			Exp_UF_S = 1'b0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:352:12
			Mant_res_norm_D = Mant_in_DI[55:3];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:353:12
			Exp_res_norm_D = Exp_subOne_D;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:354:12
			Mant_forround_D = {Mant_in_DI[2:0], {54 {1'b0}}};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:355:12
			Sign_res_D = Sign_in_DI;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:356:12
			NV_OP_S = 1'b0;
		end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:365:4
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_upper_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:366:4
	wire [53:0] Mant_upperRounded_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:367:4
	reg Mant_roundUp_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:368:4
	wire Mant_rounded_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:370:3
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:372:7
		if (FP32_SI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:374:11
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:29], {29 {1'b0}}};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:375:11
			Mant_lower_D = Mant_res_norm_D[28:27];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:376:11
			Mant_sticky_bit_D = |Mant_res_norm_D[26:0];
		end
		else if (FP64_SI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:380:11
			Mant_upper_D = Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:0];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:381:11
			Mant_lower_D = Mant_forround_D[56:55];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:382:11
			Mant_sticky_bit_D = |Mant_forround_D[55:0];
		end
		else if (FP16_SI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:386:11
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:42], {42 {1'b0}}};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:387:11
			Mant_lower_D = Mant_res_norm_D[41:40];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:388:11
			Mant_sticky_bit_D = |Mant_res_norm_D[39:30];
		end
		else begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:392:11
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:45], {45 {1'b0}}};
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:393:11
			Mant_lower_D = Mant_res_norm_D[44:43];
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:394:11
			Mant_sticky_bit_D = |Mant_res_norm_D[42:30];
		end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:398:4
	assign Mant_rounded_S = |Mant_lower_D | Mant_sticky_bit_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:403:4
	localparam defs_div_sqrt_mvp_C_RM_MINUSINF = 3'h3;
	localparam defs_div_sqrt_mvp_C_RM_NEAREST = 3'h0;
	localparam defs_div_sqrt_mvp_C_RM_PLUSINF = 3'h2;
	localparam defs_div_sqrt_mvp_C_RM_TRUNC = 3'h1;
	always @(*) begin
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:405:9
		Mant_roundUp_S = 1'b0;
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:406:9
		case (RM_SI)
			defs_div_sqrt_mvp_C_RM_NEAREST:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:408:13
				Mant_roundUp_S = Mant_lower_D[1] && ((Mant_lower_D[0] | Mant_sticky_bit_D) | ((((FP32_SI && Mant_upper_D[29]) | (FP64_SI && Mant_upper_D[0])) | (FP16_SI && Mant_upper_D[42])) | (FP16ALT_SI && Mant_upper_D[45])));
			defs_div_sqrt_mvp_C_RM_TRUNC:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:410:13
				Mant_roundUp_S = 0;
			defs_div_sqrt_mvp_C_RM_PLUSINF:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:412:13
				Mant_roundUp_S = Mant_rounded_S & ~Sign_in_DI;
			defs_div_sqrt_mvp_C_RM_MINUSINF:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:414:13
				Mant_roundUp_S = Mant_rounded_S & Sign_in_DI;
			default:
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:416:13
				Mant_roundUp_S = 0;
		endcase
	end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:420:3
	wire Mant_renorm_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:421:3
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_roundUp_Vector_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:423:3
	assign Mant_roundUp_Vector_S = {7'h00, FP16ALT_SI && Mant_roundUp_S, 2'h0, FP16_SI && Mant_roundUp_S, 12'h000, FP32_SI && Mant_roundUp_S, 28'h0000000, FP64_SI && Mant_roundUp_S};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:426:3
	assign Mant_upperRounded_D = Mant_upper_D + Mant_roundUp_Vector_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:427:3
	assign Mant_renorm_S = Mant_upperRounded_D[53];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:432:3
	wire [51:0] Mant_res_round_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:433:3
	wire [10:0] Exp_res_round_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:436:3
	assign Mant_res_round_D = (Mant_renorm_S ? Mant_upperRounded_D[defs_div_sqrt_mvp_C_MANT_FP64:1] : Mant_upperRounded_D[51:0]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:437:3
	assign Exp_res_round_D = Exp_res_norm_D + Mant_renorm_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:442:3
	wire [51:0] Mant_before_format_ctl_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:443:3
	wire [10:0] Exp_before_format_ctl_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:444:3
	assign Mant_before_format_ctl_D = (Full_precision_SI ? Mant_res_round_D : Mant_res_norm_D);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:445:3
	assign Exp_before_format_ctl_D = (Full_precision_SI ? Exp_res_round_D : Exp_res_norm_D);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:447:3
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:449:7
		if (FP32_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:451:13
			Result_DO = {32'hffffffff, Sign_res_D, Exp_before_format_ctl_D[7:0], Mant_before_format_ctl_D[51:29]};
		else if (FP64_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:455:13
			Result_DO = {Sign_res_D, Exp_before_format_ctl_D[10:0], Mant_before_format_ctl_D[51:0]};
		else if (FP16_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:459:13
			Result_DO = {48'hffffffffffff, Sign_res_D, Exp_before_format_ctl_D[4:0], Mant_before_format_ctl_D[51:42]};
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:463:13
			Result_DO = {48'hffffffffffff, Sign_res_D, Exp_before_format_ctl_D[7:0], Mant_before_format_ctl_D[51:45]};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:467:1
	assign In_Exact_S = ~Full_precision_SI | Mant_rounded_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/norm_div_sqrt_mvp.sv:468:1
	assign Fflags_SO = {NV_OP_S, Div_Zero_S, Exp_OF_S, Exp_UF_S, In_Exact_S};
endmodule
// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:34:1
// removed ["import defs_div_sqrt_mvp::*;"]
module nrbd_nrsc_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Start_SI,
	Kill_SI,
	Special_case_SBI,
	Special_case_dly_SBI,
	Precision_ctl_SI,
	Format_sel_SI,
	Mant_a_DI,
	Mant_b_DI,
	Exp_a_DI,
	Exp_b_DI,
	Div_enable_SO,
	Sqrt_enable_SO,
	Full_precision_SO,
	FP32_SO,
	FP64_SO,
	FP16_SO,
	FP16ALT_SO,
	Ready_SO,
	Done_SO,
	Mant_z_DO,
	Exp_z_DO
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:39:4
	input wire Clk_CI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:40:4
	input wire Rst_RBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:41:4
	input wire Div_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:42:4
	input wire Sqrt_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:43:4
	input wire Start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:44:4
	input wire Kill_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:45:4
	input wire Special_case_SBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:46:4
	input wire Special_case_dly_SBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:47:4
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:48:4
	input wire [1:0] Format_sel_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:49:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:50:4
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:51:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:52:4
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:54:4
	output wire Div_enable_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:55:4
	output wire Sqrt_enable_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:57:4
	output wire Full_precision_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:58:4
	output wire FP32_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:59:4
	output wire FP64_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:60:4
	output wire FP16_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:61:4
	output wire FP16ALT_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:62:4
	output wire Ready_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:63:4
	output wire Done_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:64:4
	output wire [56:0] Mant_z_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:65:4
	output wire [12:0] Exp_z_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:69:5
	wire Div_start_dly_S;
	wire Sqrt_start_dly_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/nrbd_nrsc_mvp.sv:72:1
	control_mvp control_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Start_SI(Start_SI),
		.Kill_SI(Kill_SI),
		.Special_case_SBI(Special_case_SBI),
		.Special_case_dly_SBI(Special_case_dly_SBI),
		.Precision_ctl_SI(Precision_ctl_SI),
		.Format_sel_SI(Format_sel_SI),
		.Numerator_DI(Mant_a_DI),
		.Exp_num_DI(Exp_a_DI),
		.Denominator_DI(Mant_b_DI),
		.Exp_den_DI(Exp_b_DI),
		.Div_start_dly_SO(Div_start_dly_S),
		.Sqrt_start_dly_SO(Sqrt_start_dly_S),
		.Div_enable_SO(Div_enable_SO),
		.Sqrt_enable_SO(Sqrt_enable_SO),
		.Full_precision_SO(Full_precision_SO),
		.FP32_SO(FP32_SO),
		.FP64_SO(FP64_SO),
		.FP16_SO(FP16_SO),
		.FP16ALT_SO(FP16ALT_SO),
		.Ready_SO(Ready_SO),
		.Done_SO(Done_SO),
		.Mant_result_prenorm_DO(Mant_z_DO),
		.Exp_result_prenorm_DO(Exp_z_DO)
	);
endmodule
// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:35:1
// removed ["import defs_div_sqrt_mvp::*;"]
module preprocess_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Ready_SI,
	Operand_a_DI,
	Operand_b_DI,
	RM_SI,
	Format_sel_SI,
	Start_SO,
	Exp_a_DO_norm,
	Exp_b_DO_norm,
	Mant_a_DO_norm,
	Mant_b_DO_norm,
	RM_dly_SO,
	Sign_z_DO,
	Inf_a_SO,
	Inf_b_SO,
	Zero_a_SO,
	Zero_b_SO,
	NaN_a_SO,
	NaN_b_SO,
	SNaN_SO,
	Special_case_SBO,
	Special_case_dly_SBO
);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:39:4
	input wire Clk_CI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:40:4
	input wire Rst_RBI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:41:4
	input wire Div_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:42:4
	input wire Sqrt_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:43:4
	input wire Ready_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:45:4
	localparam defs_div_sqrt_mvp_C_OP_FP64 = 64;
	input wire [63:0] Operand_a_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:46:4
	input wire [63:0] Operand_b_DI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:47:4
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:48:4
	localparam defs_div_sqrt_mvp_C_FS = 2;
	input wire [1:0] Format_sel_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:51:4
	output wire Start_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:52:4
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	output wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_DO_norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:53:4
	output wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_DO_norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:54:4
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	output wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_DO_norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:55:4
	output wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_DO_norm;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:57:4
	output wire [2:0] RM_dly_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:59:4
	output wire Sign_z_DO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:60:4
	output wire Inf_a_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:61:4
	output wire Inf_b_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:62:4
	output wire Zero_a_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:63:4
	output wire Zero_b_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:64:4
	output wire NaN_a_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:65:4
	output wire NaN_b_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:66:4
	output wire SNaN_SO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:67:4
	output wire Special_case_SBO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:68:4
	output reg Special_case_dly_SBO;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:72:4
	wire Hb_a_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:73:4
	wire Hb_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:75:4
	reg [10:0] Exp_a_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:76:4
	reg [10:0] Exp_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:77:4
	reg [51:0] Mant_a_NonH_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:78:4
	reg [51:0] Mant_b_NonH_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:79:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:80:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:85:4
	reg Sign_a_D;
	reg Sign_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:86:4
	wire Start_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:88:6
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	localparam defs_div_sqrt_mvp_C_OP_FP16 = 16;
	localparam defs_div_sqrt_mvp_C_OP_FP16ALT = 16;
	localparam defs_div_sqrt_mvp_C_OP_FP32 = 32;
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:90:10
		case (Format_sel_SI)
			2'b00: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:93:16
				Sign_a_D = Operand_a_DI[31];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:94:16
				Sign_b_D = Operand_b_DI[31];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:95:16
				Exp_a_D = {3'h0, Operand_a_DI[30:defs_div_sqrt_mvp_C_MANT_FP32]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:96:16
				Exp_b_D = {3'h0, Operand_b_DI[30:defs_div_sqrt_mvp_C_MANT_FP32]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:97:16
				Mant_a_NonH_D = {Operand_a_DI[22:0], 29'h00000000};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:98:16
				Mant_b_NonH_D = {Operand_b_DI[22:0], 29'h00000000};
			end
			2'b01: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:102:16
				Sign_a_D = Operand_a_DI[63];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:103:16
				Sign_b_D = Operand_b_DI[63];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:104:16
				Exp_a_D = Operand_a_DI[62:defs_div_sqrt_mvp_C_MANT_FP64];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:105:16
				Exp_b_D = Operand_b_DI[62:defs_div_sqrt_mvp_C_MANT_FP64];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:106:16
				Mant_a_NonH_D = Operand_a_DI[51:0];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:107:16
				Mant_b_NonH_D = Operand_b_DI[51:0];
			end
			2'b10: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:111:16
				Sign_a_D = Operand_a_DI[15];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:112:16
				Sign_b_D = Operand_b_DI[15];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:113:16
				Exp_a_D = {6'h00, Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:114:16
				Exp_b_D = {6'h00, Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:115:16
				Mant_a_NonH_D = {Operand_a_DI[9:0], 42'h00000000000};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:116:16
				Mant_b_NonH_D = {Operand_b_DI[9:0], 42'h00000000000};
			end
			2'b11: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:120:16
				Sign_a_D = Operand_a_DI[15];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:121:16
				Sign_b_D = Operand_b_DI[15];
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:122:16
				Exp_a_D = {3'h0, Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:123:16
				Exp_b_D = {3'h0, Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT]};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:124:16
				Mant_a_NonH_D = {Operand_a_DI[6:0], 45'h000000000000};
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:125:16
				Mant_b_NonH_D = {Operand_b_DI[6:0], 45'h000000000000};
			end
		endcase
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:131:4
	assign Mant_a_D = {Hb_a_D, Mant_a_NonH_D};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:132:4
	assign Mant_b_D = {Hb_b_D, Mant_b_NonH_D};
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:134:4
	assign Hb_a_D = |Exp_a_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:135:4
	assign Hb_b_D = |Exp_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:137:4
	assign Start_S = Div_start_SI | Sqrt_start_SI;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:145:4
	reg Mant_a_prenorm_zero_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:146:4
	reg Mant_b_prenorm_zero_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:148:4
	wire Exp_a_prenorm_zero_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:149:4
	wire Exp_b_prenorm_zero_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:150:4
	assign Exp_a_prenorm_zero_S = ~Hb_a_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:151:4
	assign Exp_b_prenorm_zero_S = ~Hb_b_D;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:153:4
	reg Exp_a_prenorm_Inf_NaN_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:154:4
	reg Exp_b_prenorm_Inf_NaN_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:156:4
	wire Mant_a_prenorm_QNaN_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:157:4
	wire Mant_a_prenorm_SNaN_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:158:4
	wire Mant_b_prenorm_QNaN_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:159:4
	wire Mant_b_prenorm_SNaN_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:161:4
	assign Mant_a_prenorm_QNaN_S = Mant_a_NonH_D[51] && ~(|Mant_a_NonH_D[50:0]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:162:4
	assign Mant_a_prenorm_SNaN_S = ~Mant_a_NonH_D[51] && |Mant_a_NonH_D[50:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:163:4
	assign Mant_b_prenorm_QNaN_S = Mant_b_NonH_D[51] && ~(|Mant_b_NonH_D[50:0]);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:164:4
	assign Mant_b_prenorm_SNaN_S = ~Mant_b_NonH_D[51] && |Mant_b_NonH_D[50:0];
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:166:6
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP16 = 5'h1f;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP16ALT = 8'hff;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP32 = 8'hff;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP64 = 11'h7ff;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP16 = 10'h000;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT = 7'h00;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP32 = 23'h000000;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP64 = 52'h0000000000000;
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:168:10
		case (Format_sel_SI)
			2'b00: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:171:16
				Mant_a_prenorm_zero_S = Operand_a_DI[22:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP32;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:172:16
				Mant_b_prenorm_zero_S = Operand_b_DI[22:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP32;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:173:16
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[30:defs_div_sqrt_mvp_C_MANT_FP32] == defs_div_sqrt_mvp_C_EXP_INF_FP32;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:174:16
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[30:defs_div_sqrt_mvp_C_MANT_FP32] == defs_div_sqrt_mvp_C_EXP_INF_FP32;
			end
			2'b01: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:178:16
				Mant_a_prenorm_zero_S = Operand_a_DI[51:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP64;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:179:16
				Mant_b_prenorm_zero_S = Operand_b_DI[51:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP64;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:180:16
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[62:defs_div_sqrt_mvp_C_MANT_FP64] == defs_div_sqrt_mvp_C_EXP_INF_FP64;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:181:16
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[62:defs_div_sqrt_mvp_C_MANT_FP64] == defs_div_sqrt_mvp_C_EXP_INF_FP64;
			end
			2'b10: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:185:16
				Mant_a_prenorm_zero_S = Operand_a_DI[9:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:186:16
				Mant_b_prenorm_zero_S = Operand_b_DI[9:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:187:16
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16] == defs_div_sqrt_mvp_C_EXP_INF_FP16;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:188:16
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16] == defs_div_sqrt_mvp_C_EXP_INF_FP16;
			end
			2'b11: begin
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:192:16
				Mant_a_prenorm_zero_S = Operand_a_DI[6:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:193:16
				Mant_b_prenorm_zero_S = Operand_b_DI[6:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:194:16
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT] == defs_div_sqrt_mvp_C_EXP_INF_FP16ALT;
				// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:195:16
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT] == defs_div_sqrt_mvp_C_EXP_INF_FP16ALT;
			end
		endcase
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:203:4
	wire Zero_a_SN;
	reg Zero_a_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:204:4
	wire Zero_b_SN;
	reg Zero_b_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:205:4
	wire Inf_a_SN;
	reg Inf_a_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:206:4
	wire Inf_b_SN;
	reg Inf_b_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:207:4
	wire NaN_a_SN;
	reg NaN_a_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:208:4
	wire NaN_b_SN;
	reg NaN_b_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:209:4
	wire SNaN_SN;
	reg SNaN_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:211:4
	assign Zero_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_zero_S && Mant_a_prenorm_zero_S : Zero_a_SP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:212:4
	assign Zero_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_zero_S && Mant_b_prenorm_zero_S : Zero_b_SP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:213:4
	assign Inf_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_Inf_NaN_S && Mant_a_prenorm_zero_S : Inf_a_SP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:214:4
	assign Inf_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_Inf_NaN_S && Mant_b_prenorm_zero_S : Inf_b_SP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:215:4
	assign NaN_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_Inf_NaN_S && ~Mant_a_prenorm_zero_S : NaN_a_SP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:216:4
	assign NaN_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_Inf_NaN_S && ~Mant_b_prenorm_zero_S : NaN_b_SP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:217:4
	assign SNaN_SN = (Start_S && Ready_SI ? (Mant_a_prenorm_SNaN_S && NaN_a_SN) | (Mant_b_prenorm_SNaN_S && NaN_b_SN) : SNaN_SP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:219:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:221:9
		if (~Rst_RBI) begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:223:13
			Zero_a_SP <= 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:224:13
			Zero_b_SP <= 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:225:13
			Inf_a_SP <= 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:226:13
			Inf_b_SP <= 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:227:13
			NaN_a_SP <= 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:228:13
			NaN_b_SP <= 1'sb0;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:229:13
			SNaN_SP <= 1'sb0;
		end
		else begin
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:233:12
			Inf_a_SP <= Inf_a_SN;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:234:12
			Inf_b_SP <= Inf_b_SN;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:235:12
			Zero_a_SP <= Zero_a_SN;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:236:12
			Zero_b_SP <= Zero_b_SN;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:237:12
			NaN_a_SP <= NaN_a_SN;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:238:12
			NaN_b_SP <= NaN_b_SN;
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:239:12
			SNaN_SP <= SNaN_SN;
		end
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:247:4
	assign Special_case_SBO = ~{(Div_start_SI ? ((((Zero_a_SN | Zero_b_SN) | Inf_a_SN) | Inf_b_SN) | NaN_a_SN) | NaN_b_SN : ((Zero_a_SN | Inf_a_SN) | NaN_a_SN) | Sign_a_D)} && (Start_S && Ready_SI);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:250:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:252:8
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:254:13
			Special_case_dly_SBO <= 1'sb0;
		else if (Start_S && Ready_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:258:13
			Special_case_dly_SBO <= Special_case_SBO;
		else if (Special_case_dly_SBO)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:262:10
			Special_case_dly_SBO <= 1'b1;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:266:13
			Special_case_dly_SBO <= 1'sb0;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:274:4
	reg Sign_z_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:275:4
	reg Sign_z_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:277:4
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:279:8
		if (Div_start_SI && Ready_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:280:12
			Sign_z_DN = Sign_a_D ^ Sign_b_D;
		else if (Sqrt_start_SI && Ready_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:282:12
			Sign_z_DN = Sign_a_D;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:284:12
			Sign_z_DN = Sign_z_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:287:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:289:8
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:291:13
			Sign_z_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:295:13
			Sign_z_DP <= Sign_z_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:299:4
	reg [2:0] RM_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:300:4
	reg [2:0] RM_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:302:4
	always @(*)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:304:8
		if (Start_S && Ready_SI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:305:12
			RM_DN = RM_SI;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:307:12
			RM_DN = RM_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:310:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:312:8
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:314:13
			RM_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:318:13
			RM_DP <= RM_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:321:4
	assign RM_dly_SO = RM_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:323:4
	wire [5:0] Mant_leadingOne_a;
	wire [5:0] Mant_leadingOne_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:324:4
	wire Mant_zero_S_a;
	wire Mant_zero_S_b;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:326:3
	lzc #(
		.WIDTH(53),
		.MODE(1)
	) LOD_Ua(
		.in_i(Mant_a_D),
		.cnt_o(Mant_leadingOne_a),
		.empty_o(Mant_zero_S_a)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:335:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_norm_DN;
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_norm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:337:4
	assign Mant_a_norm_DN = (Start_S && Ready_SI ? Mant_a_D << Mant_leadingOne_a : Mant_a_norm_DP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:339:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:341:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:343:13
			Mant_a_norm_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:347:13
			Mant_a_norm_DP <= Mant_a_norm_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:351:4
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_norm_DN;
	reg [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_norm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:352:4
	assign Exp_a_norm_DN = (Start_S && Ready_SI ? (Exp_a_D - Mant_leadingOne_a) + |Mant_leadingOne_a : Exp_a_norm_DP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:354:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:356:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:358:13
			Exp_a_norm_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:362:13
			Exp_a_norm_DP <= Exp_a_norm_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:366:3
	lzc #(
		.WIDTH(53),
		.MODE(1)
	) LOD_Ub(
		.in_i(Mant_b_D),
		.cnt_o(Mant_leadingOne_b),
		.empty_o(Mant_zero_S_b)
	);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:376:4
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_norm_DN;
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_norm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:378:4
	assign Mant_b_norm_DN = (Start_S && Ready_SI ? Mant_b_D << Mant_leadingOne_b : Mant_b_norm_DP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:380:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:382:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:384:13
			Mant_b_norm_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:388:13
			Mant_b_norm_DP <= Mant_b_norm_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:392:4
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_norm_DN;
	reg [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_norm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:393:4
	assign Exp_b_norm_DN = (Start_S && Ready_SI ? (Exp_b_D - Mant_leadingOne_b) + |Mant_leadingOne_b : Exp_b_norm_DP);
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:395:4
	always @(posedge Clk_CI or negedge Rst_RBI)
		// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:397:9
		if (~Rst_RBI)
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:399:13
			Exp_b_norm_DP <= 1'sb0;
		else
			// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:403:13
			Exp_b_norm_DP <= Exp_b_norm_DN;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:411:4
	assign Start_SO = Start_S;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:412:4
	assign Exp_a_DO_norm = Exp_a_norm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:413:4
	assign Exp_b_DO_norm = Exp_b_norm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:414:4
	assign Mant_a_DO_norm = Mant_a_norm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:415:4
	assign Mant_b_DO_norm = Mant_b_norm_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:416:4
	assign Sign_z_DO = Sign_z_DP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:417:4
	assign Inf_a_SO = Inf_a_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:418:4
	assign Inf_b_SO = Inf_b_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:419:4
	assign Zero_a_SO = Zero_a_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:420:4
	assign Zero_b_SO = Zero_b_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:421:4
	assign NaN_a_SO = NaN_a_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:422:4
	assign NaN_b_SO = NaN_b_SP;
	// Trace: ../../rtl/../../third_party/fpnew/src/fpu_div_sqrt_mvp/hdl/preprocess_mvp.sv:423:4
	assign SNaN_SO = SNaN_SP;
endmodule
