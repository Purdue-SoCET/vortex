/*
    socet115 / zlagpaca@purdue.edu
    Zach Lagpacan

    module for faking memory with basic register file which can interface with Vortex memory interface
*/

`include "VX_define.vh"

module ram_fake_reg_file #(
    parameter WORD_W = 32;
)(
    // seq
    input clk, reset,

    // Memory Request:
    // vortex outputs
    input logic                             mem_req_valid;
    input logic                             mem_req_rw;
    input logic [`VX_MEM_BYTEEN_WIDTH-1:0]  mem_req_byteen;    
    input logic [`VX_MEM_ADDR_WIDTH-1:0]    mem_req_addr;
    input logic [`VX_MEM_DATA_WIDTH-1:0]    mem_req_data;
    input logic [`VX_MEM_TAG_WIDTH-1:0]     mem_req_tag;
    // vortex inputs
    output logic                            mem_req_ready;

    // Memory response:
    // vortex inputs
    output logic                            mem_rsp_valid;        
    output logic [`VX_MEM_DATA_WIDTH-1:0]   mem_rsp_data;
    output logic [`VX_MEM_TAG_WIDTH-1:0]    mem_rsp_tag;
    // vortex outputs
    input logic                             mem_rsp_ready;

    // Status:
    // vortex outputs
    input logic                             busy;

    // tb:
    output logic                            tb_addr_out_of_bounds;  
);
    // register file instances
    
    // chunk 0
    logic wen_0_80000000;
    logic [9-1:0] wsel_0_80000000;
    logic [32-1:0] wdata_0_80000000;
    logic [9-1:0] rsel_0_80000000;
    logic [32-1:0] rdata_0_80000000;
    
    reg_file #(
        .WORD_W (32),
        .NUM_WORDS (512),
        .SEL_W (9),
        .RESET_WORDS ({
            32'h6F008004, 32'h732F2034, 32'h930F8000, 32'h6308FF03, 32'h930F9000, 32'h6304FF03, 32'h930FB000, 32'h6300FF03, 32'h130F0000, 32'h63040F00, 32'h67000F00, 32'h732F2034, 32'h63540F00, 32'h6F004000, 32'h93E19153, 32'h171F0000, 32'h23223FFC, 32'h6FF09FFF, 32'h93000000, 32'h13010000, 32'h93010000, 32'h13020000, 32'h93020000, 32'h13030000, 32'h93030000, 32'h13040000, 32'h93040000, 32'h13050000, 32'h93050000, 32'h13060000, 32'h93060000, 32'h13070000, 32'h93070000, 32'h13080000, 32'h93080000, 32'h13090000, 32'h93090000, 32'h130A0000, 32'h930A0000, 32'h130B0000, 32'h930B0000, 32'h130C0000, 32'h930C0000, 32'h130D0000, 32'h930D0000, 32'h130E0000, 32'h930E0000, 32'h130F0000, 32'h930F0000, 32'h732540F1, 32'h63100500, 32'h97020000, 32'h93820201, 32'h73905230, 32'h73500018, 32'h97020000, 32'h93820202, 32'h73905230, 32'hB7020080, 32'h9382F2FF, 32'h7390023B, 32'h9302F001, 32'h7390023A, 32'h73504030, 32'h97020000, 32'h93824201, 32'h73905230, 32'h73502030, 32'h73503030, 32'h93010000, 32'h97020000, 32'h9382C2EE, 32'h73905230, 32'h13051000, 32'h1315F501, 32'h634C0500, 32'h0F00F00F, 32'h93011000, 32'h9308D005, 32'h13050000, 32'h73000000, 32'h93020000, 32'h638A0200, 32'h73905210, 32'hB7B20000, 32'h93829210, 32'h73902230, 32'h73500030, 32'h37250000, 32'h73200530, 32'h73503000, 32'h97020000, 32'h93824201, 32'h73901234, 32'h732540F1, 32'h73002030, 32'h93012000, 32'h17250000, 32'h1305C5E7, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD3711002, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13060000, 32'h631AD526, 32'h63187326, 32'h6396C526, 32'h93013000, 32'h17250000, 32'h130585E5, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD3711002, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13061000, 32'h6318D522, 32'h63167322, 32'h6394C522, 32'h93014000, 32'h17250000, 32'h130545E3, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD3711002, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13061000, 32'h6316D51E, 32'h6314731E, 32'h6392C51E, 32'h93015000, 32'h17250000, 32'h130505E1, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD371100A, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13060000, 32'h6314D51A, 32'h6312731A, 32'h6390C51A, 32'h93016000, 32'h17250000, 32'h1305C5DE, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD371100A, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13061000, 32'h6312D516, 32'h63107316, 32'h639EC514, 32'h93017000, 32'h17250000, 32'h130585DC, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD371100A, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13061000, 32'h6310D512, 32'h631E7310, 32'h639CC510, 32'h93018000, 32'h17250000, 32'h130545DA, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD3711012, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13060000, 32'h631ED50C, 32'h631C730C, 32'h639AC50C, 32'h93019000, 32'h17250000, 32'h130505D8, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD3711012, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13061000, 32'h631CD508, 32'h631A7308, 32'h6398C508, 32'h9301A000, 32'h17250000, 32'h1305C5D5, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD3711012, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13061000, 32'h631AD504, 32'h63187304, 32'h6396C504, 32'h9301B000, 32'h17250000, 32'h130585D3, 32'h07300500, 32'h87308500, 32'h07310501, 32'h83268501, 32'h0323C501, 32'hD371100A, 32'h27303500, 32'h83234500, 32'h03250500, 32'hF3151000, 32'h13060001, 32'h6318D500, 32'h63167300, 32'h6394C500, 32'h63103002, 32'h0F00F00F, 32'h63800100, 32'h93911100, 32'h93E11100, 32'h9308D005, 32'h13850100, 32'h73000000, 32'h0F00F00F, 32'h93011000, 32'h9308D005, 32'h13050000, 32'h73000000, 32'h731000C0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000
        })
    ) reg_file_0_80000000 (
        .clk (clk), .reset (reset),
        .wen (wen_0_80000000),
        .wsel (wsel_0_80000000),
        .wdata (wdata_0_80000000),
        .rsel (rsel_0_80000000),
        .rdata (rdata_0_80000000)
    );
    
    // chunk 1
    logic wen_1_80001000;
    logic [5-1:0] wsel_1_80001000;
    logic [32-1:0] wdata_1_80001000;
    logic [5-1:0] rsel_1_80001000;
    logic [32-1:0] rdata_1_80001000;
    
    reg_file #(
        .WORD_W (32),
        .NUM_WORDS (32),
        .SEL_W (5),
        .RESET_WORDS ({
            32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000
        })
    ) reg_file_1_80001000 (
        .clk (clk), .reset (reset),
        .wen (wen_1_80001000),
        .wsel (wsel_1_80001000),
        .wdata (wdata_1_80001000),
        .rsel (rsel_1_80001000),
        .rdata (rdata_1_80001000)
    );
    
    // chunk 2
    logic wen_2_80002000;
    logic [7-1:0] wsel_2_80002000;
    logic [32-1:0] wdata_2_80002000;
    logic [7-1:0] rsel_2_80002000;
    logic [32-1:0] rdata_2_80002000;
    
    reg_file #(
        .WORD_W (32),
        .NUM_WORDS (128),
        .SEL_W (7),
        .RESET_WORDS ({
            32'h00000000, 32'h00000440, 32'h00000000, 32'h0000F03F, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000C40, 32'h66666666, 32'h664C93C0, 32'h9A999999, 32'h9999F13F, 32'h00000000, 32'h00000000, 32'h00000000, 32'h004893C0, 32'hF1D4C853, 32'hFB210940, 32'h3A8C30E2, 32'h8E79453E, 32'h00000000, 32'h00000000, 32'hDF6D2055, 32'hFB210940, 32'h00000000, 32'h00000440, 32'h00000000, 32'h0000F03F, 32'h00000000, 32'h00000000, 32'h00000000, 32'h0000F83F, 32'h66666666, 32'h664C93C0, 32'h9A999999, 32'h9999F1BF, 32'h00000000, 32'h00000000, 32'h00000000, 32'h004893C0, 32'hF1D4C853, 32'hFB210940, 32'h3A8C30E2, 32'h8E79453E, 32'h00000000, 32'h00000000, 32'h033C7152, 32'hFB210940, 32'h00000000, 32'h00000440, 32'h00000000, 32'h0000F03F, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000440, 32'h66666666, 32'h664C93C0, 32'h9A999999, 32'h9999F1BF, 32'h00000000, 32'h00000000, 32'h3D0AD7A3, 32'h703A9540, 32'hF1D4C853, 32'hFB210940, 32'h3A8C30E2, 32'h8E79453E, 32'h00000000, 32'h00000000, 32'h09FFC1A5, 32'hC5DD603E, 32'h00000000, 32'h0000F07F, 32'h00000000, 32'h0000F07F, 32'h00000000, 32'h00000000, 32'h00000000, 32'h0000F87F, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000
        })
    ) reg_file_2_80002000 (
        .clk (clk), .reset (reset),
        .wen (wen_2_80002000),
        .wsel (wsel_2_80002000),
        .wdata (wdata_2_80002000),
        .rsel (rsel_2_80002000),
        .rdata (rdata_2_80002000)
    );
    
    // need reg file/chunk selection signal
    logic [2-1:0] chunk_sel;

    // addr hashing logic
    always_comb begin : ADDR_HASHING_LOGIC
        // bit = 1 branch
        if (mem_req_addr[18] == 1'b1)
        begin
            chunk_sel = 2
        end
        // bit = 0 branch
        else if (mem_req_addr[18] == 1'b0)
        begin
            if (mem_req_addr[19] == 1'b0)
            begin
                chunk_sel = 0
            end
            else if (mem_req_addr[19] == 1'b1)
            begin
                chunk_sel = 1
            end
        end
        else
        begin
            $display("error: got to else in high-level branch")
        end
        
        // hardwired outputs:
        // hardwiring for chunk 0
        wsel_0_80000000 = mem_req_addr[9-1:0];
        wdata_0_80000000 = mem_req_data[9-1:0];
        rsel_0_80000000 = mem_req_addr[9-1:0];
        // hardwiring for chunk 1
        wsel_1_80001000 = mem_req_addr[5-1:0];
        wdata_1_80001000 = mem_req_data[5-1:0];
        rsel_1_80001000 = mem_req_addr[5-1:0];
        // hardwiring for chunk 2
        wsel_2_80002000 = mem_req_addr[7-1:0];
        wdata_2_80002000 = mem_req_data[7-1:0];
        rsel_2_80002000 = mem_req_addr[7-1:0];
        
        // default outputs:
        mem_rsp_data = '0;
        tb_addr_out_of_bounds = 1'b0;        // chunk wen's:
        wen_0_80000000 = 1'b0;
        wen_1_80001000 = 1'b0;
        wen_2_80002000 = 1'b0;
        
        // case for routing to diff reg file chunks
        casez (chunk_sel)
        
            // select chunk 0
            0:
            begin
                // write routing
                wen_0_80000000 = mem_req_rw;
        
                // read routing
                mem_rsp_data = rdata_0_80000000;
            end
        
            // select chunk 1
            1:
            begin
                // write routing
                wen_1_80001000 = mem_req_rw;
        
                // read routing
                mem_rsp_data = rdata_1_80001000;
            end
        
            // select chunk 2
            2:
            begin
                // write routing
                wen_2_80002000 = mem_req_rw;
        
                // read routing
                mem_rsp_data = rdata_2_80002000;
            end
        
            // shouldn't get here
            default:
            begin
                mem_rsp_data = '0;
                tb_addr_out_of_bounds = 1'b1;
            end
        endcase
    end

    // other combinational logic for memory interface
    always_comb begin : OTHER_MEM_COMB_LOGIC

        mem_req_ready = 1'b1; // when read or write ready (always)
        mem_rsp_valid = 1'b1; // when read ready (always)
        mem_rsp_tag = mem_req_tag; // match req immediately
    end

    // NOTES:
    // don't know what to do with: 
        // mem_req_byteeen
        // busy

endmodule
