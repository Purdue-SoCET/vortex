/*
    socet115 / zlagpaca@purdue.edu
    Zach Lagpacan

    module for on-chip RAM fake register file with AFTx07 AHB slave interface and Vortex memory interface 
*/

// temporary include to have defined vals
// `include "local_mem.vh"
`include "../include/VX_define.vh"
// `include "VX_define.vh"

// size of register file (128 Kb -> 16 KB -> 16*2^10 B -> 2^14 B -> 0x4000 B worth of byte address space)
`define REG_FILE_BYTE_WIDTH = 14
`define REG_FILE_BYTE_SIZE = 2**REG_FILE_BYTE_WIDTH

//////////////////////////////////
// Generic Bus Interface (AHB): //
//////////////////////////////////

`ifndef GENERIC_BUS_IF_VH
`define GENERIC_BUS_IF_VH

typedef logic [WORD_SIZE-1:0] word_t;

interface generic_bus_if ();
    // import rv32i_types_pkg::*;

    // logic [RAM_ADDR_SIZE-1:0] addr;
    logic [32-1:0] addr;                // RAM_ADDR_SIZE = 32
    word_t wdata;
    word_t rdata;
    logic ren,wen;
    logic busy;
    logic [3:0] byte_en;

    modport generic_bus (
        input addr, ren, wen, wdata, byte_en,
        output rdata, busy
    );

    modport cpu (
        input rdata, busy,
        output addr, ren, wen, wdata, byte_en
    );

endinterface

`endif //GENERIC_BUS_IF_VH

module Vortex_mem_slave #(
)(
    /////////////////
    // Sequential: //
    /////////////////
    input clk, reset,

    ///////////////////////
    // Memory Interface: //
    ///////////////////////

    // Memory Request:
    // vortex outputs
    input logic                             mem_req_valid,
    input logic                             mem_req_rw,
    input logic [`VX_MEM_BYTEEN_WIDTH-1:0]  mem_req_byteen, // 64 (512 / 8)
    input logic [`VX_MEM_ADDR_WIDTH-1:0]    mem_req_addr,   // 26
    input logic [`VX_MEM_DATA_WIDTH-1:0]    mem_req_data,   // 512
    input logic [`VX_MEM_TAG_WIDTH-1:0]     mem_req_tag,    // 56 (55 for SM disabled)
    // vortex inputs
    output logic                            mem_req_ready,

    // Memory response:
    // vortex inputs
    output logic                            mem_rsp_valid,        
    output logic [`VX_MEM_DATA_WIDTH-1:0]   mem_rsp_data,   // 512
    output logic [`VX_MEM_TAG_WIDTH-1:0]    mem_rsp_tag,    // 56 (55 for SM disabled)
    // vortex outputs
    input logic                             mem_rsp_ready,

    // Status:
    // vortex outputs
    input logic                             busy,

    // tb:
    output logic                            tb_addr_out_of_bounds,

    //////////////////////////////////
    // Generic Bus Interface (AHB): //
    //////////////////////////////////

    generic_bus_if.generic_bus              gbif
);
    // internal signals:
    // reg file signals (bytewise)
    logic [7:0] reg_file        [REG_FILE_BYTE_SIZE-1:0];
    logic [7:0] next_reg_file   [REG_FILE_BYTE_SIZE-1:0];

    // reg file instance
    always_ff @ (posedge clk) begin : REG_FILE_FF_LOGIC
        if (reset)
        begin
            reg_file[0] <= 8'h73
            reg_file[1] <= 8'h25
            reg_file[2] <= 8'h10
            reg_file[3] <= 8'hFC
            reg_file[4] <= 8'h97
            reg_file[5] <= 8'h05
            reg_file[6] <= 8'h00
            reg_file[7] <= 8'h00
            reg_file[8] <= 8'h93
            reg_file[9] <= 8'h85
            reg_file[10] <= 8'hC5
            reg_file[11] <= 8'h09
            reg_file[12] <= 8'h6B
            reg_file[13] <= 8'h10
            reg_file[14] <= 8'hB5
            reg_file[15] <= 8'h00
            reg_file[16] <= 8'hEF
            reg_file[17] <= 8'h00
            reg_file[18] <= 8'h00
            reg_file[19] <= 8'h09
            reg_file[20] <= 8'h13
            reg_file[21] <= 8'h05
            reg_file[22] <= 8'h10
            reg_file[23] <= 8'h00
            reg_file[24] <= 8'h6B
            reg_file[25] <= 8'h00
            reg_file[26] <= 8'h05
            reg_file[27] <= 8'h00
            reg_file[28] <= 8'h73
            reg_file[29] <= 8'h25
            reg_file[30] <= 8'h10
            reg_file[31] <= 8'hFC
            reg_file[32] <= 8'h97
            reg_file[33] <= 8'h05
            reg_file[34] <= 8'h00
            reg_file[35] <= 8'h00
            reg_file[36] <= 8'h93
            reg_file[37] <= 8'h85
            reg_file[38] <= 8'h05
            reg_file[39] <= 8'h12
            reg_file[40] <= 8'h6B
            reg_file[41] <= 8'h10
            reg_file[42] <= 8'hB5
            reg_file[43] <= 8'h00
            reg_file[44] <= 8'hEF
            reg_file[45] <= 8'h00
            reg_file[46] <= 8'h40
            reg_file[47] <= 8'h11
            reg_file[48] <= 8'h13
            reg_file[49] <= 8'h05
            reg_file[50] <= 8'h10
            reg_file[51] <= 8'h00
            reg_file[52] <= 8'h6B
            reg_file[53] <= 8'h00
            reg_file[54] <= 8'h05
            reg_file[55] <= 8'h00
            reg_file[56] <= 8'h17
            reg_file[57] <= 8'h15
            reg_file[58] <= 8'h00
            reg_file[59] <= 8'h00
            reg_file[60] <= 8'h13
            reg_file[61] <= 8'h05
            reg_file[62] <= 8'h85
            reg_file[63] <= 8'h40
            reg_file[64] <= 8'h17
            reg_file[65] <= 8'h16
            reg_file[66] <= 8'h00
            reg_file[67] <= 8'h00
            reg_file[68] <= 8'h13
            reg_file[69] <= 8'h06
            reg_file[70] <= 8'h06
            reg_file[71] <= 8'h48
            reg_file[72] <= 8'h33
            reg_file[73] <= 8'h06
            reg_file[74] <= 8'hA6
            reg_file[75] <= 8'h40
            reg_file[76] <= 8'h93
            reg_file[77] <= 8'h05
            reg_file[78] <= 8'h00
            reg_file[79] <= 8'h00
            reg_file[80] <= 8'hEF
            reg_file[81] <= 8'h00
            reg_file[82] <= 8'hD0
            reg_file[83] <= 8'h29
            reg_file[84] <= 8'h17
            reg_file[85] <= 8'h05
            reg_file[86] <= 8'h00
            reg_file[87] <= 8'h00
            reg_file[88] <= 8'h13
            reg_file[89] <= 8'h05
            reg_file[90] <= 8'hC5
            reg_file[91] <= 8'h1D
            reg_file[92] <= 8'hEF
            reg_file[93] <= 8'h00
            reg_file[94] <= 8'hD0
            reg_file[95] <= 8'h12
            reg_file[96] <= 8'hEF
            reg_file[97] <= 8'h00
            reg_file[98] <= 8'hC0
            reg_file[99] <= 8'h13
            reg_file[100] <= 8'hEF
            reg_file[101] <= 8'h00
            reg_file[102] <= 8'h80
            reg_file[103] <= 8'h00
            reg_file[104] <= 8'h6F
            reg_file[105] <= 8'h00
            reg_file[106] <= 8'h50
            reg_file[107] <= 8'h13
            reg_file[108] <= 8'h93
            reg_file[109] <= 8'h07
            reg_file[110] <= 8'hF0
            reg_file[111] <= 8'hFF
            reg_file[112] <= 8'h6B
            reg_file[113] <= 8'h80
            reg_file[114] <= 8'h07
            reg_file[115] <= 8'h00
            reg_file[116] <= 8'h13
            reg_file[117] <= 8'h05
            reg_file[118] <= 8'h00
            reg_file[119] <= 8'h00
            reg_file[120] <= 8'h67
            reg_file[121] <= 8'h80
            reg_file[122] <= 8'h00
            reg_file[123] <= 8'h00
            reg_file[124] <= 8'h93
            reg_file[125] <= 8'h07
            reg_file[126] <= 8'h00
            reg_file[127] <= 8'h00
            reg_file[128] <= 8'h63
            reg_file[129] <= 8'h88
            reg_file[130] <= 8'h07
            reg_file[131] <= 8'h00
            reg_file[132] <= 8'h37
            reg_file[133] <= 8'h05
            reg_file[134] <= 8'h00
            reg_file[135] <= 8'h80
            reg_file[136] <= 8'h13
            reg_file[137] <= 8'h05
            reg_file[138] <= 8'h05
            reg_file[139] <= 8'h23
            reg_file[140] <= 8'h6F
            reg_file[141] <= 8'h00
            reg_file[142] <= 8'hD0
            reg_file[143] <= 8'h0F
            reg_file[144] <= 8'h67
            reg_file[145] <= 8'h80
            reg_file[146] <= 8'h00
            reg_file[147] <= 8'h00
            reg_file[148] <= 8'h93
            reg_file[149] <= 8'h01
            reg_file[150] <= 8'h04
            reg_file[151] <= 8'h00
            reg_file[152] <= 8'h13
            reg_file[153] <= 8'h05
            reg_file[154] <= 8'h00
            reg_file[155] <= 8'h00
            reg_file[156] <= 8'h6B
            reg_file[157] <= 8'h00
            reg_file[158] <= 8'h05
            reg_file[159] <= 8'h00
            reg_file[160] <= 8'h13
            reg_file[161] <= 8'h05
            reg_file[162] <= 8'hF0
            reg_file[163] <= 8'hFF
            reg_file[164] <= 8'h6B
            reg_file[165] <= 8'h00
            reg_file[166] <= 8'h05
            reg_file[167] <= 8'h00
            reg_file[168] <= 8'h97
            reg_file[169] <= 8'h11
            reg_file[170] <= 8'h00
            reg_file[171] <= 8'h00
            reg_file[172] <= 8'h93
            reg_file[173] <= 8'h81
            reg_file[174] <= 8'h01
            reg_file[175] <= 8'h76
            reg_file[176] <= 8'h37
            reg_file[177] <= 8'h01
            reg_file[178] <= 8'h00
            reg_file[179] <= 8'hFF
            reg_file[180] <= 8'h73
            reg_file[181] <= 8'h25
            reg_file[182] <= 8'h10
            reg_file[183] <= 8'hCC
            reg_file[184] <= 8'h93
            reg_file[185] <= 8'h15
            reg_file[186] <= 8'hA5
            reg_file[187] <= 8'h00
            reg_file[188] <= 8'h33
            reg_file[189] <= 8'h01
            reg_file[190] <= 8'hB1
            reg_file[191] <= 8'h40
            reg_file[192] <= 8'h93
            reg_file[193] <= 8'h05
            reg_file[194] <= 8'h00
            reg_file[195] <= 8'h00
            reg_file[196] <= 8'h33
            reg_file[197] <= 8'h05
            reg_file[198] <= 8'hB5
            reg_file[199] <= 8'h02
            reg_file[200] <= 8'h17
            reg_file[201] <= 8'h12
            reg_file[202] <= 8'h00
            reg_file[203] <= 8'h00
            reg_file[204] <= 8'h13
            reg_file[205] <= 8'h02
            reg_file[206] <= 8'h72
            reg_file[207] <= 8'h43
            reg_file[208] <= 8'h33
            reg_file[209] <= 8'h02
            reg_file[210] <= 8'hA2
            reg_file[211] <= 8'h00
            reg_file[212] <= 8'h13
            reg_file[213] <= 8'h72
            reg_file[214] <= 8'h02
            reg_file[215] <= 8'hFC
            reg_file[216] <= 8'hF3
            reg_file[217] <= 8'h26
            reg_file[218] <= 8'h30
            reg_file[219] <= 8'hCC
            reg_file[220] <= 8'h63
            reg_file[221] <= 8'h86
            reg_file[222] <= 8'h06
            reg_file[223] <= 8'h00
            reg_file[224] <= 8'h13
            reg_file[225] <= 8'h05
            reg_file[226] <= 8'h00
            reg_file[227] <= 8'h00
            reg_file[228] <= 8'h6B
            reg_file[229] <= 8'h00
            reg_file[230] <= 8'h05
            reg_file[231] <= 8'h00
            reg_file[232] <= 8'h67
            reg_file[233] <= 8'h80
            reg_file[234] <= 8'h00
            reg_file[235] <= 8'h00
            reg_file[236] <= 8'h13
            reg_file[237] <= 8'h05
            reg_file[238] <= 8'hF0
            reg_file[239] <= 8'hFF
            reg_file[240] <= 8'h67
            reg_file[241] <= 8'h80
            reg_file[242] <= 8'h00
            reg_file[243] <= 8'h00
            reg_file[244] <= 8'h13
            reg_file[245] <= 8'h05
            reg_file[246] <= 8'hF0
            reg_file[247] <= 8'hFF
            reg_file[248] <= 8'h67
            reg_file[249] <= 8'h80
            reg_file[250] <= 8'h00
            reg_file[251] <= 8'h00
            reg_file[252] <= 8'h13
            reg_file[253] <= 8'h05
            reg_file[254] <= 8'h00
            reg_file[255] <= 8'h00
            reg_file[256] <= 8'h67
            reg_file[257] <= 8'h80
            reg_file[258] <= 8'h00
            reg_file[259] <= 8'h00
            reg_file[260] <= 8'h13
            reg_file[261] <= 8'h05
            reg_file[262] <= 8'h00
            reg_file[263] <= 8'h00
            reg_file[264] <= 8'h67
            reg_file[265] <= 8'h80
            reg_file[266] <= 8'h00
            reg_file[267] <= 8'h00
            reg_file[268] <= 8'h13
            reg_file[269] <= 8'h05
            reg_file[270] <= 8'hF0
            reg_file[271] <= 8'hFF
            reg_file[272] <= 8'h67
            reg_file[273] <= 8'h80
            reg_file[274] <= 8'h00
            reg_file[275] <= 8'h00
            reg_file[276] <= 8'h13
            reg_file[277] <= 8'h05
            reg_file[278] <= 8'hF0
            reg_file[279] <= 8'hFF
            reg_file[280] <= 8'h67
            reg_file[281] <= 8'h80
            reg_file[282] <= 8'h00
            reg_file[283] <= 8'h00
            reg_file[284] <= 8'h73
            reg_file[285] <= 8'h00
            reg_file[286] <= 8'h10
            reg_file[287] <= 8'h00
            reg_file[288] <= 8'h13
            reg_file[289] <= 8'h05
            reg_file[290] <= 8'h00
            reg_file[291] <= 8'h00
            reg_file[292] <= 8'h67
            reg_file[293] <= 8'h80
            reg_file[294] <= 8'h00
            reg_file[295] <= 8'h00
            reg_file[296] <= 8'h13
            reg_file[297] <= 8'h05
            reg_file[298] <= 8'h06
            reg_file[299] <= 8'h00
            reg_file[300] <= 8'h67
            reg_file[301] <= 8'h80
            reg_file[302] <= 8'h00
            reg_file[303] <= 8'h00
            reg_file[304] <= 8'h13
            reg_file[305] <= 8'h05
            reg_file[306] <= 8'hF0
            reg_file[307] <= 8'hFF
            reg_file[308] <= 8'h67
            reg_file[309] <= 8'h80
            reg_file[310] <= 8'h00
            reg_file[311] <= 8'h00
            reg_file[312] <= 8'h73
            reg_file[313] <= 8'h25
            reg_file[314] <= 8'h40
            reg_file[315] <= 8'hF1
            reg_file[316] <= 8'h67
            reg_file[317] <= 8'h80
            reg_file[318] <= 8'h00
            reg_file[319] <= 8'h00
            reg_file[320] <= 8'h13
            reg_file[321] <= 8'h01
            reg_file[322] <= 8'h01
            reg_file[323] <= 8'hFF
            reg_file[324] <= 8'h23
            reg_file[325] <= 8'h26
            reg_file[326] <= 8'h11
            reg_file[327] <= 8'h00
            reg_file[328] <= 8'h23
            reg_file[329] <= 8'h24
            reg_file[330] <= 8'h81
            reg_file[331] <= 8'h00
            reg_file[332] <= 8'h93
            reg_file[333] <= 8'h07
            reg_file[334] <= 8'hF0
            reg_file[335] <= 8'hFF
            reg_file[336] <= 8'h6B
            reg_file[337] <= 8'h80
            reg_file[338] <= 8'h07
            reg_file[339] <= 8'h00
            reg_file[340] <= 8'h13
            reg_file[341] <= 8'h06
            reg_file[342] <= 8'h00
            reg_file[343] <= 8'h00
            reg_file[344] <= 8'h13
            reg_file[345] <= 8'h05
            reg_file[346] <= 8'h02
            reg_file[347] <= 8'h00
            reg_file[348] <= 8'h97
            reg_file[349] <= 8'h15
            reg_file[350] <= 8'h00
            reg_file[351] <= 8'h00
            reg_file[352] <= 8'h93
            reg_file[353] <= 8'h85
            reg_file[354] <= 8'h45
            reg_file[355] <= 8'hEA
            reg_file[356] <= 8'h13
            reg_file[357] <= 8'h04
            reg_file[358] <= 8'h02
            reg_file[359] <= 8'h00
            reg_file[360] <= 8'hEF
            reg_file[361] <= 8'h00
            reg_file[362] <= 8'h90
            reg_file[363] <= 8'h06
            reg_file[364] <= 8'h13
            reg_file[365] <= 8'h05
            reg_file[366] <= 8'h00
            reg_file[367] <= 8'h00
            reg_file[368] <= 8'h13
            reg_file[369] <= 8'h06
            reg_file[370] <= 8'h00
            reg_file[371] <= 8'h00
            reg_file[372] <= 8'h93
            reg_file[373] <= 8'h05
            reg_file[374] <= 8'h00
            reg_file[375] <= 8'h00
            reg_file[376] <= 8'h33
            reg_file[377] <= 8'h05
            reg_file[378] <= 8'hA4
            reg_file[379] <= 8'h00
            reg_file[380] <= 8'hEF
            reg_file[381] <= 8'h00
            reg_file[382] <= 8'h10
            reg_file[383] <= 8'h17
            reg_file[384] <= 8'hF3
            reg_file[385] <= 8'h27
            reg_file[386] <= 8'h30
            reg_file[387] <= 8'hCC
            reg_file[388] <= 8'h93
            reg_file[389] <= 8'hB7
            reg_file[390] <= 8'h17
            reg_file[391] <= 8'h00
            reg_file[392] <= 8'h6B
            reg_file[393] <= 8'h80
            reg_file[394] <= 8'h07
            reg_file[395] <= 8'h00
            reg_file[396] <= 8'h83
            reg_file[397] <= 8'h20
            reg_file[398] <= 8'hC1
            reg_file[399] <= 8'h00
            reg_file[400] <= 8'h03
            reg_file[401] <= 8'h24
            reg_file[402] <= 8'h81
            reg_file[403] <= 8'h00
            reg_file[404] <= 8'h13
            reg_file[405] <= 8'h01
            reg_file[406] <= 8'h01
            reg_file[407] <= 8'h01
            reg_file[408] <= 8'h67
            reg_file[409] <= 8'h80
            reg_file[410] <= 8'h00
            reg_file[411] <= 8'h00
            reg_file[412] <= 8'h13
            reg_file[413] <= 8'h01
            reg_file[414] <= 8'h01
            reg_file[415] <= 8'hFF
            reg_file[416] <= 8'h23
            reg_file[417] <= 8'h24
            reg_file[418] <= 8'h81
            reg_file[419] <= 8'h00
            reg_file[420] <= 8'h23
            reg_file[421] <= 8'h20
            reg_file[422] <= 8'h21
            reg_file[423] <= 8'h01
            reg_file[424] <= 8'h17
            reg_file[425] <= 8'h14
            reg_file[426] <= 8'h00
            reg_file[427] <= 8'h00
            reg_file[428] <= 8'h13
            reg_file[429] <= 8'h04
            reg_file[430] <= 8'h84
            reg_file[431] <= 8'hE5
            reg_file[432] <= 8'h17
            reg_file[433] <= 8'h19
            reg_file[434] <= 8'h00
            reg_file[435] <= 8'h00
            reg_file[436] <= 8'h13
            reg_file[437] <= 8'h09
            reg_file[438] <= 8'h09
            reg_file[439] <= 8'hE5
            reg_file[440] <= 8'h33
            reg_file[441] <= 8'h09
            reg_file[442] <= 8'h89
            reg_file[443] <= 8'h40
            reg_file[444] <= 8'h23
            reg_file[445] <= 8'h26
            reg_file[446] <= 8'h11
            reg_file[447] <= 8'h00
            reg_file[448] <= 8'h23
            reg_file[449] <= 8'h22
            reg_file[450] <= 8'h91
            reg_file[451] <= 8'h00
            reg_file[452] <= 8'h13
            reg_file[453] <= 8'h59
            reg_file[454] <= 8'h29
            reg_file[455] <= 8'h40
            reg_file[456] <= 8'h63
            reg_file[457] <= 8'h0E
            reg_file[458] <= 8'h09
            reg_file[459] <= 8'h00
            reg_file[460] <= 8'h93
            reg_file[461] <= 8'h04
            reg_file[462] <= 8'h00
            reg_file[463] <= 8'h00
            reg_file[464] <= 8'h83
            reg_file[465] <= 8'h27
            reg_file[466] <= 8'h04
            reg_file[467] <= 8'h00
            reg_file[468] <= 8'h93
            reg_file[469] <= 8'h84
            reg_file[470] <= 8'h14
            reg_file[471] <= 8'h00
            reg_file[472] <= 8'h13
            reg_file[473] <= 8'h04
            reg_file[474] <= 8'h44
            reg_file[475] <= 8'h00
            reg_file[476] <= 8'hE7
            reg_file[477] <= 8'h80
            reg_file[478] <= 8'h07
            reg_file[479] <= 8'h00
            reg_file[480] <= 8'hE3
            reg_file[481] <= 8'h18
            reg_file[482] <= 8'h99
            reg_file[483] <= 8'hFE
            reg_file[484] <= 8'h17
            reg_file[485] <= 8'h14
            reg_file[486] <= 8'h00
            reg_file[487] <= 8'h00
            reg_file[488] <= 8'h13
            reg_file[489] <= 8'h04
            reg_file[490] <= 8'hC4
            reg_file[491] <= 8'hE1
            reg_file[492] <= 8'h17
            reg_file[493] <= 8'h19
            reg_file[494] <= 8'h00
            reg_file[495] <= 8'h00
            reg_file[496] <= 8'h13
            reg_file[497] <= 8'h09
            reg_file[498] <= 8'h89
            reg_file[499] <= 8'hE1
            reg_file[500] <= 8'h33
            reg_file[501] <= 8'h09
            reg_file[502] <= 8'h89
            reg_file[503] <= 8'h40
            reg_file[504] <= 8'h13
            reg_file[505] <= 8'h59
            reg_file[506] <= 8'h29
            reg_file[507] <= 8'h40
            reg_file[508] <= 8'h63
            reg_file[509] <= 8'h0E
            reg_file[510] <= 8'h09
            reg_file[511] <= 8'h00
            reg_file[512] <= 8'h93
            reg_file[513] <= 8'h04
            reg_file[514] <= 8'h00
            reg_file[515] <= 8'h00
            reg_file[516] <= 8'h83
            reg_file[517] <= 8'h27
            reg_file[518] <= 8'h04
            reg_file[519] <= 8'h00
            reg_file[520] <= 8'h93
            reg_file[521] <= 8'h84
            reg_file[522] <= 8'h14
            reg_file[523] <= 8'h00
            reg_file[524] <= 8'h13
            reg_file[525] <= 8'h04
            reg_file[526] <= 8'h44
            reg_file[527] <= 8'h00
            reg_file[528] <= 8'hE7
            reg_file[529] <= 8'h80
            reg_file[530] <= 8'h07
            reg_file[531] <= 8'h00
            reg_file[532] <= 8'hE3
            reg_file[533] <= 8'h18
            reg_file[534] <= 8'h99
            reg_file[535] <= 8'hFE
            reg_file[536] <= 8'h83
            reg_file[537] <= 8'h20
            reg_file[538] <= 8'hC1
            reg_file[539] <= 8'h00
            reg_file[540] <= 8'h03
            reg_file[541] <= 8'h24
            reg_file[542] <= 8'h81
            reg_file[543] <= 8'h00
            reg_file[544] <= 8'h83
            reg_file[545] <= 8'h24
            reg_file[546] <= 8'h41
            reg_file[547] <= 8'h00
            reg_file[548] <= 8'h03
            reg_file[549] <= 8'h29
            reg_file[550] <= 8'h01
            reg_file[551] <= 8'h00
            reg_file[552] <= 8'h13
            reg_file[553] <= 8'h01
            reg_file[554] <= 8'h01
            reg_file[555] <= 8'h01
            reg_file[556] <= 8'h67
            reg_file[557] <= 8'h80
            reg_file[558] <= 8'h00
            reg_file[559] <= 8'h00
            reg_file[560] <= 8'h13
            reg_file[561] <= 8'h01
            reg_file[562] <= 8'h01
            reg_file[563] <= 8'hFF
            reg_file[564] <= 8'h23
            reg_file[565] <= 8'h24
            reg_file[566] <= 8'h81
            reg_file[567] <= 8'h00
            reg_file[568] <= 8'h97
            reg_file[569] <= 8'h17
            reg_file[570] <= 8'h00
            reg_file[571] <= 8'h00
            reg_file[572] <= 8'h93
            reg_file[573] <= 8'h87
            reg_file[574] <= 8'hC7
            reg_file[575] <= 8'hDC
            reg_file[576] <= 8'h17
            reg_file[577] <= 8'h14
            reg_file[578] <= 8'h00
            reg_file[579] <= 8'h00
            reg_file[580] <= 8'h13
            reg_file[581] <= 8'h04
            reg_file[582] <= 8'h44
            reg_file[583] <= 8'hDC
            reg_file[584] <= 8'hB3
            reg_file[585] <= 8'h87
            reg_file[586] <= 8'h87
            reg_file[587] <= 8'h40
            reg_file[588] <= 8'h23
            reg_file[589] <= 8'h22
            reg_file[590] <= 8'h91
            reg_file[591] <= 8'h00
            reg_file[592] <= 8'h23
            reg_file[593] <= 8'h26
            reg_file[594] <= 8'h11
            reg_file[595] <= 8'h00
            reg_file[596] <= 8'h93
            reg_file[597] <= 8'hD4
            reg_file[598] <= 8'h27
            reg_file[599] <= 8'h40
            reg_file[600] <= 8'h63
            reg_file[601] <= 8'h80
            reg_file[602] <= 8'h04
            reg_file[603] <= 8'h02
            reg_file[604] <= 8'h93
            reg_file[605] <= 8'h87
            reg_file[606] <= 8'hC7
            reg_file[607] <= 8'hFF
            reg_file[608] <= 8'h33
            reg_file[609] <= 8'h84
            reg_file[610] <= 8'h87
            reg_file[611] <= 8'h00
            reg_file[612] <= 8'h83
            reg_file[613] <= 8'h27
            reg_file[614] <= 8'h04
            reg_file[615] <= 8'h00
            reg_file[616] <= 8'h93
            reg_file[617] <= 8'h84
            reg_file[618] <= 8'hF4
            reg_file[619] <= 8'hFF
            reg_file[620] <= 8'h13
            reg_file[621] <= 8'h04
            reg_file[622] <= 8'hC4
            reg_file[623] <= 8'hFF
            reg_file[624] <= 8'hE7
            reg_file[625] <= 8'h80
            reg_file[626] <= 8'h07
            reg_file[627] <= 8'h00
            reg_file[628] <= 8'hE3
            reg_file[629] <= 8'h98
            reg_file[630] <= 8'h04
            reg_file[631] <= 8'hFE
            reg_file[632] <= 8'h83
            reg_file[633] <= 8'h20
            reg_file[634] <= 8'hC1
            reg_file[635] <= 8'h00
            reg_file[636] <= 8'h03
            reg_file[637] <= 8'h24
            reg_file[638] <= 8'h81
            reg_file[639] <= 8'h00
            reg_file[640] <= 8'h83
            reg_file[641] <= 8'h24
            reg_file[642] <= 8'h41
            reg_file[643] <= 8'h00
            reg_file[644] <= 8'h13
            reg_file[645] <= 8'h01
            reg_file[646] <= 8'h01
            reg_file[647] <= 8'h01
            reg_file[648] <= 8'h67
            reg_file[649] <= 8'h80
            reg_file[650] <= 8'h00
            reg_file[651] <= 8'h00
            reg_file[652] <= 8'h13
            reg_file[653] <= 8'h01
            reg_file[654] <= 8'h01
            reg_file[655] <= 8'hFF
            reg_file[656] <= 8'h23
            reg_file[657] <= 8'h26
            reg_file[658] <= 8'h11
            reg_file[659] <= 8'h00
            reg_file[660] <= 8'h23
            reg_file[661] <= 8'h24
            reg_file[662] <= 8'h81
            reg_file[663] <= 8'h00
            reg_file[664] <= 8'h23
            reg_file[665] <= 8'h22
            reg_file[666] <= 8'h91
            reg_file[667] <= 8'h00
            reg_file[668] <= 8'h23
            reg_file[669] <= 8'h20
            reg_file[670] <= 8'h21
            reg_file[671] <= 8'h01
            reg_file[672] <= 8'hF3
            reg_file[673] <= 8'h27
            reg_file[674] <= 8'h50
            reg_file[675] <= 8'hCC
            reg_file[676] <= 8'h73
            reg_file[677] <= 8'h27
            reg_file[678] <= 8'h30
            reg_file[679] <= 8'hCC
            reg_file[680] <= 8'hF3
            reg_file[681] <= 8'h26
            reg_file[682] <= 8'h00
            reg_file[683] <= 8'hCC
            reg_file[684] <= 8'hF3
            reg_file[685] <= 8'h25
            reg_file[686] <= 8'h00
            reg_file[687] <= 8'hFC
            reg_file[688] <= 8'h13
            reg_file[689] <= 8'h96
            reg_file[690] <= 8'h27
            reg_file[691] <= 8'h00
            reg_file[692] <= 8'h97
            reg_file[693] <= 8'h17
            reg_file[694] <= 8'h00
            reg_file[695] <= 8'h00
            reg_file[696] <= 8'h93
            reg_file[697] <= 8'h87
            reg_file[698] <= 8'hC7
            reg_file[699] <= 8'h18
            reg_file[700] <= 8'hB3
            reg_file[701] <= 8'h87
            reg_file[702] <= 8'hC7
            reg_file[703] <= 8'h00
            reg_file[704] <= 8'h83
            reg_file[705] <= 8'hA4
            reg_file[706] <= 8'h07
            reg_file[707] <= 8'h00
            reg_file[708] <= 8'h03
            reg_file[709] <= 8'hA4
            reg_file[710] <= 8'h04
            reg_file[711] <= 8'h01
            reg_file[712] <= 8'h03
            reg_file[713] <= 8'hA6
            reg_file[714] <= 8'hC4
            reg_file[715] <= 8'h00
            reg_file[716] <= 8'h33
            reg_file[717] <= 8'h29
            reg_file[718] <= 8'h87
            reg_file[719] <= 8'h00
            reg_file[720] <= 8'h93
            reg_file[721] <= 8'h07
            reg_file[722] <= 8'h04
            reg_file[723] <= 8'h00
            reg_file[724] <= 8'h33
            reg_file[725] <= 8'h09
            reg_file[726] <= 8'hC9
            reg_file[727] <= 8'h00
            reg_file[728] <= 8'h33
            reg_file[729] <= 8'h04
            reg_file[730] <= 8'hE6
            reg_file[731] <= 8'h02
            reg_file[732] <= 8'h63
            reg_file[733] <= 8'h54
            reg_file[734] <= 8'hF7
            reg_file[735] <= 8'h00
            reg_file[736] <= 8'h93
            reg_file[737] <= 8'h07
            reg_file[738] <= 8'h07
            reg_file[739] <= 8'h00
            reg_file[740] <= 8'h33
            reg_file[741] <= 8'h04
            reg_file[742] <= 8'hF4
            reg_file[743] <= 8'h00
            reg_file[744] <= 8'h03
            reg_file[745] <= 8'hA7
            reg_file[746] <= 8'h84
            reg_file[747] <= 8'h00
            reg_file[748] <= 8'h33
            reg_file[749] <= 8'h04
            reg_file[750] <= 8'hB4
            reg_file[751] <= 8'h02
            reg_file[752] <= 8'hB3
            reg_file[753] <= 8'h07
            reg_file[754] <= 8'hD9
            reg_file[755] <= 8'h02
            reg_file[756] <= 8'h33
            reg_file[757] <= 8'h04
            reg_file[758] <= 8'hE4
            reg_file[759] <= 8'h00
            reg_file[760] <= 8'h33
            reg_file[761] <= 8'h04
            reg_file[762] <= 8'hF4
            reg_file[763] <= 8'h00
            reg_file[764] <= 8'h33
            reg_file[765] <= 8'h09
            reg_file[766] <= 8'h89
            reg_file[767] <= 8'h00
            reg_file[768] <= 8'h63
            reg_file[769] <= 8'h5E
            reg_file[770] <= 8'h24
            reg_file[771] <= 8'h01
            reg_file[772] <= 8'h83
            reg_file[773] <= 8'hA7
            reg_file[774] <= 8'h04
            reg_file[775] <= 8'h00
            reg_file[776] <= 8'h83
            reg_file[777] <= 8'hA5
            reg_file[778] <= 8'h44
            reg_file[779] <= 8'h00
            reg_file[780] <= 8'h13
            reg_file[781] <= 8'h05
            reg_file[782] <= 8'h04
            reg_file[783] <= 8'h00
            reg_file[784] <= 8'h13
            reg_file[785] <= 8'h04
            reg_file[786] <= 8'h14
            reg_file[787] <= 8'h00
            reg_file[788] <= 8'hE7
            reg_file[789] <= 8'h80
            reg_file[790] <= 8'h07
            reg_file[791] <= 8'h00
            reg_file[792] <= 8'hE3
            reg_file[793] <= 8'h16
            reg_file[794] <= 8'h89
            reg_file[795] <= 8'hFE
            reg_file[796] <= 8'h03
            reg_file[797] <= 8'hA7
            reg_file[798] <= 8'h44
            reg_file[799] <= 8'h01
            reg_file[800] <= 8'h93
            reg_file[801] <= 8'h07
            reg_file[802] <= 8'h00
            reg_file[803] <= 8'h00
            reg_file[804] <= 8'h6B
            reg_file[805] <= 8'hC0
            reg_file[806] <= 8'hE7
            reg_file[807] <= 8'h00
            reg_file[808] <= 8'h83
            reg_file[809] <= 8'h20
            reg_file[810] <= 8'hC1
            reg_file[811] <= 8'h00
            reg_file[812] <= 8'h03
            reg_file[813] <= 8'h24
            reg_file[814] <= 8'h81
            reg_file[815] <= 8'h00
            reg_file[816] <= 8'h83
            reg_file[817] <= 8'h24
            reg_file[818] <= 8'h41
            reg_file[819] <= 8'h00
            reg_file[820] <= 8'h03
            reg_file[821] <= 8'h29
            reg_file[822] <= 8'h01
            reg_file[823] <= 8'h00
            reg_file[824] <= 8'h13
            reg_file[825] <= 8'h01
            reg_file[826] <= 8'h01
            reg_file[827] <= 8'h01
            reg_file[828] <= 8'h67
            reg_file[829] <= 8'h80
            reg_file[830] <= 8'h00
            reg_file[831] <= 8'h00
            reg_file[832] <= 8'hF3
            reg_file[833] <= 8'h27
            reg_file[834] <= 8'h50
            reg_file[835] <= 8'hCC
            reg_file[836] <= 8'h73
            reg_file[837] <= 8'h25
            reg_file[838] <= 8'h20
            reg_file[839] <= 8'hCC
            reg_file[840] <= 8'h13
            reg_file[841] <= 8'h97
            reg_file[842] <= 8'h27
            reg_file[843] <= 8'h00
            reg_file[844] <= 8'h97
            reg_file[845] <= 8'h17
            reg_file[846] <= 8'h00
            reg_file[847] <= 8'h00
            reg_file[848] <= 8'h93
            reg_file[849] <= 8'h87
            reg_file[850] <= 8'h47
            reg_file[851] <= 8'h0F
            reg_file[852] <= 8'hB3
            reg_file[853] <= 8'h87
            reg_file[854] <= 8'hE7
            reg_file[855] <= 8'h00
            reg_file[856] <= 8'h83
            reg_file[857] <= 8'hA7
            reg_file[858] <= 8'h07
            reg_file[859] <= 8'h00
            reg_file[860] <= 8'h03
            reg_file[861] <= 8'hA7
            reg_file[862] <= 8'h87
            reg_file[863] <= 8'h00
            reg_file[864] <= 8'h03
            reg_file[865] <= 8'hA3
            reg_file[866] <= 8'h07
            reg_file[867] <= 8'h00
            reg_file[868] <= 8'h83
            reg_file[869] <= 8'hA5
            reg_file[870] <= 8'h47
            reg_file[871] <= 8'h00
            reg_file[872] <= 8'h33
            reg_file[873] <= 8'h05
            reg_file[874] <= 8'hE5
            reg_file[875] <= 8'h00
            reg_file[876] <= 8'h67
            reg_file[877] <= 8'h00
            reg_file[878] <= 8'h03
            reg_file[879] <= 8'h00
            reg_file[880] <= 8'h13
            reg_file[881] <= 8'h01
            reg_file[882] <= 8'h01
            reg_file[883] <= 8'hFF
            reg_file[884] <= 8'h23
            reg_file[885] <= 8'h26
            reg_file[886] <= 8'h11
            reg_file[887] <= 8'h00
            reg_file[888] <= 8'h93
            reg_file[889] <= 8'h07
            reg_file[890] <= 8'hF0
            reg_file[891] <= 8'hFF
            reg_file[892] <= 8'h6B
            reg_file[893] <= 8'h80
            reg_file[894] <= 8'h07
            reg_file[895] <= 8'h00
            reg_file[896] <= 8'hEF
            reg_file[897] <= 8'hF0
            reg_file[898] <= 8'hDF
            reg_file[899] <= 8'hF0
            reg_file[900] <= 8'hF3
            reg_file[901] <= 8'h27
            reg_file[902] <= 8'h30
            reg_file[903] <= 8'hCC
            reg_file[904] <= 8'h93
            reg_file[905] <= 8'hB7
            reg_file[906] <= 8'h17
            reg_file[907] <= 8'h00
            reg_file[908] <= 8'h6B
            reg_file[909] <= 8'h80
            reg_file[910] <= 8'h07
            reg_file[911] <= 8'h00
            reg_file[912] <= 8'h83
            reg_file[913] <= 8'h20
            reg_file[914] <= 8'hC1
            reg_file[915] <= 8'h00
            reg_file[916] <= 8'h13
            reg_file[917] <= 8'h01
            reg_file[918] <= 8'h01
            reg_file[919] <= 8'h01
            reg_file[920] <= 8'h67
            reg_file[921] <= 8'h80
            reg_file[922] <= 8'h00
            reg_file[923] <= 8'h00
            reg_file[924] <= 8'h13
            reg_file[925] <= 8'h01
            reg_file[926] <= 8'h01
            reg_file[927] <= 8'hFE
            reg_file[928] <= 8'h23
            reg_file[929] <= 8'h2E
            reg_file[930] <= 8'h11
            reg_file[931] <= 8'h00
            reg_file[932] <= 8'h23
            reg_file[933] <= 8'h2C
            reg_file[934] <= 8'h81
            reg_file[935] <= 8'h00
            reg_file[936] <= 8'h23
            reg_file[937] <= 8'h2A
            reg_file[938] <= 8'h91
            reg_file[939] <= 8'h00
            reg_file[940] <= 8'h23
            reg_file[941] <= 8'h28
            reg_file[942] <= 8'h21
            reg_file[943] <= 8'h01
            reg_file[944] <= 8'h23
            reg_file[945] <= 8'h26
            reg_file[946] <= 8'h31
            reg_file[947] <= 8'h01
            reg_file[948] <= 8'h23
            reg_file[949] <= 8'h24
            reg_file[950] <= 8'h41
            reg_file[951] <= 8'h01
            reg_file[952] <= 8'hF3
            reg_file[953] <= 8'h27
            reg_file[954] <= 8'h50
            reg_file[955] <= 8'hCC
            reg_file[956] <= 8'h73
            reg_file[957] <= 8'h27
            reg_file[958] <= 8'h30
            reg_file[959] <= 8'hCC
            reg_file[960] <= 8'hF3
            reg_file[961] <= 8'h26
            reg_file[962] <= 8'h00
            reg_file[963] <= 8'hCC
            reg_file[964] <= 8'h73
            reg_file[965] <= 8'h25
            reg_file[966] <= 8'h00
            reg_file[967] <= 8'hFC
            reg_file[968] <= 8'h13
            reg_file[969] <= 8'h96
            reg_file[970] <= 8'h27
            reg_file[971] <= 8'h00
            reg_file[972] <= 8'h97
            reg_file[973] <= 8'h17
            reg_file[974] <= 8'h00
            reg_file[975] <= 8'h00
            reg_file[976] <= 8'h93
            reg_file[977] <= 8'h87
            reg_file[978] <= 8'h47
            reg_file[979] <= 8'h07
            reg_file[980] <= 8'hB3
            reg_file[981] <= 8'h87
            reg_file[982] <= 8'hC7
            reg_file[983] <= 8'h00
            reg_file[984] <= 8'h03
            reg_file[985] <= 8'hA4
            reg_file[986] <= 8'h07
            reg_file[987] <= 8'h00
            reg_file[988] <= 8'h83
            reg_file[989] <= 8'h24
            reg_file[990] <= 8'h44
            reg_file[991] <= 8'h01
            reg_file[992] <= 8'h03
            reg_file[993] <= 8'h26
            reg_file[994] <= 8'h04
            reg_file[995] <= 8'h01
            reg_file[996] <= 8'h33
            reg_file[997] <= 8'h2A
            reg_file[998] <= 8'h97
            reg_file[999] <= 8'h00
            reg_file[1000] <= 8'h93
            reg_file[1001] <= 8'h87
            reg_file[1002] <= 8'h04
            reg_file[1003] <= 8'h00
            reg_file[1004] <= 8'h33
            reg_file[1005] <= 8'h0A
            reg_file[1006] <= 8'hCA
            reg_file[1007] <= 8'h00
            reg_file[1008] <= 8'hB3
            reg_file[1009] <= 8'h04
            reg_file[1010] <= 8'hE6
            reg_file[1011] <= 8'h02
            reg_file[1012] <= 8'h63
            reg_file[1013] <= 8'h54
            reg_file[1014] <= 8'hF7
            reg_file[1015] <= 8'h00
            reg_file[1016] <= 8'h93
            reg_file[1017] <= 8'h07
            reg_file[1018] <= 8'h07
            reg_file[1019] <= 8'h00
            reg_file[1020] <= 8'hB3
            reg_file[1021] <= 8'h84
            reg_file[1022] <= 8'hF4
            reg_file[1023] <= 8'h00
            reg_file[1024] <= 8'h83
            reg_file[1025] <= 8'h25
            reg_file[1026] <= 8'h04
            reg_file[1027] <= 8'h00
            reg_file[1028] <= 8'h03
            reg_file[1029] <= 8'h27
            reg_file[1030] <= 8'hC4
            reg_file[1031] <= 8'h00
            reg_file[1032] <= 8'h03
            reg_file[1033] <= 8'hA9
            reg_file[1034] <= 8'h05
            reg_file[1035] <= 8'h00
            reg_file[1036] <= 8'h83
            reg_file[1037] <= 8'hA9
            reg_file[1038] <= 8'h45
            reg_file[1039] <= 8'h00
            reg_file[1040] <= 8'hB3
            reg_file[1041] <= 8'h84
            reg_file[1042] <= 8'hA4
            reg_file[1043] <= 8'h02
            reg_file[1044] <= 8'hB3
            reg_file[1045] <= 8'h07
            reg_file[1046] <= 8'hDA
            reg_file[1047] <= 8'h02
            reg_file[1048] <= 8'hB3
            reg_file[1049] <= 8'h84
            reg_file[1050] <= 8'hE4
            reg_file[1051] <= 8'h00
            reg_file[1052] <= 8'hB3
            reg_file[1053] <= 8'h84
            reg_file[1054] <= 8'hF4
            reg_file[1055] <= 8'h00
            reg_file[1056] <= 8'h33
            reg_file[1057] <= 8'h0A
            reg_file[1058] <= 8'h9A
            reg_file[1059] <= 8'h00
            reg_file[1060] <= 8'hB3
            reg_file[1061] <= 8'h09
            reg_file[1062] <= 8'h39
            reg_file[1063] <= 8'h03
            reg_file[1064] <= 8'h63
            reg_file[1065] <= 8'hC0
            reg_file[1066] <= 8'h44
            reg_file[1067] <= 8'h07
            reg_file[1068] <= 8'h6F
            reg_file[1069] <= 8'h00
            reg_file[1070] <= 8'h00
            reg_file[1071] <= 8'h08
            reg_file[1072] <= 8'h03
            reg_file[1073] <= 8'h47
            reg_file[1074] <= 8'hE4
            reg_file[1075] <= 8'h01
            reg_file[1076] <= 8'h83
            reg_file[1077] <= 8'h46
            reg_file[1078] <= 8'hD4
            reg_file[1079] <= 8'h01
            reg_file[1080] <= 8'h33
            reg_file[1081] <= 8'hD7
            reg_file[1082] <= 8'hE4
            reg_file[1083] <= 8'h40
            reg_file[1084] <= 8'hB3
            reg_file[1085] <= 8'h07
            reg_file[1086] <= 8'h37
            reg_file[1087] <= 8'h03
            reg_file[1088] <= 8'hB3
            reg_file[1089] <= 8'h87
            reg_file[1090] <= 8'hF4
            reg_file[1091] <= 8'h40
            reg_file[1092] <= 8'h63
            reg_file[1093] <= 8'h80
            reg_file[1094] <= 8'h06
            reg_file[1095] <= 8'h06
            reg_file[1096] <= 8'h83
            reg_file[1097] <= 8'h46
            reg_file[1098] <= 8'hF4
            reg_file[1099] <= 8'h01
            reg_file[1100] <= 8'hB3
            reg_file[1101] <= 8'hD6
            reg_file[1102] <= 8'hD7
            reg_file[1103] <= 8'h40
            reg_file[1104] <= 8'hB3
            reg_file[1105] <= 8'h88
            reg_file[1106] <= 8'h26
            reg_file[1107] <= 8'h03
            reg_file[1108] <= 8'h03
            reg_file[1109] <= 8'hAE
            reg_file[1110] <= 8'h45
            reg_file[1111] <= 8'h01
            reg_file[1112] <= 8'h03
            reg_file[1113] <= 8'hA3
            reg_file[1114] <= 8'h05
            reg_file[1115] <= 8'h01
            reg_file[1116] <= 8'h03
            reg_file[1117] <= 8'hA6
            reg_file[1118] <= 8'hC5
            reg_file[1119] <= 8'h00
            reg_file[1120] <= 8'h03
            reg_file[1121] <= 8'h28
            reg_file[1122] <= 8'h44
            reg_file[1123] <= 8'h00
            reg_file[1124] <= 8'h03
            reg_file[1125] <= 8'h25
            reg_file[1126] <= 8'h84
            reg_file[1127] <= 8'h00
            reg_file[1128] <= 8'h93
            reg_file[1129] <= 8'h84
            reg_file[1130] <= 8'h14
            reg_file[1131] <= 8'h00
            reg_file[1132] <= 8'h33
            reg_file[1133] <= 8'h07
            reg_file[1134] <= 8'hC7
            reg_file[1135] <= 8'h01
            reg_file[1136] <= 8'hB3
            reg_file[1137] <= 8'h86
            reg_file[1138] <= 8'h66
            reg_file[1139] <= 8'h00
            reg_file[1140] <= 8'hB3
            reg_file[1141] <= 8'h87
            reg_file[1142] <= 8'h17
            reg_file[1143] <= 8'h41
            reg_file[1144] <= 8'h33
            reg_file[1145] <= 8'h86
            reg_file[1146] <= 8'hC7
            reg_file[1147] <= 8'h00
            reg_file[1148] <= 8'hE7
            reg_file[1149] <= 8'h00
            reg_file[1150] <= 8'h08
            reg_file[1151] <= 8'h00
            reg_file[1152] <= 8'h63
            reg_file[1153] <= 8'h06
            reg_file[1154] <= 8'h9A
            reg_file[1155] <= 8'h02
            reg_file[1156] <= 8'h83
            reg_file[1157] <= 8'h25
            reg_file[1158] <= 8'h04
            reg_file[1159] <= 8'h00
            reg_file[1160] <= 8'h83
            reg_file[1161] <= 8'h47
            reg_file[1162] <= 8'hC4
            reg_file[1163] <= 8'h01
            reg_file[1164] <= 8'hE3
            reg_file[1165] <= 8'h92
            reg_file[1166] <= 8'h07
            reg_file[1167] <= 8'hFA
            reg_file[1168] <= 8'h33
            reg_file[1169] <= 8'hC7
            reg_file[1170] <= 8'h34
            reg_file[1171] <= 8'h03
            reg_file[1172] <= 8'h83
            reg_file[1173] <= 8'h46
            reg_file[1174] <= 8'hD4
            reg_file[1175] <= 8'h01
            reg_file[1176] <= 8'hB3
            reg_file[1177] <= 8'h07
            reg_file[1178] <= 8'h37
            reg_file[1179] <= 8'h03
            reg_file[1180] <= 8'hB3
            reg_file[1181] <= 8'h87
            reg_file[1182] <= 8'hF4
            reg_file[1183] <= 8'h40
            reg_file[1184] <= 8'hE3
            reg_file[1185] <= 8'h94
            reg_file[1186] <= 8'h06
            reg_file[1187] <= 8'hFA
            reg_file[1188] <= 8'hB3
            reg_file[1189] <= 8'hC6
            reg_file[1190] <= 8'h27
            reg_file[1191] <= 8'h03
            reg_file[1192] <= 8'h6F
            reg_file[1193] <= 8'hF0
            reg_file[1194] <= 8'h9F
            reg_file[1195] <= 8'hFA
            reg_file[1196] <= 8'h03
            reg_file[1197] <= 8'h27
            reg_file[1198] <= 8'h84
            reg_file[1199] <= 8'h01
            reg_file[1200] <= 8'h93
            reg_file[1201] <= 8'h07
            reg_file[1202] <= 8'h00
            reg_file[1203] <= 8'h00
            reg_file[1204] <= 8'h6B
            reg_file[1205] <= 8'hC0
            reg_file[1206] <= 8'hE7
            reg_file[1207] <= 8'h00
            reg_file[1208] <= 8'h83
            reg_file[1209] <= 8'h20
            reg_file[1210] <= 8'hC1
            reg_file[1211] <= 8'h01
            reg_file[1212] <= 8'h03
            reg_file[1213] <= 8'h24
            reg_file[1214] <= 8'h81
            reg_file[1215] <= 8'h01
            reg_file[1216] <= 8'h83
            reg_file[1217] <= 8'h24
            reg_file[1218] <= 8'h41
            reg_file[1219] <= 8'h01
            reg_file[1220] <= 8'h03
            reg_file[1221] <= 8'h29
            reg_file[1222] <= 8'h01
            reg_file[1223] <= 8'h01
            reg_file[1224] <= 8'h83
            reg_file[1225] <= 8'h29
            reg_file[1226] <= 8'hC1
            reg_file[1227] <= 8'h00
            reg_file[1228] <= 8'h03
            reg_file[1229] <= 8'h2A
            reg_file[1230] <= 8'h81
            reg_file[1231] <= 8'h00
            reg_file[1232] <= 8'h13
            reg_file[1233] <= 8'h01
            reg_file[1234] <= 8'h01
            reg_file[1235] <= 8'h02
            reg_file[1236] <= 8'h67
            reg_file[1237] <= 8'h80
            reg_file[1238] <= 8'h00
            reg_file[1239] <= 8'h00
            reg_file[1240] <= 8'h73
            reg_file[1241] <= 8'h27
            reg_file[1242] <= 8'h50
            reg_file[1243] <= 8'hCC
            reg_file[1244] <= 8'hF3
            reg_file[1245] <= 8'h27
            reg_file[1246] <= 8'h20
            reg_file[1247] <= 8'hCC
            reg_file[1248] <= 8'h93
            reg_file[1249] <= 8'h16
            reg_file[1250] <= 8'h27
            reg_file[1251] <= 8'h00
            reg_file[1252] <= 8'h17
            reg_file[1253] <= 8'h17
            reg_file[1254] <= 8'h00
            reg_file[1255] <= 8'h00
            reg_file[1256] <= 8'h13
            reg_file[1257] <= 8'h07
            reg_file[1258] <= 8'hC7
            reg_file[1259] <= 8'hF5
            reg_file[1260] <= 8'h33
            reg_file[1261] <= 8'h07
            reg_file[1262] <= 8'hD7
            reg_file[1263] <= 8'h00
            reg_file[1264] <= 8'h03
            reg_file[1265] <= 8'h25
            reg_file[1266] <= 8'h07
            reg_file[1267] <= 8'h00
            reg_file[1268] <= 8'h83
            reg_file[1269] <= 8'h25
            reg_file[1270] <= 8'h05
            reg_file[1271] <= 8'h00
            reg_file[1272] <= 8'h83
            reg_file[1273] <= 8'h26
            reg_file[1274] <= 8'hC5
            reg_file[1275] <= 8'h00
            reg_file[1276] <= 8'h03
            reg_file[1277] <= 8'h47
            reg_file[1278] <= 8'hC5
            reg_file[1279] <= 8'h01
            reg_file[1280] <= 8'h83
            reg_file[1281] <= 8'hA8
            reg_file[1282] <= 8'h05
            reg_file[1283] <= 8'h00
            reg_file[1284] <= 8'h03
            reg_file[1285] <= 8'hA6
            reg_file[1286] <= 8'h45
            reg_file[1287] <= 8'h00
            reg_file[1288] <= 8'hB3
            reg_file[1289] <= 8'h87
            reg_file[1290] <= 8'hD7
            reg_file[1291] <= 8'h00
            reg_file[1292] <= 8'h33
            reg_file[1293] <= 8'h86
            reg_file[1294] <= 8'hC8
            reg_file[1295] <= 8'h02
            reg_file[1296] <= 8'h63
            reg_file[1297] <= 8'h08
            reg_file[1298] <= 8'h07
            reg_file[1299] <= 8'h04
            reg_file[1300] <= 8'h03
            reg_file[1301] <= 8'h47
            reg_file[1302] <= 8'hE5
            reg_file[1303] <= 8'h01
            reg_file[1304] <= 8'h83
            reg_file[1305] <= 8'h46
            reg_file[1306] <= 8'hD5
            reg_file[1307] <= 8'h01
            reg_file[1308] <= 8'h33
            reg_file[1309] <= 8'hD7
            reg_file[1310] <= 8'hE7
            reg_file[1311] <= 8'h40
            reg_file[1312] <= 8'h33
            reg_file[1313] <= 8'h06
            reg_file[1314] <= 8'hC7
            reg_file[1315] <= 8'h02
            reg_file[1316] <= 8'hB3
            reg_file[1317] <= 8'h87
            reg_file[1318] <= 8'hC7
            reg_file[1319] <= 8'h40
            reg_file[1320] <= 8'h63
            reg_file[1321] <= 8'h86
            reg_file[1322] <= 8'h06
            reg_file[1323] <= 8'h04
            reg_file[1324] <= 8'h83
            reg_file[1325] <= 8'h46
            reg_file[1326] <= 8'hF5
            reg_file[1327] <= 8'h01
            reg_file[1328] <= 8'h33
            reg_file[1329] <= 8'hD8
            reg_file[1330] <= 8'hD7
            reg_file[1331] <= 8'h40
            reg_file[1332] <= 8'h83
            reg_file[1333] <= 8'hA6
            reg_file[1334] <= 8'h05
            reg_file[1335] <= 8'h01
            reg_file[1336] <= 8'h03
            reg_file[1337] <= 8'hAE
            reg_file[1338] <= 8'h45
            reg_file[1339] <= 8'h01
            reg_file[1340] <= 8'h03
            reg_file[1341] <= 8'hA6
            reg_file[1342] <= 8'hC5
            reg_file[1343] <= 8'h00
            reg_file[1344] <= 8'hB3
            reg_file[1345] <= 8'h06
            reg_file[1346] <= 8'hD8
            reg_file[1347] <= 8'h00
            reg_file[1348] <= 8'h33
            reg_file[1349] <= 8'h08
            reg_file[1350] <= 8'h18
            reg_file[1351] <= 8'h03
            reg_file[1352] <= 8'h03
            reg_file[1353] <= 8'h23
            reg_file[1354] <= 8'h45
            reg_file[1355] <= 8'h00
            reg_file[1356] <= 8'h03
            reg_file[1357] <= 8'h25
            reg_file[1358] <= 8'h85
            reg_file[1359] <= 8'h00
            reg_file[1360] <= 8'h33
            reg_file[1361] <= 8'h07
            reg_file[1362] <= 8'hC7
            reg_file[1363] <= 8'h01
            reg_file[1364] <= 8'hB3
            reg_file[1365] <= 8'h87
            reg_file[1366] <= 8'h07
            reg_file[1367] <= 8'h41
            reg_file[1368] <= 8'h33
            reg_file[1369] <= 8'h86
            reg_file[1370] <= 8'hC7
            reg_file[1371] <= 8'h00
            reg_file[1372] <= 8'h67
            reg_file[1373] <= 8'h00
            reg_file[1374] <= 8'h03
            reg_file[1375] <= 8'h00
            reg_file[1376] <= 8'h33
            reg_file[1377] <= 8'hC7
            reg_file[1378] <= 8'hC7
            reg_file[1379] <= 8'h02
            reg_file[1380] <= 8'h83
            reg_file[1381] <= 8'h46
            reg_file[1382] <= 8'hD5
            reg_file[1383] <= 8'h01
            reg_file[1384] <= 8'h33
            reg_file[1385] <= 8'h06
            reg_file[1386] <= 8'hC7
            reg_file[1387] <= 8'h02
            reg_file[1388] <= 8'hB3
            reg_file[1389] <= 8'h87
            reg_file[1390] <= 8'hC7
            reg_file[1391] <= 8'h40
            reg_file[1392] <= 8'hE3
            reg_file[1393] <= 8'h9E
            reg_file[1394] <= 8'h06
            reg_file[1395] <= 8'hFA
            reg_file[1396] <= 8'h33
            reg_file[1397] <= 8'hC8
            reg_file[1398] <= 8'h17
            reg_file[1399] <= 8'h03
            reg_file[1400] <= 8'h6F
            reg_file[1401] <= 8'hF0
            reg_file[1402] <= 8'hDF
            reg_file[1403] <= 8'hFB
            reg_file[1404] <= 8'h13
            reg_file[1405] <= 8'h01
            reg_file[1406] <= 8'h01
            reg_file[1407] <= 8'hFF
            reg_file[1408] <= 8'h23
            reg_file[1409] <= 8'h26
            reg_file[1410] <= 8'h11
            reg_file[1411] <= 8'h00
            reg_file[1412] <= 8'h93
            reg_file[1413] <= 8'h07
            reg_file[1414] <= 8'hF0
            reg_file[1415] <= 8'hFF
            reg_file[1416] <= 8'h6B
            reg_file[1417] <= 8'h80
            reg_file[1418] <= 8'h07
            reg_file[1419] <= 8'h00
            reg_file[1420] <= 8'hEF
            reg_file[1421] <= 8'hF0
            reg_file[1422] <= 8'h1F
            reg_file[1423] <= 8'hE1
            reg_file[1424] <= 8'hF3
            reg_file[1425] <= 8'h27
            reg_file[1426] <= 8'h30
            reg_file[1427] <= 8'hCC
            reg_file[1428] <= 8'h93
            reg_file[1429] <= 8'hB7
            reg_file[1430] <= 8'h17
            reg_file[1431] <= 8'h00
            reg_file[1432] <= 8'h6B
            reg_file[1433] <= 8'h80
            reg_file[1434] <= 8'h07
            reg_file[1435] <= 8'h00
            reg_file[1436] <= 8'h83
            reg_file[1437] <= 8'h20
            reg_file[1438] <= 8'hC1
            reg_file[1439] <= 8'h00
            reg_file[1440] <= 8'h13
            reg_file[1441] <= 8'h01
            reg_file[1442] <= 8'h01
            reg_file[1443] <= 8'h01
            reg_file[1444] <= 8'h67
            reg_file[1445] <= 8'h80
            reg_file[1446] <= 8'h00
            reg_file[1447] <= 8'h00
            reg_file[1448] <= 8'h13
            reg_file[1449] <= 8'h01
            reg_file[1450] <= 8'h01
            reg_file[1451] <= 8'hFD
            reg_file[1452] <= 8'h23
            reg_file[1453] <= 8'h26
            reg_file[1454] <= 8'h11
            reg_file[1455] <= 8'h02
            reg_file[1456] <= 8'h23
            reg_file[1457] <= 8'h24
            reg_file[1458] <= 8'h81
            reg_file[1459] <= 8'h02
            reg_file[1460] <= 8'h23
            reg_file[1461] <= 8'h22
            reg_file[1462] <= 8'h91
            reg_file[1463] <= 8'h02
            reg_file[1464] <= 8'h23
            reg_file[1465] <= 8'h20
            reg_file[1466] <= 8'h21
            reg_file[1467] <= 8'h03
            reg_file[1468] <= 8'hF3
            reg_file[1469] <= 8'h26
            reg_file[1470] <= 8'h20
            reg_file[1471] <= 8'hFC
            reg_file[1472] <= 8'hF3
            reg_file[1473] <= 8'h28
            reg_file[1474] <= 8'h10
            reg_file[1475] <= 8'hFC
            reg_file[1476] <= 8'hF3
            reg_file[1477] <= 8'h24
            reg_file[1478] <= 8'h00
            reg_file[1479] <= 8'hFC
            reg_file[1480] <= 8'hF3
            reg_file[1481] <= 8'h27
            reg_file[1482] <= 8'h50
            reg_file[1483] <= 8'hCC
            reg_file[1484] <= 8'h13
            reg_file[1485] <= 8'h07
            reg_file[1486] <= 8'hF0
            reg_file[1487] <= 8'h01
            reg_file[1488] <= 8'h63
            reg_file[1489] <= 8'h48
            reg_file[1490] <= 8'hF7
            reg_file[1491] <= 8'h08
            reg_file[1492] <= 8'h33
            reg_file[1493] <= 8'h88
            reg_file[1494] <= 8'h14
            reg_file[1495] <= 8'h03
            reg_file[1496] <= 8'h13
            reg_file[1497] <= 8'h07
            reg_file[1498] <= 8'h10
            reg_file[1499] <= 8'h00
            reg_file[1500] <= 8'h63
            reg_file[1501] <= 8'h54
            reg_file[1502] <= 8'hA8
            reg_file[1503] <= 8'h00
            reg_file[1504] <= 8'h33
            reg_file[1505] <= 8'h47
            reg_file[1506] <= 8'h05
            reg_file[1507] <= 8'h03
            reg_file[1508] <= 8'h63
            reg_file[1509] <= 8'hCA
            reg_file[1510] <= 8'hE6
            reg_file[1511] <= 8'h08
            reg_file[1512] <= 8'h63
            reg_file[1513] <= 8'hDC
            reg_file[1514] <= 8'hE7
            reg_file[1515] <= 8'h06
            reg_file[1516] <= 8'h93
            reg_file[1517] <= 8'h86
            reg_file[1518] <= 8'hF6
            reg_file[1519] <= 8'hFF
            reg_file[1520] <= 8'h33
            reg_file[1521] <= 8'h43
            reg_file[1522] <= 8'hE5
            reg_file[1523] <= 8'h02
            reg_file[1524] <= 8'h13
            reg_file[1525] <= 8'h08
            reg_file[1526] <= 8'h03
            reg_file[1527] <= 8'h00
            reg_file[1528] <= 8'h63
            reg_file[1529] <= 8'h96
            reg_file[1530] <= 8'hF6
            reg_file[1531] <= 8'h00
            reg_file[1532] <= 8'h33
            reg_file[1533] <= 8'h65
            reg_file[1534] <= 8'hE5
            reg_file[1535] <= 8'h02
            reg_file[1536] <= 8'h33
            reg_file[1537] <= 8'h08
            reg_file[1538] <= 8'h65
            reg_file[1539] <= 8'h00
            reg_file[1540] <= 8'h33
            reg_file[1541] <= 8'h49
            reg_file[1542] <= 8'h98
            reg_file[1543] <= 8'h02
            reg_file[1544] <= 8'h33
            reg_file[1545] <= 8'h64
            reg_file[1546] <= 8'h98
            reg_file[1547] <= 8'h02
            reg_file[1548] <= 8'h63
            reg_file[1549] <= 8'h4C
            reg_file[1550] <= 8'h19
            reg_file[1551] <= 8'h07
            reg_file[1552] <= 8'h13
            reg_file[1553] <= 8'h05
            reg_file[1554] <= 8'h10
            reg_file[1555] <= 8'h00
            reg_file[1556] <= 8'hB3
            reg_file[1557] <= 8'h46
            reg_file[1558] <= 8'h19
            reg_file[1559] <= 8'h03
            reg_file[1560] <= 8'h63
            reg_file[1561] <= 8'h86
            reg_file[1562] <= 8'h06
            reg_file[1563] <= 8'h00
            reg_file[1564] <= 8'h13
            reg_file[1565] <= 8'h85
            reg_file[1566] <= 8'h06
            reg_file[1567] <= 8'h00
            reg_file[1568] <= 8'hB3
            reg_file[1569] <= 8'h66
            reg_file[1570] <= 8'h19
            reg_file[1571] <= 8'h03
            reg_file[1572] <= 8'h17
            reg_file[1573] <= 8'h17
            reg_file[1574] <= 8'h00
            reg_file[1575] <= 8'h00
            reg_file[1576] <= 8'h13
            reg_file[1577] <= 8'h07
            reg_file[1578] <= 8'hC7
            reg_file[1579] <= 8'hE1
            reg_file[1580] <= 8'h23
            reg_file[1581] <= 8'h24
            reg_file[1582] <= 8'hB1
            reg_file[1583] <= 8'h00
            reg_file[1584] <= 8'h23
            reg_file[1585] <= 8'h26
            reg_file[1586] <= 8'hC1
            reg_file[1587] <= 8'h00
            reg_file[1588] <= 8'h23
            reg_file[1589] <= 8'h2A
            reg_file[1590] <= 8'hA1
            reg_file[1591] <= 8'h00
            reg_file[1592] <= 8'h23
            reg_file[1593] <= 8'h2C
            reg_file[1594] <= 8'hD1
            reg_file[1595] <= 8'h00
            reg_file[1596] <= 8'h23
            reg_file[1597] <= 8'h2E
            reg_file[1598] <= 8'h01
            reg_file[1599] <= 8'h00
            reg_file[1600] <= 8'h33
            reg_file[1601] <= 8'h03
            reg_file[1602] <= 8'hF3
            reg_file[1603] <= 8'h02
            reg_file[1604] <= 8'h93
            reg_file[1605] <= 8'h97
            reg_file[1606] <= 8'h27
            reg_file[1607] <= 8'h00
            reg_file[1608] <= 8'hB3
            reg_file[1609] <= 8'h07
            reg_file[1610] <= 8'hF7
            reg_file[1611] <= 8'h00
            reg_file[1612] <= 8'h13
            reg_file[1613] <= 8'h07
            reg_file[1614] <= 8'h81
            reg_file[1615] <= 8'h00
            reg_file[1616] <= 8'h23
            reg_file[1617] <= 8'hA0
            reg_file[1618] <= 8'hE7
            reg_file[1619] <= 8'h00
            reg_file[1620] <= 8'h23
            reg_file[1621] <= 8'h28
            reg_file[1622] <= 8'h61
            reg_file[1623] <= 8'h00
            reg_file[1624] <= 8'h63
            reg_file[1625] <= 8'h4C
            reg_file[1626] <= 8'h20
            reg_file[1627] <= 8'h03
            reg_file[1628] <= 8'h63
            reg_file[1629] <= 8'h16
            reg_file[1630] <= 8'h04
            reg_file[1631] <= 8'h06
            reg_file[1632] <= 8'h83
            reg_file[1633] <= 8'h20
            reg_file[1634] <= 8'hC1
            reg_file[1635] <= 8'h02
            reg_file[1636] <= 8'h03
            reg_file[1637] <= 8'h24
            reg_file[1638] <= 8'h81
            reg_file[1639] <= 8'h02
            reg_file[1640] <= 8'h83
            reg_file[1641] <= 8'h24
            reg_file[1642] <= 8'h41
            reg_file[1643] <= 8'h02
            reg_file[1644] <= 8'h03
            reg_file[1645] <= 8'h29
            reg_file[1646] <= 8'h01
            reg_file[1647] <= 8'h02
            reg_file[1648] <= 8'h13
            reg_file[1649] <= 8'h01
            reg_file[1650] <= 8'h01
            reg_file[1651] <= 8'h03
            reg_file[1652] <= 8'h67
            reg_file[1653] <= 8'h80
            reg_file[1654] <= 8'h00
            reg_file[1655] <= 8'h00
            reg_file[1656] <= 8'h13
            reg_file[1657] <= 8'h87
            reg_file[1658] <= 8'h06
            reg_file[1659] <= 8'h00
            reg_file[1660] <= 8'hE3
            reg_file[1661] <= 8'hC8
            reg_file[1662] <= 8'hE7
            reg_file[1663] <= 8'hF6
            reg_file[1664] <= 8'h6F
            reg_file[1665] <= 8'hF0
            reg_file[1666] <= 8'h1F
            reg_file[1667] <= 8'hFE
            reg_file[1668] <= 8'h93
            reg_file[1669] <= 8'h06
            reg_file[1670] <= 8'h00
            reg_file[1671] <= 8'h00
            reg_file[1672] <= 8'h13
            reg_file[1673] <= 8'h05
            reg_file[1674] <= 8'h10
            reg_file[1675] <= 8'h00
            reg_file[1676] <= 8'h6F
            reg_file[1677] <= 8'hF0
            reg_file[1678] <= 8'h9F
            reg_file[1679] <= 8'hF9
            reg_file[1680] <= 8'h93
            reg_file[1681] <= 8'h07
            reg_file[1682] <= 8'h09
            reg_file[1683] <= 8'h00
            reg_file[1684] <= 8'h63
            reg_file[1685] <= 8'hD4
            reg_file[1686] <= 8'h28
            reg_file[1687] <= 8'h01
            reg_file[1688] <= 8'h93
            reg_file[1689] <= 8'h87
            reg_file[1690] <= 8'h08
            reg_file[1691] <= 8'h00
            reg_file[1692] <= 8'h23
            reg_file[1693] <= 8'h2E
            reg_file[1694] <= 8'hF1
            reg_file[1695] <= 8'h00
            reg_file[1696] <= 8'h17
            reg_file[1697] <= 8'h07
            reg_file[1698] <= 8'h00
            reg_file[1699] <= 8'h00
            reg_file[1700] <= 8'h13
            reg_file[1701] <= 8'h07
            reg_file[1702] <= 8'h07
            reg_file[1703] <= 8'hCD
            reg_file[1704] <= 8'h6B
            reg_file[1705] <= 8'h90
            reg_file[1706] <= 8'hE7
            reg_file[1707] <= 8'h00
            reg_file[1708] <= 8'h93
            reg_file[1709] <= 8'h07
            reg_file[1710] <= 8'hF0
            reg_file[1711] <= 8'hFF
            reg_file[1712] <= 8'h6B
            reg_file[1713] <= 8'h80
            reg_file[1714] <= 8'h07
            reg_file[1715] <= 8'h00
            reg_file[1716] <= 8'hEF
            reg_file[1717] <= 8'hF0
            reg_file[1718] <= 8'h9F
            reg_file[1719] <= 8'hBD
            reg_file[1720] <= 8'hF3
            reg_file[1721] <= 8'h27
            reg_file[1722] <= 8'h30
            reg_file[1723] <= 8'hCC
            reg_file[1724] <= 8'h93
            reg_file[1725] <= 8'hB7
            reg_file[1726] <= 8'h17
            reg_file[1727] <= 8'h00
            reg_file[1728] <= 8'h6B
            reg_file[1729] <= 8'h80
            reg_file[1730] <= 8'h07
            reg_file[1731] <= 8'h00
            reg_file[1732] <= 8'hE3
            reg_file[1733] <= 8'h0E
            reg_file[1734] <= 8'h04
            reg_file[1735] <= 8'hF8
            reg_file[1736] <= 8'hB3
            reg_file[1737] <= 8'h04
            reg_file[1738] <= 8'h99
            reg_file[1739] <= 8'h02
            reg_file[1740] <= 8'h13
            reg_file[1741] <= 8'h09
            reg_file[1742] <= 8'h10
            reg_file[1743] <= 8'h00
            reg_file[1744] <= 8'h33
            reg_file[1745] <= 8'h18
            reg_file[1746] <= 8'h89
            reg_file[1747] <= 8'h00
            reg_file[1748] <= 8'h13
            reg_file[1749] <= 8'h08
            reg_file[1750] <= 8'hF8
            reg_file[1751] <= 8'hFF
            reg_file[1752] <= 8'h23
            reg_file[1753] <= 8'h28
            reg_file[1754] <= 8'h91
            reg_file[1755] <= 8'h00
            reg_file[1756] <= 8'h6B
            reg_file[1757] <= 8'h00
            reg_file[1758] <= 8'h08
            reg_file[1759] <= 8'h00
            reg_file[1760] <= 8'hEF
            reg_file[1761] <= 8'hF0
            reg_file[1762] <= 8'h1F
            reg_file[1763] <= 8'hC6
            reg_file[1764] <= 8'h6B
            reg_file[1765] <= 8'h00
            reg_file[1766] <= 8'h09
            reg_file[1767] <= 8'h00
            reg_file[1768] <= 8'h83
            reg_file[1769] <= 8'h20
            reg_file[1770] <= 8'hC1
            reg_file[1771] <= 8'h02
            reg_file[1772] <= 8'h03
            reg_file[1773] <= 8'h24
            reg_file[1774] <= 8'h81
            reg_file[1775] <= 8'h02
            reg_file[1776] <= 8'h83
            reg_file[1777] <= 8'h24
            reg_file[1778] <= 8'h41
            reg_file[1779] <= 8'h02
            reg_file[1780] <= 8'h03
            reg_file[1781] <= 8'h29
            reg_file[1782] <= 8'h01
            reg_file[1783] <= 8'h02
            reg_file[1784] <= 8'h13
            reg_file[1785] <= 8'h01
            reg_file[1786] <= 8'h01
            reg_file[1787] <= 8'h03
            reg_file[1788] <= 8'h67
            reg_file[1789] <= 8'h80
            reg_file[1790] <= 8'h00
            reg_file[1791] <= 8'h00
            reg_file[1792] <= 8'h13
            reg_file[1793] <= 8'h01
            reg_file[1794] <= 8'h01
            reg_file[1795] <= 8'hFD
            reg_file[1796] <= 8'h23
            reg_file[1797] <= 8'h26
            reg_file[1798] <= 8'h11
            reg_file[1799] <= 8'h02
            reg_file[1800] <= 8'h23
            reg_file[1801] <= 8'h24
            reg_file[1802] <= 8'h81
            reg_file[1803] <= 8'h02
            reg_file[1804] <= 8'h23
            reg_file[1805] <= 8'h22
            reg_file[1806] <= 8'h91
            reg_file[1807] <= 8'h02
            reg_file[1808] <= 8'h23
            reg_file[1809] <= 8'h20
            reg_file[1810] <= 8'h21
            reg_file[1811] <= 8'h03
            reg_file[1812] <= 8'hF3
            reg_file[1813] <= 8'h28
            reg_file[1814] <= 8'h20
            reg_file[1815] <= 8'hFC
            reg_file[1816] <= 8'h73
            reg_file[1817] <= 8'h23
            reg_file[1818] <= 8'h10
            reg_file[1819] <= 8'hFC
            reg_file[1820] <= 8'hF3
            reg_file[1821] <= 8'h24
            reg_file[1822] <= 8'h00
            reg_file[1823] <= 8'hFC
            reg_file[1824] <= 8'hF3
            reg_file[1825] <= 8'h27
            reg_file[1826] <= 8'h50
            reg_file[1827] <= 8'hCC
            reg_file[1828] <= 8'h13
            reg_file[1829] <= 8'h07
            reg_file[1830] <= 8'hF0
            reg_file[1831] <= 8'h01
            reg_file[1832] <= 8'h63
            reg_file[1833] <= 8'h46
            reg_file[1834] <= 8'hF7
            reg_file[1835] <= 8'h0E
            reg_file[1836] <= 8'h03
            reg_file[1837] <= 8'h2E
            reg_file[1838] <= 8'h05
            reg_file[1839] <= 8'h00
            reg_file[1840] <= 8'h83
            reg_file[1841] <= 8'h26
            reg_file[1842] <= 8'h45
            reg_file[1843] <= 8'h00
            reg_file[1844] <= 8'h03
            reg_file[1845] <= 8'h28
            reg_file[1846] <= 8'h85
            reg_file[1847] <= 8'h00
            reg_file[1848] <= 8'hB3
            reg_file[1849] <= 8'h0E
            reg_file[1850] <= 8'h93
            reg_file[1851] <= 8'h02
            reg_file[1852] <= 8'h13
            reg_file[1853] <= 8'h07
            reg_file[1854] <= 8'h10
            reg_file[1855] <= 8'h00
            reg_file[1856] <= 8'hB3
            reg_file[1857] <= 8'h06
            reg_file[1858] <= 8'hDE
            reg_file[1859] <= 8'h02
            reg_file[1860] <= 8'h33
            reg_file[1861] <= 8'h88
            reg_file[1862] <= 8'h06
            reg_file[1863] <= 8'h03
            reg_file[1864] <= 8'h63
            reg_file[1865] <= 8'hD4
            reg_file[1866] <= 8'h0E
            reg_file[1867] <= 8'h01
            reg_file[1868] <= 8'h33
            reg_file[1869] <= 8'h47
            reg_file[1870] <= 8'hD8
            reg_file[1871] <= 8'h03
            reg_file[1872] <= 8'h63
            reg_file[1873] <= 8'hCE
            reg_file[1874] <= 8'hE8
            reg_file[1875] <= 8'h0C
            reg_file[1876] <= 8'h63
            reg_file[1877] <= 8'hD0
            reg_file[1878] <= 8'hE7
            reg_file[1879] <= 8'h0C
            reg_file[1880] <= 8'h93
            reg_file[1881] <= 8'h88
            reg_file[1882] <= 8'hF8
            reg_file[1883] <= 8'hFF
            reg_file[1884] <= 8'h33
            reg_file[1885] <= 8'h4F
            reg_file[1886] <= 8'hE8
            reg_file[1887] <= 8'h02
            reg_file[1888] <= 8'h13
            reg_file[1889] <= 8'h04
            reg_file[1890] <= 8'h0F
            reg_file[1891] <= 8'h00
            reg_file[1892] <= 8'h63
            reg_file[1893] <= 8'h96
            reg_file[1894] <= 8'hF8
            reg_file[1895] <= 8'h00
            reg_file[1896] <= 8'h33
            reg_file[1897] <= 8'h67
            reg_file[1898] <= 8'hE8
            reg_file[1899] <= 8'h02
            reg_file[1900] <= 8'h33
            reg_file[1901] <= 8'h04
            reg_file[1902] <= 8'hE7
            reg_file[1903] <= 8'h01
            reg_file[1904] <= 8'h33
            reg_file[1905] <= 8'h49
            reg_file[1906] <= 8'h94
            reg_file[1907] <= 8'h02
            reg_file[1908] <= 8'h33
            reg_file[1909] <= 8'h64
            reg_file[1910] <= 8'h94
            reg_file[1911] <= 8'h02
            reg_file[1912] <= 8'h63
            reg_file[1913] <= 8'h40
            reg_file[1914] <= 8'h69
            reg_file[1915] <= 8'h0C
            reg_file[1916] <= 8'h93
            reg_file[1917] <= 8'h02
            reg_file[1918] <= 8'h10
            reg_file[1919] <= 8'h00
            reg_file[1920] <= 8'hB3
            reg_file[1921] <= 8'h4F
            reg_file[1922] <= 8'h69
            reg_file[1923] <= 8'h02
            reg_file[1924] <= 8'h63
            reg_file[1925] <= 8'h86
            reg_file[1926] <= 8'h0F
            reg_file[1927] <= 8'h00
            reg_file[1928] <= 8'h93
            reg_file[1929] <= 8'h82
            reg_file[1930] <= 8'h0F
            reg_file[1931] <= 8'h00
            reg_file[1932] <= 8'hB3
            reg_file[1933] <= 8'h6F
            reg_file[1934] <= 8'h69
            reg_file[1935] <= 8'h02
            reg_file[1936] <= 8'hD3
            reg_file[1937] <= 8'hF7
            reg_file[1938] <= 8'h06
            reg_file[1939] <= 8'hD0
            reg_file[1940] <= 8'h93
            reg_file[1941] <= 8'h08
            reg_file[1942] <= 8'hFE
            reg_file[1943] <= 8'hFF
            reg_file[1944] <= 8'h93
            reg_file[1945] <= 8'h8E
            reg_file[1946] <= 8'hF6
            reg_file[1947] <= 8'hFF
            reg_file[1948] <= 8'h53
            reg_file[1949] <= 8'h88
            reg_file[1950] <= 8'h07
            reg_file[1951] <= 8'hE0
            reg_file[1952] <= 8'hD3
            reg_file[1953] <= 8'h77
            reg_file[1954] <= 8'h0E
            reg_file[1955] <= 8'hD0
            reg_file[1956] <= 8'hB3
            reg_file[1957] <= 8'hF6
            reg_file[1958] <= 8'hDE
            reg_file[1959] <= 8'h00
            reg_file[1960] <= 8'h33
            reg_file[1961] <= 8'hFE
            reg_file[1962] <= 8'hC8
            reg_file[1963] <= 8'h01
            reg_file[1964] <= 8'h53
            reg_file[1965] <= 8'h87
            reg_file[1966] <= 8'h07
            reg_file[1967] <= 8'hE0
            reg_file[1968] <= 8'h13
            reg_file[1969] <= 8'h58
            reg_file[1970] <= 8'h78
            reg_file[1971] <= 8'h41
            reg_file[1972] <= 8'h97
            reg_file[1973] <= 8'h18
            reg_file[1974] <= 8'h00
            reg_file[1975] <= 8'h00
            reg_file[1976] <= 8'h93
            reg_file[1977] <= 8'h88
            reg_file[1978] <= 8'hC8
            reg_file[1979] <= 8'hC8
            reg_file[1980] <= 8'h13
            reg_file[1981] <= 8'h57
            reg_file[1982] <= 8'h77
            reg_file[1983] <= 8'h41
            reg_file[1984] <= 8'h93
            reg_file[1985] <= 8'hB6
            reg_file[1986] <= 8'h16
            reg_file[1987] <= 8'h00
            reg_file[1988] <= 8'h13
            reg_file[1989] <= 8'h3E
            reg_file[1990] <= 8'h1E
            reg_file[1991] <= 8'h00
            reg_file[1992] <= 8'h13
            reg_file[1993] <= 8'h08
            reg_file[1994] <= 8'h18
            reg_file[1995] <= 8'hF8
            reg_file[1996] <= 8'h13
            reg_file[1997] <= 8'h07
            reg_file[1998] <= 8'h17
            reg_file[1999] <= 8'hF8
            reg_file[2000] <= 8'h23
            reg_file[2001] <= 8'h20
            reg_file[2002] <= 8'hA1
            reg_file[2003] <= 8'h00
            reg_file[2004] <= 8'h23
            reg_file[2005] <= 8'h22
            reg_file[2006] <= 8'hB1
            reg_file[2007] <= 8'h00
            reg_file[2008] <= 8'h23
            reg_file[2009] <= 8'h24
            reg_file[2010] <= 8'hC1
            reg_file[2011] <= 8'h00
            reg_file[2012] <= 8'h23
            reg_file[2013] <= 8'h28
            reg_file[2014] <= 8'h51
            reg_file[2015] <= 8'h00
            reg_file[2016] <= 8'h23
            reg_file[2017] <= 8'h2A
            reg_file[2018] <= 8'hF1
            reg_file[2019] <= 8'h01
            reg_file[2020] <= 8'h23
            reg_file[2021] <= 8'h2C
            reg_file[2022] <= 8'h01
            reg_file[2023] <= 8'h00
            reg_file[2024] <= 8'h23
            reg_file[2025] <= 8'h0E
            reg_file[2026] <= 8'hD1
            reg_file[2027] <= 8'h00
            reg_file[2028] <= 8'hA3
            reg_file[2029] <= 8'h0E
            reg_file[2030] <= 8'hC1
            reg_file[2031] <= 8'h01
            reg_file[2032] <= 8'h23
            reg_file[2033] <= 8'h0F
            reg_file[2034] <= 8'h01
            reg_file[2035] <= 8'h01
            reg_file[2036] <= 8'hA3
            reg_file[2037] <= 8'h0F
            reg_file[2038] <= 8'hE1
            reg_file[2039] <= 8'h00
            reg_file[2040] <= 8'h33
            reg_file[2041] <= 8'h0F
            reg_file[2042] <= 8'hFF
            reg_file[2043] <= 8'h02
            reg_file[2044] <= 8'h93
            reg_file[2045] <= 8'h97
            reg_file[2046] <= 8'h27
            reg_file[2047] <= 8'h00
            reg_file[2048] <= 8'hB3
            reg_file[2049] <= 8'h87
            reg_file[2050] <= 8'hF8
            reg_file[2051] <= 8'h00
            reg_file[2052] <= 8'h23
            reg_file[2053] <= 8'hA0
            reg_file[2054] <= 8'h27
            reg_file[2055] <= 8'h00
            reg_file[2056] <= 8'h23
            reg_file[2057] <= 8'h26
            reg_file[2058] <= 8'hE1
            reg_file[2059] <= 8'h01
            reg_file[2060] <= 8'h63
            reg_file[2061] <= 8'h4C
            reg_file[2062] <= 8'h20
            reg_file[2063] <= 8'h03
            reg_file[2064] <= 8'h63
            reg_file[2065] <= 8'h16
            reg_file[2066] <= 8'h04
            reg_file[2067] <= 8'h06
            reg_file[2068] <= 8'h83
            reg_file[2069] <= 8'h20
            reg_file[2070] <= 8'hC1
            reg_file[2071] <= 8'h02
            reg_file[2072] <= 8'h03
            reg_file[2073] <= 8'h24
            reg_file[2074] <= 8'h81
            reg_file[2075] <= 8'h02
            reg_file[2076] <= 8'h83
            reg_file[2077] <= 8'h24
            reg_file[2078] <= 8'h41
            reg_file[2079] <= 8'h02
            reg_file[2080] <= 8'h03
            reg_file[2081] <= 8'h29
            reg_file[2082] <= 8'h01
            reg_file[2083] <= 8'h02
            reg_file[2084] <= 8'h13
            reg_file[2085] <= 8'h01
            reg_file[2086] <= 8'h01
            reg_file[2087] <= 8'h03
            reg_file[2088] <= 8'h67
            reg_file[2089] <= 8'h80
            reg_file[2090] <= 8'h00
            reg_file[2091] <= 8'h00
            reg_file[2092] <= 8'h13
            reg_file[2093] <= 8'h87
            reg_file[2094] <= 8'h08
            reg_file[2095] <= 8'h00
            reg_file[2096] <= 8'hE3
            reg_file[2097] <= 8'hC4
            reg_file[2098] <= 8'hE7
            reg_file[2099] <= 8'hF2
            reg_file[2100] <= 8'h6F
            reg_file[2101] <= 8'hF0
            reg_file[2102] <= 8'h1F
            reg_file[2103] <= 8'hFE
            reg_file[2104] <= 8'h93
            reg_file[2105] <= 8'h0F
            reg_file[2106] <= 8'h00
            reg_file[2107] <= 8'h00
            reg_file[2108] <= 8'h93
            reg_file[2109] <= 8'h02
            reg_file[2110] <= 8'h10
            reg_file[2111] <= 8'h00
            reg_file[2112] <= 8'h6F
            reg_file[2113] <= 8'hF0
            reg_file[2114] <= 8'h1F
            reg_file[2115] <= 8'hF5
            reg_file[2116] <= 8'h93
            reg_file[2117] <= 8'h07
            reg_file[2118] <= 8'h09
            reg_file[2119] <= 8'h00
            reg_file[2120] <= 8'h63
            reg_file[2121] <= 8'h54
            reg_file[2122] <= 8'h23
            reg_file[2123] <= 8'h01
            reg_file[2124] <= 8'h93
            reg_file[2125] <= 8'h07
            reg_file[2126] <= 8'h03
            reg_file[2127] <= 8'h00
            reg_file[2128] <= 8'h23
            reg_file[2129] <= 8'h2C
            reg_file[2130] <= 8'hF1
            reg_file[2131] <= 8'h00
            reg_file[2132] <= 8'h17
            reg_file[2133] <= 8'h07
            reg_file[2134] <= 8'h00
            reg_file[2135] <= 8'h00
            reg_file[2136] <= 8'h13
            reg_file[2137] <= 8'h07
            reg_file[2138] <= 8'h87
            reg_file[2139] <= 8'hD2
            reg_file[2140] <= 8'h6B
            reg_file[2141] <= 8'h90
            reg_file[2142] <= 8'hE7
            reg_file[2143] <= 8'h00
            reg_file[2144] <= 8'h93
            reg_file[2145] <= 8'h07
            reg_file[2146] <= 8'hF0
            reg_file[2147] <= 8'hFF
            reg_file[2148] <= 8'h6B
            reg_file[2149] <= 8'h80
            reg_file[2150] <= 8'h07
            reg_file[2151] <= 8'h00
            reg_file[2152] <= 8'hEF
            reg_file[2153] <= 8'hF0
            reg_file[2154] <= 8'h5F
            reg_file[2155] <= 8'hB3
            reg_file[2156] <= 8'hF3
            reg_file[2157] <= 8'h27
            reg_file[2158] <= 8'h30
            reg_file[2159] <= 8'hCC
            reg_file[2160] <= 8'h93
            reg_file[2161] <= 8'hB7
            reg_file[2162] <= 8'h17
            reg_file[2163] <= 8'h00
            reg_file[2164] <= 8'h6B
            reg_file[2165] <= 8'h80
            reg_file[2166] <= 8'h07
            reg_file[2167] <= 8'h00
            reg_file[2168] <= 8'hE3
            reg_file[2169] <= 8'h0E
            reg_file[2170] <= 8'h04
            reg_file[2171] <= 8'hF8
            reg_file[2172] <= 8'hB3
            reg_file[2173] <= 8'h04
            reg_file[2174] <= 8'h99
            reg_file[2175] <= 8'h02
            reg_file[2176] <= 8'h13
            reg_file[2177] <= 8'h09
            reg_file[2178] <= 8'h10
            reg_file[2179] <= 8'h00
            reg_file[2180] <= 8'h33
            reg_file[2181] <= 8'h14
            reg_file[2182] <= 8'h89
            reg_file[2183] <= 8'h00
            reg_file[2184] <= 8'h13
            reg_file[2185] <= 8'h04
            reg_file[2186] <= 8'hF4
            reg_file[2187] <= 8'hFF
            reg_file[2188] <= 8'h23
            reg_file[2189] <= 8'h26
            reg_file[2190] <= 8'h91
            reg_file[2191] <= 8'h00
            reg_file[2192] <= 8'h6B
            reg_file[2193] <= 8'h00
            reg_file[2194] <= 8'h04
            reg_file[2195] <= 8'h00
            reg_file[2196] <= 8'hEF
            reg_file[2197] <= 8'hF0
            reg_file[2198] <= 8'h5F
            reg_file[2199] <= 8'hC4
            reg_file[2200] <= 8'h6B
            reg_file[2201] <= 8'h00
            reg_file[2202] <= 8'h09
            reg_file[2203] <= 8'h00
            reg_file[2204] <= 8'h83
            reg_file[2205] <= 8'h20
            reg_file[2206] <= 8'hC1
            reg_file[2207] <= 8'h02
            reg_file[2208] <= 8'h03
            reg_file[2209] <= 8'h24
            reg_file[2210] <= 8'h81
            reg_file[2211] <= 8'h02
            reg_file[2212] <= 8'h83
            reg_file[2213] <= 8'h24
            reg_file[2214] <= 8'h41
            reg_file[2215] <= 8'h02
            reg_file[2216] <= 8'h03
            reg_file[2217] <= 8'h29
            reg_file[2218] <= 8'h01
            reg_file[2219] <= 8'h02
            reg_file[2220] <= 8'h13
            reg_file[2221] <= 8'h01
            reg_file[2222] <= 8'h01
            reg_file[2223] <= 8'h03
            reg_file[2224] <= 8'h67
            reg_file[2225] <= 8'h80
            reg_file[2226] <= 8'h00
            reg_file[2227] <= 8'h00
            reg_file[2228] <= 8'h13
            reg_file[2229] <= 8'h01
            reg_file[2230] <= 8'h81
            reg_file[2231] <= 8'hFE
            reg_file[2232] <= 8'h23
            reg_file[2233] <= 8'h2A
            reg_file[2234] <= 8'h11
            reg_file[2235] <= 8'h00
            reg_file[2236] <= 8'h23
            reg_file[2237] <= 8'h28
            reg_file[2238] <= 8'h41
            reg_file[2239] <= 8'h01
            reg_file[2240] <= 8'h23
            reg_file[2241] <= 8'h26
            reg_file[2242] <= 8'h31
            reg_file[2243] <= 8'h01
            reg_file[2244] <= 8'h23
            reg_file[2245] <= 8'h24
            reg_file[2246] <= 8'h21
            reg_file[2247] <= 8'h01
            reg_file[2248] <= 8'h23
            reg_file[2249] <= 8'h22
            reg_file[2250] <= 8'h91
            reg_file[2251] <= 8'h00
            reg_file[2252] <= 8'h23
            reg_file[2253] <= 8'h20
            reg_file[2254] <= 8'h81
            reg_file[2255] <= 8'h00
            reg_file[2256] <= 8'h13
            reg_file[2257] <= 8'h0A
            reg_file[2258] <= 8'h05
            reg_file[2259] <= 8'h00
            reg_file[2260] <= 8'h93
            reg_file[2261] <= 8'h89
            reg_file[2262] <= 8'h05
            reg_file[2263] <= 8'h00
            reg_file[2264] <= 8'h73
            reg_file[2265] <= 8'h29
            reg_file[2266] <= 8'h00
            reg_file[2267] <= 8'hFC
            reg_file[2268] <= 8'hF3
            reg_file[2269] <= 8'h24
            reg_file[2270] <= 8'h00
            reg_file[2271] <= 8'hCC
            reg_file[2272] <= 8'h13
            reg_file[2273] <= 8'h04
            reg_file[2274] <= 8'h00
            reg_file[2275] <= 8'h00
            reg_file[2276] <= 8'hB3
            reg_file[2277] <= 8'h02
            reg_file[2278] <= 8'h94
            reg_file[2279] <= 8'h40
            reg_file[2280] <= 8'h13
            reg_file[2281] <= 8'hB3
            reg_file[2282] <= 8'h12
            reg_file[2283] <= 8'h00
            reg_file[2284] <= 8'h6B
            reg_file[2285] <= 8'h20
            reg_file[2286] <= 8'h03
            reg_file[2287] <= 8'h00
            reg_file[2288] <= 8'h63
            reg_file[2289] <= 8'h96
            reg_file[2290] <= 8'h02
            reg_file[2291] <= 8'h00
            reg_file[2292] <= 8'h13
            reg_file[2293] <= 8'h85
            reg_file[2294] <= 8'h09
            reg_file[2295] <= 8'h00
            reg_file[2296] <= 8'hE7
            reg_file[2297] <= 8'h00
            reg_file[2298] <= 8'h0A
            reg_file[2299] <= 8'h00
            reg_file[2300] <= 8'h6B
            reg_file[2301] <= 8'h30
            reg_file[2302] <= 8'h00
            reg_file[2303] <= 8'h00
            reg_file[2304] <= 8'h13
            reg_file[2305] <= 8'h04
            reg_file[2306] <= 8'h14
            reg_file[2307] <= 8'h00
            reg_file[2308] <= 8'hE3
            reg_file[2309] <= 8'h40
            reg_file[2310] <= 8'h24
            reg_file[2311] <= 8'hFF
            reg_file[2312] <= 8'h83
            reg_file[2313] <= 8'h20
            reg_file[2314] <= 8'h41
            reg_file[2315] <= 8'h01
            reg_file[2316] <= 8'h03
            reg_file[2317] <= 8'h2A
            reg_file[2318] <= 8'h01
            reg_file[2319] <= 8'h01
            reg_file[2320] <= 8'h83
            reg_file[2321] <= 8'h29
            reg_file[2322] <= 8'hC1
            reg_file[2323] <= 8'h00
            reg_file[2324] <= 8'h03
            reg_file[2325] <= 8'h29
            reg_file[2326] <= 8'h81
            reg_file[2327] <= 8'h00
            reg_file[2328] <= 8'h83
            reg_file[2329] <= 8'h24
            reg_file[2330] <= 8'h41
            reg_file[2331] <= 8'h00
            reg_file[2332] <= 8'h03
            reg_file[2333] <= 8'h24
            reg_file[2334] <= 8'h01
            reg_file[2335] <= 8'h00
            reg_file[2336] <= 8'h13
            reg_file[2337] <= 8'h01
            reg_file[2338] <= 8'h81
            reg_file[2339] <= 8'h01
            reg_file[2340] <= 8'h67
            reg_file[2341] <= 8'h80
            reg_file[2342] <= 8'h00
            reg_file[2343] <= 8'h00
            reg_file[2344] <= 8'h13
            reg_file[2345] <= 8'h05
            reg_file[2346] <= 8'hF0
            reg_file[2347] <= 8'hFF
            reg_file[2348] <= 8'h67
            reg_file[2349] <= 8'h80
            reg_file[2350] <= 8'h00
            reg_file[2351] <= 8'h00
            reg_file[2352] <= 8'h13
            reg_file[2353] <= 8'h05
            reg_file[2354] <= 8'hF0
            reg_file[2355] <= 8'hFF
            reg_file[2356] <= 8'h67
            reg_file[2357] <= 8'h80
            reg_file[2358] <= 8'h00
            reg_file[2359] <= 8'h00
            reg_file[2360] <= 8'h13
            reg_file[2361] <= 8'h05
            reg_file[2362] <= 8'hF0
            reg_file[2363] <= 8'hFF
            reg_file[2364] <= 8'h67
            reg_file[2365] <= 8'h80
            reg_file[2366] <= 8'h00
            reg_file[2367] <= 8'h00
            reg_file[2368] <= 8'h13
            reg_file[2369] <= 8'h05
            reg_file[2370] <= 8'hF0
            reg_file[2371] <= 8'hFF
            reg_file[2372] <= 8'h67
            reg_file[2373] <= 8'h80
            reg_file[2374] <= 8'h00
            reg_file[2375] <= 8'h00
            reg_file[2376] <= 8'h13
            reg_file[2377] <= 8'h05
            reg_file[2378] <= 8'hF0
            reg_file[2379] <= 8'hFF
            reg_file[2380] <= 8'h67
            reg_file[2381] <= 8'h80
            reg_file[2382] <= 8'h00
            reg_file[2383] <= 8'h00
            reg_file[2384] <= 8'h13
            reg_file[2385] <= 8'h05
            reg_file[2386] <= 8'hF0
            reg_file[2387] <= 8'hFF
            reg_file[2388] <= 8'h67
            reg_file[2389] <= 8'h80
            reg_file[2390] <= 8'h00
            reg_file[2391] <= 8'h00
            reg_file[2392] <= 8'h13
            reg_file[2393] <= 8'h05
            reg_file[2394] <= 8'h00
            reg_file[2395] <= 8'h00
            reg_file[2396] <= 8'h67
            reg_file[2397] <= 8'h80
            reg_file[2398] <= 8'h00
            reg_file[2399] <= 8'h00
            reg_file[2400] <= 8'h13
            reg_file[2401] <= 8'h05
            reg_file[2402] <= 8'hF0
            reg_file[2403] <= 8'hFF
            reg_file[2404] <= 8'h67
            reg_file[2405] <= 8'h80
            reg_file[2406] <= 8'h00
            reg_file[2407] <= 8'h00
            reg_file[2408] <= 8'h13
            reg_file[2409] <= 8'h05
            reg_file[2410] <= 8'hF0
            reg_file[2411] <= 8'hFF
            reg_file[2412] <= 8'h67
            reg_file[2413] <= 8'h80
            reg_file[2414] <= 8'h00
            reg_file[2415] <= 8'h00
            reg_file[2416] <= 8'h13
            reg_file[2417] <= 8'h05
            reg_file[2418] <= 8'hF0
            reg_file[2419] <= 8'hFF
            reg_file[2420] <= 8'h67
            reg_file[2421] <= 8'h80
            reg_file[2422] <= 8'h00
            reg_file[2423] <= 8'h00
            reg_file[2424] <= 8'h13
            reg_file[2425] <= 8'h05
            reg_file[2426] <= 8'hF0
            reg_file[2427] <= 8'hFF
            reg_file[2428] <= 8'h67
            reg_file[2429] <= 8'h80
            reg_file[2430] <= 8'h00
            reg_file[2431] <= 8'h00
            reg_file[2432] <= 8'h13
            reg_file[2433] <= 8'h05
            reg_file[2434] <= 8'hF0
            reg_file[2435] <= 8'hFF
            reg_file[2436] <= 8'h67
            reg_file[2437] <= 8'h80
            reg_file[2438] <= 8'h00
            reg_file[2439] <= 8'h00
            reg_file[2440] <= 8'h93
            reg_file[2441] <= 8'h05
            reg_file[2442] <= 8'h05
            reg_file[2443] <= 8'h00
            reg_file[2444] <= 8'h93
            reg_file[2445] <= 8'h06
            reg_file[2446] <= 8'h00
            reg_file[2447] <= 8'h00
            reg_file[2448] <= 8'h13
            reg_file[2449] <= 8'h06
            reg_file[2450] <= 8'h00
            reg_file[2451] <= 8'h00
            reg_file[2452] <= 8'h13
            reg_file[2453] <= 8'h05
            reg_file[2454] <= 8'h00
            reg_file[2455] <= 8'h00
            reg_file[2456] <= 8'h6F
            reg_file[2457] <= 8'h00
            reg_file[2458] <= 8'h00
            reg_file[2459] <= 8'h23
            reg_file[2460] <= 8'h13
            reg_file[2461] <= 8'h01
            reg_file[2462] <= 8'h01
            reg_file[2463] <= 8'hFF
            reg_file[2464] <= 8'h93
            reg_file[2465] <= 8'h05
            reg_file[2466] <= 8'h00
            reg_file[2467] <= 8'h00
            reg_file[2468] <= 8'h23
            reg_file[2469] <= 8'h24
            reg_file[2470] <= 8'h81
            reg_file[2471] <= 8'h00
            reg_file[2472] <= 8'h23
            reg_file[2473] <= 8'h26
            reg_file[2474] <= 8'h11
            reg_file[2475] <= 8'h00
            reg_file[2476] <= 8'h13
            reg_file[2477] <= 8'h04
            reg_file[2478] <= 8'h05
            reg_file[2479] <= 8'h00
            reg_file[2480] <= 8'hEF
            reg_file[2481] <= 8'h00
            reg_file[2482] <= 8'h40
            reg_file[2483] <= 8'h2B
            reg_file[2484] <= 8'hB7
            reg_file[2485] <= 8'h17
            reg_file[2486] <= 8'h00
            reg_file[2487] <= 8'h80
            reg_file[2488] <= 8'h03
            reg_file[2489] <= 8'hA5
            reg_file[2490] <= 8'h87
            reg_file[2491] <= 8'h43
            reg_file[2492] <= 8'h83
            reg_file[2493] <= 8'h27
            reg_file[2494] <= 8'hC5
            reg_file[2495] <= 8'h03
            reg_file[2496] <= 8'h63
            reg_file[2497] <= 8'h84
            reg_file[2498] <= 8'h07
            reg_file[2499] <= 8'h00
            reg_file[2500] <= 8'hE7
            reg_file[2501] <= 8'h80
            reg_file[2502] <= 8'h07
            reg_file[2503] <= 8'h00
            reg_file[2504] <= 8'h13
            reg_file[2505] <= 8'h05
            reg_file[2506] <= 8'h04
            reg_file[2507] <= 8'h00
            reg_file[2508] <= 8'hEF
            reg_file[2509] <= 8'hF0
            reg_file[2510] <= 8'h8F
            reg_file[2511] <= 8'hEC
            reg_file[2512] <= 8'hB3
            reg_file[2513] <= 8'hC7
            reg_file[2514] <= 8'hA5
            reg_file[2515] <= 8'h00
            reg_file[2516] <= 8'h93
            reg_file[2517] <= 8'hF7
            reg_file[2518] <= 8'h37
            reg_file[2519] <= 8'h00
            reg_file[2520] <= 8'hB3
            reg_file[2521] <= 8'h08
            reg_file[2522] <= 8'hC5
            reg_file[2523] <= 8'h00
            reg_file[2524] <= 8'h63
            reg_file[2525] <= 8'h92
            reg_file[2526] <= 8'h07
            reg_file[2527] <= 8'h06
            reg_file[2528] <= 8'h93
            reg_file[2529] <= 8'h07
            reg_file[2530] <= 8'h30
            reg_file[2531] <= 8'h00
            reg_file[2532] <= 8'h63
            reg_file[2533] <= 8'hFE
            reg_file[2534] <= 8'hC7
            reg_file[2535] <= 8'h04
            reg_file[2536] <= 8'h93
            reg_file[2537] <= 8'h77
            reg_file[2538] <= 8'h35
            reg_file[2539] <= 8'h00
            reg_file[2540] <= 8'h13
            reg_file[2541] <= 8'h07
            reg_file[2542] <= 8'h05
            reg_file[2543] <= 8'h00
            reg_file[2544] <= 8'h63
            reg_file[2545] <= 8'h98
            reg_file[2546] <= 8'h07
            reg_file[2547] <= 8'h06
            reg_file[2548] <= 8'h13
            reg_file[2549] <= 8'hF6
            reg_file[2550] <= 8'hC8
            reg_file[2551] <= 8'hFF
            reg_file[2552] <= 8'h93
            reg_file[2553] <= 8'h07
            reg_file[2554] <= 8'h06
            reg_file[2555] <= 8'hFE
            reg_file[2556] <= 8'h63
            reg_file[2557] <= 8'h6C
            reg_file[2558] <= 8'hF7
            reg_file[2559] <= 8'h08
            reg_file[2560] <= 8'h63
            reg_file[2561] <= 8'h7C
            reg_file[2562] <= 8'hC7
            reg_file[2563] <= 8'h02
            reg_file[2564] <= 8'h93
            reg_file[2565] <= 8'h86
            reg_file[2566] <= 8'h05
            reg_file[2567] <= 8'h00
            reg_file[2568] <= 8'h93
            reg_file[2569] <= 8'h07
            reg_file[2570] <= 8'h07
            reg_file[2571] <= 8'h00
            reg_file[2572] <= 8'h03
            reg_file[2573] <= 8'hA8
            reg_file[2574] <= 8'h06
            reg_file[2575] <= 8'h00
            reg_file[2576] <= 8'h93
            reg_file[2577] <= 8'h87
            reg_file[2578] <= 8'h47
            reg_file[2579] <= 8'h00
            reg_file[2580] <= 8'h93
            reg_file[2581] <= 8'h86
            reg_file[2582] <= 8'h46
            reg_file[2583] <= 8'h00
            reg_file[2584] <= 8'h23
            reg_file[2585] <= 8'hAE
            reg_file[2586] <= 8'h07
            reg_file[2587] <= 8'hFF
            reg_file[2588] <= 8'hE3
            reg_file[2589] <= 8'hE8
            reg_file[2590] <= 8'hC7
            reg_file[2591] <= 8'hFE
            reg_file[2592] <= 8'h93
            reg_file[2593] <= 8'h07
            reg_file[2594] <= 8'hF6
            reg_file[2595] <= 8'hFF
            reg_file[2596] <= 8'hB3
            reg_file[2597] <= 8'h87
            reg_file[2598] <= 8'hE7
            reg_file[2599] <= 8'h40
            reg_file[2600] <= 8'h93
            reg_file[2601] <= 8'hF7
            reg_file[2602] <= 8'hC7
            reg_file[2603] <= 8'hFF
            reg_file[2604] <= 8'h93
            reg_file[2605] <= 8'h87
            reg_file[2606] <= 8'h47
            reg_file[2607] <= 8'h00
            reg_file[2608] <= 8'h33
            reg_file[2609] <= 8'h07
            reg_file[2610] <= 8'hF7
            reg_file[2611] <= 8'h00
            reg_file[2612] <= 8'hB3
            reg_file[2613] <= 8'h85
            reg_file[2614] <= 8'hF5
            reg_file[2615] <= 8'h00
            reg_file[2616] <= 8'h63
            reg_file[2617] <= 8'h68
            reg_file[2618] <= 8'h17
            reg_file[2619] <= 8'h01
            reg_file[2620] <= 8'h67
            reg_file[2621] <= 8'h80
            reg_file[2622] <= 8'h00
            reg_file[2623] <= 8'h00
            reg_file[2624] <= 8'h13
            reg_file[2625] <= 8'h07
            reg_file[2626] <= 8'h05
            reg_file[2627] <= 8'h00
            reg_file[2628] <= 8'hE3
            reg_file[2629] <= 8'h7C
            reg_file[2630] <= 8'h15
            reg_file[2631] <= 8'hFF
            reg_file[2632] <= 8'h83
            reg_file[2633] <= 8'hC7
            reg_file[2634] <= 8'h05
            reg_file[2635] <= 8'h00
            reg_file[2636] <= 8'h13
            reg_file[2637] <= 8'h07
            reg_file[2638] <= 8'h17
            reg_file[2639] <= 8'h00
            reg_file[2640] <= 8'h93
            reg_file[2641] <= 8'h85
            reg_file[2642] <= 8'h15
            reg_file[2643] <= 8'h00
            reg_file[2644] <= 8'hA3
            reg_file[2645] <= 8'h0F
            reg_file[2646] <= 8'hF7
            reg_file[2647] <= 8'hFE
            reg_file[2648] <= 8'hE3
            reg_file[2649] <= 8'h68
            reg_file[2650] <= 8'h17
            reg_file[2651] <= 8'hFF
            reg_file[2652] <= 8'h67
            reg_file[2653] <= 8'h80
            reg_file[2654] <= 8'h00
            reg_file[2655] <= 8'h00
            reg_file[2656] <= 8'h83
            reg_file[2657] <= 8'hC6
            reg_file[2658] <= 8'h05
            reg_file[2659] <= 8'h00
            reg_file[2660] <= 8'h13
            reg_file[2661] <= 8'h07
            reg_file[2662] <= 8'h17
            reg_file[2663] <= 8'h00
            reg_file[2664] <= 8'h93
            reg_file[2665] <= 8'h77
            reg_file[2666] <= 8'h37
            reg_file[2667] <= 8'h00
            reg_file[2668] <= 8'hA3
            reg_file[2669] <= 8'h0F
            reg_file[2670] <= 8'hD7
            reg_file[2671] <= 8'hFE
            reg_file[2672] <= 8'h93
            reg_file[2673] <= 8'h85
            reg_file[2674] <= 8'h15
            reg_file[2675] <= 8'h00
            reg_file[2676] <= 8'hE3
            reg_file[2677] <= 8'h80
            reg_file[2678] <= 8'h07
            reg_file[2679] <= 8'hF8
            reg_file[2680] <= 8'h83
            reg_file[2681] <= 8'hC6
            reg_file[2682] <= 8'h05
            reg_file[2683] <= 8'h00
            reg_file[2684] <= 8'h13
            reg_file[2685] <= 8'h07
            reg_file[2686] <= 8'h17
            reg_file[2687] <= 8'h00
            reg_file[2688] <= 8'h93
            reg_file[2689] <= 8'h77
            reg_file[2690] <= 8'h37
            reg_file[2691] <= 8'h00
            reg_file[2692] <= 8'hA3
            reg_file[2693] <= 8'h0F
            reg_file[2694] <= 8'hD7
            reg_file[2695] <= 8'hFE
            reg_file[2696] <= 8'h93
            reg_file[2697] <= 8'h85
            reg_file[2698] <= 8'h15
            reg_file[2699] <= 8'h00
            reg_file[2700] <= 8'hE3
            reg_file[2701] <= 8'h9A
            reg_file[2702] <= 8'h07
            reg_file[2703] <= 8'hFC
            reg_file[2704] <= 8'h6F
            reg_file[2705] <= 8'hF0
            reg_file[2706] <= 8'h5F
            reg_file[2707] <= 8'hF6
            reg_file[2708] <= 8'h83
            reg_file[2709] <= 8'hA6
            reg_file[2710] <= 8'h45
            reg_file[2711] <= 8'h00
            reg_file[2712] <= 8'h83
            reg_file[2713] <= 8'hA2
            reg_file[2714] <= 8'h05
            reg_file[2715] <= 8'h00
            reg_file[2716] <= 8'h83
            reg_file[2717] <= 8'hAF
            reg_file[2718] <= 8'h85
            reg_file[2719] <= 8'h00
            reg_file[2720] <= 8'h03
            reg_file[2721] <= 8'hAF
            reg_file[2722] <= 8'hC5
            reg_file[2723] <= 8'h00
            reg_file[2724] <= 8'h83
            reg_file[2725] <= 8'hAE
            reg_file[2726] <= 8'h05
            reg_file[2727] <= 8'h01
            reg_file[2728] <= 8'h03
            reg_file[2729] <= 8'hAE
            reg_file[2730] <= 8'h45
            reg_file[2731] <= 8'h01
            reg_file[2732] <= 8'h03
            reg_file[2733] <= 8'hA3
            reg_file[2734] <= 8'h85
            reg_file[2735] <= 8'h01
            reg_file[2736] <= 8'h03
            reg_file[2737] <= 8'hA8
            reg_file[2738] <= 8'hC5
            reg_file[2739] <= 8'h01
            reg_file[2740] <= 8'h23
            reg_file[2741] <= 8'h22
            reg_file[2742] <= 8'hD7
            reg_file[2743] <= 8'h00
            reg_file[2744] <= 8'h83
            reg_file[2745] <= 8'hA6
            reg_file[2746] <= 8'h05
            reg_file[2747] <= 8'h02
            reg_file[2748] <= 8'h23
            reg_file[2749] <= 8'h20
            reg_file[2750] <= 8'h57
            reg_file[2751] <= 8'h00
            reg_file[2752] <= 8'h23
            reg_file[2753] <= 8'h24
            reg_file[2754] <= 8'hF7
            reg_file[2755] <= 8'h01
            reg_file[2756] <= 8'h23
            reg_file[2757] <= 8'h26
            reg_file[2758] <= 8'hE7
            reg_file[2759] <= 8'h01
            reg_file[2760] <= 8'h23
            reg_file[2761] <= 8'h28
            reg_file[2762] <= 8'hD7
            reg_file[2763] <= 8'h01
            reg_file[2764] <= 8'h23
            reg_file[2765] <= 8'h2A
            reg_file[2766] <= 8'hC7
            reg_file[2767] <= 8'h01
            reg_file[2768] <= 8'h23
            reg_file[2769] <= 8'h2C
            reg_file[2770] <= 8'h67
            reg_file[2771] <= 8'h00
            reg_file[2772] <= 8'h23
            reg_file[2773] <= 8'h2E
            reg_file[2774] <= 8'h07
            reg_file[2775] <= 8'h01
            reg_file[2776] <= 8'h23
            reg_file[2777] <= 8'h20
            reg_file[2778] <= 8'hD7
            reg_file[2779] <= 8'h02
            reg_file[2780] <= 8'h13
            reg_file[2781] <= 8'h07
            reg_file[2782] <= 8'h47
            reg_file[2783] <= 8'h02
            reg_file[2784] <= 8'h93
            reg_file[2785] <= 8'h85
            reg_file[2786] <= 8'h45
            reg_file[2787] <= 8'h02
            reg_file[2788] <= 8'hE3
            reg_file[2789] <= 8'h68
            reg_file[2790] <= 8'hF7
            reg_file[2791] <= 8'hFA
            reg_file[2792] <= 8'h6F
            reg_file[2793] <= 8'hF0
            reg_file[2794] <= 8'h9F
            reg_file[2795] <= 8'hF1
            reg_file[2796] <= 8'h13
            reg_file[2797] <= 8'h03
            reg_file[2798] <= 8'hF0
            reg_file[2799] <= 8'h00
            reg_file[2800] <= 8'h13
            reg_file[2801] <= 8'h07
            reg_file[2802] <= 8'h05
            reg_file[2803] <= 8'h00
            reg_file[2804] <= 8'h63
            reg_file[2805] <= 8'h7E
            reg_file[2806] <= 8'hC3
            reg_file[2807] <= 8'h02
            reg_file[2808] <= 8'h93
            reg_file[2809] <= 8'h77
            reg_file[2810] <= 8'hF7
            reg_file[2811] <= 8'h00
            reg_file[2812] <= 8'h63
            reg_file[2813] <= 8'h90
            reg_file[2814] <= 8'h07
            reg_file[2815] <= 8'h0A
            reg_file[2816] <= 8'h63
            reg_file[2817] <= 8'h92
            reg_file[2818] <= 8'h05
            reg_file[2819] <= 8'h08
            reg_file[2820] <= 8'h93
            reg_file[2821] <= 8'h76
            reg_file[2822] <= 8'h06
            reg_file[2823] <= 8'hFF
            reg_file[2824] <= 8'h13
            reg_file[2825] <= 8'h76
            reg_file[2826] <= 8'hF6
            reg_file[2827] <= 8'h00
            reg_file[2828] <= 8'hB3
            reg_file[2829] <= 8'h86
            reg_file[2830] <= 8'hE6
            reg_file[2831] <= 8'h00
            reg_file[2832] <= 8'h23
            reg_file[2833] <= 8'h20
            reg_file[2834] <= 8'hB7
            reg_file[2835] <= 8'h00
            reg_file[2836] <= 8'h23
            reg_file[2837] <= 8'h22
            reg_file[2838] <= 8'hB7
            reg_file[2839] <= 8'h00
            reg_file[2840] <= 8'h23
            reg_file[2841] <= 8'h24
            reg_file[2842] <= 8'hB7
            reg_file[2843] <= 8'h00
            reg_file[2844] <= 8'h23
            reg_file[2845] <= 8'h26
            reg_file[2846] <= 8'hB7
            reg_file[2847] <= 8'h00
            reg_file[2848] <= 8'h13
            reg_file[2849] <= 8'h07
            reg_file[2850] <= 8'h07
            reg_file[2851] <= 8'h01
            reg_file[2852] <= 8'hE3
            reg_file[2853] <= 8'h66
            reg_file[2854] <= 8'hD7
            reg_file[2855] <= 8'hFE
            reg_file[2856] <= 8'h63
            reg_file[2857] <= 8'h14
            reg_file[2858] <= 8'h06
            reg_file[2859] <= 8'h00
            reg_file[2860] <= 8'h67
            reg_file[2861] <= 8'h80
            reg_file[2862] <= 8'h00
            reg_file[2863] <= 8'h00
            reg_file[2864] <= 8'hB3
            reg_file[2865] <= 8'h06
            reg_file[2866] <= 8'hC3
            reg_file[2867] <= 8'h40
            reg_file[2868] <= 8'h93
            reg_file[2869] <= 8'h96
            reg_file[2870] <= 8'h26
            reg_file[2871] <= 8'h00
            reg_file[2872] <= 8'h97
            reg_file[2873] <= 8'h02
            reg_file[2874] <= 8'h00
            reg_file[2875] <= 8'h00
            reg_file[2876] <= 8'hB3
            reg_file[2877] <= 8'h86
            reg_file[2878] <= 8'h56
            reg_file[2879] <= 8'h00
            reg_file[2880] <= 8'h67
            reg_file[2881] <= 8'h80
            reg_file[2882] <= 8'hC6
            reg_file[2883] <= 8'h00
            reg_file[2884] <= 8'h23
            reg_file[2885] <= 8'h07
            reg_file[2886] <= 8'hB7
            reg_file[2887] <= 8'h00
            reg_file[2888] <= 8'hA3
            reg_file[2889] <= 8'h06
            reg_file[2890] <= 8'hB7
            reg_file[2891] <= 8'h00
            reg_file[2892] <= 8'h23
            reg_file[2893] <= 8'h06
            reg_file[2894] <= 8'hB7
            reg_file[2895] <= 8'h00
            reg_file[2896] <= 8'hA3
            reg_file[2897] <= 8'h05
            reg_file[2898] <= 8'hB7
            reg_file[2899] <= 8'h00
            reg_file[2900] <= 8'h23
            reg_file[2901] <= 8'h05
            reg_file[2902] <= 8'hB7
            reg_file[2903] <= 8'h00
            reg_file[2904] <= 8'hA3
            reg_file[2905] <= 8'h04
            reg_file[2906] <= 8'hB7
            reg_file[2907] <= 8'h00
            reg_file[2908] <= 8'h23
            reg_file[2909] <= 8'h04
            reg_file[2910] <= 8'hB7
            reg_file[2911] <= 8'h00
            reg_file[2912] <= 8'hA3
            reg_file[2913] <= 8'h03
            reg_file[2914] <= 8'hB7
            reg_file[2915] <= 8'h00
            reg_file[2916] <= 8'h23
            reg_file[2917] <= 8'h03
            reg_file[2918] <= 8'hB7
            reg_file[2919] <= 8'h00
            reg_file[2920] <= 8'hA3
            reg_file[2921] <= 8'h02
            reg_file[2922] <= 8'hB7
            reg_file[2923] <= 8'h00
            reg_file[2924] <= 8'h23
            reg_file[2925] <= 8'h02
            reg_file[2926] <= 8'hB7
            reg_file[2927] <= 8'h00
            reg_file[2928] <= 8'hA3
            reg_file[2929] <= 8'h01
            reg_file[2930] <= 8'hB7
            reg_file[2931] <= 8'h00
            reg_file[2932] <= 8'h23
            reg_file[2933] <= 8'h01
            reg_file[2934] <= 8'hB7
            reg_file[2935] <= 8'h00
            reg_file[2936] <= 8'hA3
            reg_file[2937] <= 8'h00
            reg_file[2938] <= 8'hB7
            reg_file[2939] <= 8'h00
            reg_file[2940] <= 8'h23
            reg_file[2941] <= 8'h00
            reg_file[2942] <= 8'hB7
            reg_file[2943] <= 8'h00
            reg_file[2944] <= 8'h67
            reg_file[2945] <= 8'h80
            reg_file[2946] <= 8'h00
            reg_file[2947] <= 8'h00
            reg_file[2948] <= 8'h93
            reg_file[2949] <= 8'hF5
            reg_file[2950] <= 8'hF5
            reg_file[2951] <= 8'h0F
            reg_file[2952] <= 8'h93
            reg_file[2953] <= 8'h96
            reg_file[2954] <= 8'h85
            reg_file[2955] <= 8'h00
            reg_file[2956] <= 8'hB3
            reg_file[2957] <= 8'hE5
            reg_file[2958] <= 8'hD5
            reg_file[2959] <= 8'h00
            reg_file[2960] <= 8'h93
            reg_file[2961] <= 8'h96
            reg_file[2962] <= 8'h05
            reg_file[2963] <= 8'h01
            reg_file[2964] <= 8'hB3
            reg_file[2965] <= 8'hE5
            reg_file[2966] <= 8'hD5
            reg_file[2967] <= 8'h00
            reg_file[2968] <= 8'h6F
            reg_file[2969] <= 8'hF0
            reg_file[2970] <= 8'hDF
            reg_file[2971] <= 8'hF6
            reg_file[2972] <= 8'h93
            reg_file[2973] <= 8'h96
            reg_file[2974] <= 8'h27
            reg_file[2975] <= 8'h00
            reg_file[2976] <= 8'h97
            reg_file[2977] <= 8'h02
            reg_file[2978] <= 8'h00
            reg_file[2979] <= 8'h00
            reg_file[2980] <= 8'hB3
            reg_file[2981] <= 8'h86
            reg_file[2982] <= 8'h56
            reg_file[2983] <= 8'h00
            reg_file[2984] <= 8'h93
            reg_file[2985] <= 8'h82
            reg_file[2986] <= 8'h00
            reg_file[2987] <= 8'h00
            reg_file[2988] <= 8'hE7
            reg_file[2989] <= 8'h80
            reg_file[2990] <= 8'h06
            reg_file[2991] <= 8'hFA
            reg_file[2992] <= 8'h93
            reg_file[2993] <= 8'h80
            reg_file[2994] <= 8'h02
            reg_file[2995] <= 8'h00
            reg_file[2996] <= 8'h93
            reg_file[2997] <= 8'h87
            reg_file[2998] <= 8'h07
            reg_file[2999] <= 8'hFF
            reg_file[3000] <= 8'h33
            reg_file[3001] <= 8'h07
            reg_file[3002] <= 8'hF7
            reg_file[3003] <= 8'h40
            reg_file[3004] <= 8'h33
            reg_file[3005] <= 8'h06
            reg_file[3006] <= 8'hF6
            reg_file[3007] <= 8'h00
            reg_file[3008] <= 8'hE3
            reg_file[3009] <= 8'h78
            reg_file[3010] <= 8'hC3
            reg_file[3011] <= 8'hF6
            reg_file[3012] <= 8'h6F
            reg_file[3013] <= 8'hF0
            reg_file[3014] <= 8'hDF
            reg_file[3015] <= 8'hF3
            reg_file[3016] <= 8'hB7
            reg_file[3017] <= 8'h17
            reg_file[3018] <= 8'h00
            reg_file[3019] <= 8'h80
            reg_file[3020] <= 8'h03
            reg_file[3021] <= 8'hA7
            reg_file[3022] <= 8'h87
            reg_file[3023] <= 8'h43
            reg_file[3024] <= 8'h83
            reg_file[3025] <= 8'h27
            reg_file[3026] <= 8'h87
            reg_file[3027] <= 8'h14
            reg_file[3028] <= 8'h63
            reg_file[3029] <= 8'h8C
            reg_file[3030] <= 8'h07
            reg_file[3031] <= 8'h04
            reg_file[3032] <= 8'h03
            reg_file[3033] <= 8'hA7
            reg_file[3034] <= 8'h47
            reg_file[3035] <= 8'h00
            reg_file[3036] <= 8'h13
            reg_file[3037] <= 8'h08
            reg_file[3038] <= 8'hF0
            reg_file[3039] <= 8'h01
            reg_file[3040] <= 8'h63
            reg_file[3041] <= 8'h4E
            reg_file[3042] <= 8'hE8
            reg_file[3043] <= 8'h06
            reg_file[3044] <= 8'h13
            reg_file[3045] <= 8'h18
            reg_file[3046] <= 8'h27
            reg_file[3047] <= 8'h00
            reg_file[3048] <= 8'h63
            reg_file[3049] <= 8'h06
            reg_file[3050] <= 8'h05
            reg_file[3051] <= 8'h02
            reg_file[3052] <= 8'h33
            reg_file[3053] <= 8'h83
            reg_file[3054] <= 8'h07
            reg_file[3055] <= 8'h01
            reg_file[3056] <= 8'h23
            reg_file[3057] <= 8'h24
            reg_file[3058] <= 8'hC3
            reg_file[3059] <= 8'h08
            reg_file[3060] <= 8'h83
            reg_file[3061] <= 8'hA8
            reg_file[3062] <= 8'h87
            reg_file[3063] <= 8'h18
            reg_file[3064] <= 8'h13
            reg_file[3065] <= 8'h06
            reg_file[3066] <= 8'h10
            reg_file[3067] <= 8'h00
            reg_file[3068] <= 8'h33
            reg_file[3069] <= 8'h16
            reg_file[3070] <= 8'hE6
            reg_file[3071] <= 8'h00
            reg_file[3072] <= 8'hB3
            reg_file[3073] <= 8'hE8
            reg_file[3074] <= 8'hC8
            reg_file[3075] <= 8'h00
            reg_file[3076] <= 8'h23
            reg_file[3077] <= 8'hA4
            reg_file[3078] <= 8'h17
            reg_file[3079] <= 8'h19
            reg_file[3080] <= 8'h23
            reg_file[3081] <= 8'h24
            reg_file[3082] <= 8'hD3
            reg_file[3083] <= 8'h10
            reg_file[3084] <= 8'h93
            reg_file[3085] <= 8'h06
            reg_file[3086] <= 8'h20
            reg_file[3087] <= 8'h00
            reg_file[3088] <= 8'h63
            reg_file[3089] <= 8'h04
            reg_file[3090] <= 8'hD5
            reg_file[3091] <= 8'h02
            reg_file[3092] <= 8'h13
            reg_file[3093] <= 8'h07
            reg_file[3094] <= 8'h17
            reg_file[3095] <= 8'h00
            reg_file[3096] <= 8'h23
            reg_file[3097] <= 8'hA2
            reg_file[3098] <= 8'hE7
            reg_file[3099] <= 8'h00
            reg_file[3100] <= 8'hB3
            reg_file[3101] <= 8'h87
            reg_file[3102] <= 8'h07
            reg_file[3103] <= 8'h01
            reg_file[3104] <= 8'h23
            reg_file[3105] <= 8'hA4
            reg_file[3106] <= 8'hB7
            reg_file[3107] <= 8'h00
            reg_file[3108] <= 8'h13
            reg_file[3109] <= 8'h05
            reg_file[3110] <= 8'h00
            reg_file[3111] <= 8'h00
            reg_file[3112] <= 8'h67
            reg_file[3113] <= 8'h80
            reg_file[3114] <= 8'h00
            reg_file[3115] <= 8'h00
            reg_file[3116] <= 8'h93
            reg_file[3117] <= 8'h07
            reg_file[3118] <= 8'hC7
            reg_file[3119] <= 8'h14
            reg_file[3120] <= 8'h23
            reg_file[3121] <= 8'h24
            reg_file[3122] <= 8'hF7
            reg_file[3123] <= 8'h14
            reg_file[3124] <= 8'h6F
            reg_file[3125] <= 8'hF0
            reg_file[3126] <= 8'h5F
            reg_file[3127] <= 8'hFA
            reg_file[3128] <= 8'h83
            reg_file[3129] <= 8'hA6
            reg_file[3130] <= 8'hC7
            reg_file[3131] <= 8'h18
            reg_file[3132] <= 8'h13
            reg_file[3133] <= 8'h07
            reg_file[3134] <= 8'h17
            reg_file[3135] <= 8'h00
            reg_file[3136] <= 8'h23
            reg_file[3137] <= 8'hA2
            reg_file[3138] <= 8'hE7
            reg_file[3139] <= 8'h00
            reg_file[3140] <= 8'h33
            reg_file[3141] <= 8'hE6
            reg_file[3142] <= 8'hC6
            reg_file[3143] <= 8'h00
            reg_file[3144] <= 8'h23
            reg_file[3145] <= 8'hA6
            reg_file[3146] <= 8'hC7
            reg_file[3147] <= 8'h18
            reg_file[3148] <= 8'hB3
            reg_file[3149] <= 8'h87
            reg_file[3150] <= 8'h07
            reg_file[3151] <= 8'h01
            reg_file[3152] <= 8'h23
            reg_file[3153] <= 8'hA4
            reg_file[3154] <= 8'hB7
            reg_file[3155] <= 8'h00
            reg_file[3156] <= 8'h13
            reg_file[3157] <= 8'h05
            reg_file[3158] <= 8'h00
            reg_file[3159] <= 8'h00
            reg_file[3160] <= 8'h67
            reg_file[3161] <= 8'h80
            reg_file[3162] <= 8'h00
            reg_file[3163] <= 8'h00
            reg_file[3164] <= 8'h13
            reg_file[3165] <= 8'h05
            reg_file[3166] <= 8'hF0
            reg_file[3167] <= 8'hFF
            reg_file[3168] <= 8'h67
            reg_file[3169] <= 8'h80
            reg_file[3170] <= 8'h00
            reg_file[3171] <= 8'h00
            reg_file[3172] <= 8'h13
            reg_file[3173] <= 8'h01
            reg_file[3174] <= 8'h01
            reg_file[3175] <= 8'hFD
            reg_file[3176] <= 8'hB7
            reg_file[3177] <= 8'h17
            reg_file[3178] <= 8'h00
            reg_file[3179] <= 8'h80
            reg_file[3180] <= 8'h23
            reg_file[3181] <= 8'h2C
            reg_file[3182] <= 8'h41
            reg_file[3183] <= 8'h01
            reg_file[3184] <= 8'h03
            reg_file[3185] <= 8'hAA
            reg_file[3186] <= 8'h87
            reg_file[3187] <= 8'h43
            reg_file[3188] <= 8'h23
            reg_file[3189] <= 8'h20
            reg_file[3190] <= 8'h21
            reg_file[3191] <= 8'h03
            reg_file[3192] <= 8'h23
            reg_file[3193] <= 8'h26
            reg_file[3194] <= 8'h11
            reg_file[3195] <= 8'h02
            reg_file[3196] <= 8'h03
            reg_file[3197] <= 8'h29
            reg_file[3198] <= 8'h8A
            reg_file[3199] <= 8'h14
            reg_file[3200] <= 8'h23
            reg_file[3201] <= 8'h24
            reg_file[3202] <= 8'h81
            reg_file[3203] <= 8'h02
            reg_file[3204] <= 8'h23
            reg_file[3205] <= 8'h22
            reg_file[3206] <= 8'h91
            reg_file[3207] <= 8'h02
            reg_file[3208] <= 8'h23
            reg_file[3209] <= 8'h2E
            reg_file[3210] <= 8'h31
            reg_file[3211] <= 8'h01
            reg_file[3212] <= 8'h23
            reg_file[3213] <= 8'h2A
            reg_file[3214] <= 8'h51
            reg_file[3215] <= 8'h01
            reg_file[3216] <= 8'h23
            reg_file[3217] <= 8'h28
            reg_file[3218] <= 8'h61
            reg_file[3219] <= 8'h01
            reg_file[3220] <= 8'h23
            reg_file[3221] <= 8'h26
            reg_file[3222] <= 8'h71
            reg_file[3223] <= 8'h01
            reg_file[3224] <= 8'h23
            reg_file[3225] <= 8'h24
            reg_file[3226] <= 8'h81
            reg_file[3227] <= 8'h01
            reg_file[3228] <= 8'h63
            reg_file[3229] <= 8'h00
            reg_file[3230] <= 8'h09
            reg_file[3231] <= 8'h04
            reg_file[3232] <= 8'h13
            reg_file[3233] <= 8'h0B
            reg_file[3234] <= 8'h05
            reg_file[3235] <= 8'h00
            reg_file[3236] <= 8'h93
            reg_file[3237] <= 8'h8B
            reg_file[3238] <= 8'h05
            reg_file[3239] <= 8'h00
            reg_file[3240] <= 8'h93
            reg_file[3241] <= 8'h0A
            reg_file[3242] <= 8'h10
            reg_file[3243] <= 8'h00
            reg_file[3244] <= 8'h93
            reg_file[3245] <= 8'h09
            reg_file[3246] <= 8'hF0
            reg_file[3247] <= 8'hFF
            reg_file[3248] <= 8'h83
            reg_file[3249] <= 8'h24
            reg_file[3250] <= 8'h49
            reg_file[3251] <= 8'h00
            reg_file[3252] <= 8'h13
            reg_file[3253] <= 8'h84
            reg_file[3254] <= 8'hF4
            reg_file[3255] <= 8'hFF
            reg_file[3256] <= 8'h63
            reg_file[3257] <= 8'h42
            reg_file[3258] <= 8'h04
            reg_file[3259] <= 8'h02
            reg_file[3260] <= 8'h93
            reg_file[3261] <= 8'h94
            reg_file[3262] <= 8'h24
            reg_file[3263] <= 8'h00
            reg_file[3264] <= 8'hB3
            reg_file[3265] <= 8'h04
            reg_file[3266] <= 8'h99
            reg_file[3267] <= 8'h00
            reg_file[3268] <= 8'h63
            reg_file[3269] <= 8'h84
            reg_file[3270] <= 8'h0B
            reg_file[3271] <= 8'h04
            reg_file[3272] <= 8'h83
            reg_file[3273] <= 8'hA7
            reg_file[3274] <= 8'h44
            reg_file[3275] <= 8'h10
            reg_file[3276] <= 8'h63
            reg_file[3277] <= 8'h80
            reg_file[3278] <= 8'h77
            reg_file[3279] <= 8'h05
            reg_file[3280] <= 8'h13
            reg_file[3281] <= 8'h04
            reg_file[3282] <= 8'hF4
            reg_file[3283] <= 8'hFF
            reg_file[3284] <= 8'h93
            reg_file[3285] <= 8'h84
            reg_file[3286] <= 8'hC4
            reg_file[3287] <= 8'hFF
            reg_file[3288] <= 8'hE3
            reg_file[3289] <= 8'h16
            reg_file[3290] <= 8'h34
            reg_file[3291] <= 8'hFF
            reg_file[3292] <= 8'h83
            reg_file[3293] <= 8'h20
            reg_file[3294] <= 8'hC1
            reg_file[3295] <= 8'h02
            reg_file[3296] <= 8'h03
            reg_file[3297] <= 8'h24
            reg_file[3298] <= 8'h81
            reg_file[3299] <= 8'h02
            reg_file[3300] <= 8'h83
            reg_file[3301] <= 8'h24
            reg_file[3302] <= 8'h41
            reg_file[3303] <= 8'h02
            reg_file[3304] <= 8'h03
            reg_file[3305] <= 8'h29
            reg_file[3306] <= 8'h01
            reg_file[3307] <= 8'h02
            reg_file[3308] <= 8'h83
            reg_file[3309] <= 8'h29
            reg_file[3310] <= 8'hC1
            reg_file[3311] <= 8'h01
            reg_file[3312] <= 8'h03
            reg_file[3313] <= 8'h2A
            reg_file[3314] <= 8'h81
            reg_file[3315] <= 8'h01
            reg_file[3316] <= 8'h83
            reg_file[3317] <= 8'h2A
            reg_file[3318] <= 8'h41
            reg_file[3319] <= 8'h01
            reg_file[3320] <= 8'h03
            reg_file[3321] <= 8'h2B
            reg_file[3322] <= 8'h01
            reg_file[3323] <= 8'h01
            reg_file[3324] <= 8'h83
            reg_file[3325] <= 8'h2B
            reg_file[3326] <= 8'hC1
            reg_file[3327] <= 8'h00
            reg_file[3328] <= 8'h03
            reg_file[3329] <= 8'h2C
            reg_file[3330] <= 8'h81
            reg_file[3331] <= 8'h00
            reg_file[3332] <= 8'h13
            reg_file[3333] <= 8'h01
            reg_file[3334] <= 8'h01
            reg_file[3335] <= 8'h03
            reg_file[3336] <= 8'h67
            reg_file[3337] <= 8'h80
            reg_file[3338] <= 8'h00
            reg_file[3339] <= 8'h00
            reg_file[3340] <= 8'h83
            reg_file[3341] <= 8'h27
            reg_file[3342] <= 8'h49
            reg_file[3343] <= 8'h00
            reg_file[3344] <= 8'h83
            reg_file[3345] <= 8'hA6
            reg_file[3346] <= 8'h44
            reg_file[3347] <= 8'h00
            reg_file[3348] <= 8'h93
            reg_file[3349] <= 8'h87
            reg_file[3350] <= 8'hF7
            reg_file[3351] <= 8'hFF
            reg_file[3352] <= 8'h63
            reg_file[3353] <= 8'h8E
            reg_file[3354] <= 8'h87
            reg_file[3355] <= 8'h04
            reg_file[3356] <= 8'h23
            reg_file[3357] <= 8'hA2
            reg_file[3358] <= 8'h04
            reg_file[3359] <= 8'h00
            reg_file[3360] <= 8'hE3
            reg_file[3361] <= 8'h88
            reg_file[3362] <= 8'h06
            reg_file[3363] <= 8'hFA
            reg_file[3364] <= 8'h83
            reg_file[3365] <= 8'h27
            reg_file[3366] <= 8'h89
            reg_file[3367] <= 8'h18
            reg_file[3368] <= 8'h33
            reg_file[3369] <= 8'h97
            reg_file[3370] <= 8'h8A
            reg_file[3371] <= 8'h00
            reg_file[3372] <= 8'h03
            reg_file[3373] <= 8'h2C
            reg_file[3374] <= 8'h49
            reg_file[3375] <= 8'h00
            reg_file[3376] <= 8'hB3
            reg_file[3377] <= 8'h77
            reg_file[3378] <= 8'hF7
            reg_file[3379] <= 8'h00
            reg_file[3380] <= 8'h63
            reg_file[3381] <= 8'h92
            reg_file[3382] <= 8'h07
            reg_file[3383] <= 8'h02
            reg_file[3384] <= 8'hE7
            reg_file[3385] <= 8'h80
            reg_file[3386] <= 8'h06
            reg_file[3387] <= 8'h00
            reg_file[3388] <= 8'h03
            reg_file[3389] <= 8'h27
            reg_file[3390] <= 8'h49
            reg_file[3391] <= 8'h00
            reg_file[3392] <= 8'h83
            reg_file[3393] <= 8'h27
            reg_file[3394] <= 8'h8A
            reg_file[3395] <= 8'h14
            reg_file[3396] <= 8'h63
            reg_file[3397] <= 8'h14
            reg_file[3398] <= 8'h87
            reg_file[3399] <= 8'h01
            reg_file[3400] <= 8'hE3
            reg_file[3401] <= 8'h04
            reg_file[3402] <= 8'hF9
            reg_file[3403] <= 8'hF8
            reg_file[3404] <= 8'hE3
            reg_file[3405] <= 8'h88
            reg_file[3406] <= 8'h07
            reg_file[3407] <= 8'hF8
            reg_file[3408] <= 8'h13
            reg_file[3409] <= 8'h89
            reg_file[3410] <= 8'h07
            reg_file[3411] <= 8'h00
            reg_file[3412] <= 8'h6F
            reg_file[3413] <= 8'hF0
            reg_file[3414] <= 8'hDF
            reg_file[3415] <= 8'hF5
            reg_file[3416] <= 8'h83
            reg_file[3417] <= 8'h27
            reg_file[3418] <= 8'hC9
            reg_file[3419] <= 8'h18
            reg_file[3420] <= 8'h83
            reg_file[3421] <= 8'hA5
            reg_file[3422] <= 8'h44
            reg_file[3423] <= 8'h08
            reg_file[3424] <= 8'h33
            reg_file[3425] <= 8'h77
            reg_file[3426] <= 8'hF7
            reg_file[3427] <= 8'h00
            reg_file[3428] <= 8'h63
            reg_file[3429] <= 8'h1C
            reg_file[3430] <= 8'h07
            reg_file[3431] <= 8'h00
            reg_file[3432] <= 8'h13
            reg_file[3433] <= 8'h05
            reg_file[3434] <= 8'h0B
            reg_file[3435] <= 8'h00
            reg_file[3436] <= 8'hE7
            reg_file[3437] <= 8'h80
            reg_file[3438] <= 8'h06
            reg_file[3439] <= 8'h00
            reg_file[3440] <= 8'h6F
            reg_file[3441] <= 8'hF0
            reg_file[3442] <= 8'hDF
            reg_file[3443] <= 8'hFC
            reg_file[3444] <= 8'h23
            reg_file[3445] <= 8'h22
            reg_file[3446] <= 8'h89
            reg_file[3447] <= 8'h00
            reg_file[3448] <= 8'h6F
            reg_file[3449] <= 8'hF0
            reg_file[3450] <= 8'h9F
            reg_file[3451] <= 8'hFA
            reg_file[3452] <= 8'h13
            reg_file[3453] <= 8'h85
            reg_file[3454] <= 8'h05
            reg_file[3455] <= 8'h00
            reg_file[3456] <= 8'hE7
            reg_file[3457] <= 8'h80
            reg_file[3458] <= 8'h06
            reg_file[3459] <= 8'h00
            reg_file[3460] <= 8'h6F
            reg_file[3461] <= 8'hF0
            reg_file[3462] <= 8'h9F
            reg_file[3463] <= 8'hFB
            reg_file[3464] <= 8'h10
            reg_file[3465] <= 8'h00
            reg_file[3466] <= 8'h00
            reg_file[3467] <= 8'h00
            reg_file[3468] <= 8'h00
            reg_file[3469] <= 8'h00
            reg_file[3470] <= 8'h00
            reg_file[3471] <= 8'h00
            reg_file[3472] <= 8'h03
            reg_file[3473] <= 8'h7A
            reg_file[3474] <= 8'h52
            reg_file[3475] <= 8'h00
            reg_file[3476] <= 8'h01
            reg_file[3477] <= 8'h7C
            reg_file[3478] <= 8'h01
            reg_file[3479] <= 8'h01
            reg_file[3480] <= 8'h1B
            reg_file[3481] <= 8'h0D
            reg_file[3482] <= 8'h02
            reg_file[3483] <= 8'h00
            reg_file[3484] <= 8'h10
            reg_file[3485] <= 8'h00
            reg_file[3486] <= 8'h00
            reg_file[3487] <= 8'h00
            reg_file[3488] <= 8'h18
            reg_file[3489] <= 8'h00
            reg_file[3490] <= 8'h00
            reg_file[3491] <= 8'h00
            reg_file[3492] <= 8'h84
            reg_file[3493] <= 8'hFB
            reg_file[3494] <= 8'hFF
            reg_file[3495] <= 8'hFF
            reg_file[3496] <= 8'h08
            reg_file[3497] <= 8'h00
            reg_file[3498] <= 8'h00
            reg_file[3499] <= 8'h00
            reg_file[3500] <= 8'h00
            reg_file[3501] <= 8'h00
            reg_file[3502] <= 8'h00
            reg_file[3503] <= 8'h00
            reg_file[3504] <= 8'h10
            reg_file[3505] <= 8'h00
            reg_file[3506] <= 8'h00
            reg_file[3507] <= 8'h00
            reg_file[3508] <= 8'h2C
            reg_file[3509] <= 8'h00
            reg_file[3510] <= 8'h00
            reg_file[3511] <= 8'h00
            reg_file[3512] <= 8'h78
            reg_file[3513] <= 8'hFB
            reg_file[3514] <= 8'hFF
            reg_file[3515] <= 8'hFF
            reg_file[3516] <= 8'h08
            reg_file[3517] <= 8'h00
            reg_file[3518] <= 8'h00
            reg_file[3519] <= 8'h00
            reg_file[3520] <= 8'h00
            reg_file[3521] <= 8'h00
            reg_file[3522] <= 8'h00
            reg_file[3523] <= 8'h00
            reg_file[3524] <= 8'h10
            reg_file[3525] <= 8'h00
            reg_file[3526] <= 8'h00
            reg_file[3527] <= 8'h00
            reg_file[3528] <= 8'h40
            reg_file[3529] <= 8'h00
            reg_file[3530] <= 8'h00
            reg_file[3531] <= 8'h00
            reg_file[3532] <= 8'h6C
            reg_file[3533] <= 8'hFB
            reg_file[3534] <= 8'hFF
            reg_file[3535] <= 8'hFF
            reg_file[3536] <= 8'h08
            reg_file[3537] <= 8'h00
            reg_file[3538] <= 8'h00
            reg_file[3539] <= 8'h00
            reg_file[3540] <= 8'h00
            reg_file[3541] <= 8'h00
            reg_file[3542] <= 8'h00
            reg_file[3543] <= 8'h00
            reg_file[3544] <= 8'h10
            reg_file[3545] <= 8'h00
            reg_file[3546] <= 8'h00
            reg_file[3547] <= 8'h00
            reg_file[3548] <= 8'h54
            reg_file[3549] <= 8'h00
            reg_file[3550] <= 8'h00
            reg_file[3551] <= 8'h00
            reg_file[3552] <= 8'h60
            reg_file[3553] <= 8'hFB
            reg_file[3554] <= 8'hFF
            reg_file[3555] <= 8'hFF
            reg_file[3556] <= 8'h08
            reg_file[3557] <= 8'h00
            reg_file[3558] <= 8'h00
            reg_file[3559] <= 8'h00
            reg_file[3560] <= 8'h00
            reg_file[3561] <= 8'h00
            reg_file[3562] <= 8'h00
            reg_file[3563] <= 8'h00
            reg_file[3564] <= 8'h10
            reg_file[3565] <= 8'h00
            reg_file[3566] <= 8'h00
            reg_file[3567] <= 8'h00
            reg_file[3568] <= 8'h68
            reg_file[3569] <= 8'h00
            reg_file[3570] <= 8'h00
            reg_file[3571] <= 8'h00
            reg_file[3572] <= 8'h54
            reg_file[3573] <= 8'hFB
            reg_file[3574] <= 8'hFF
            reg_file[3575] <= 8'hFF
            reg_file[3576] <= 8'h08
            reg_file[3577] <= 8'h00
            reg_file[3578] <= 8'h00
            reg_file[3579] <= 8'h00
            reg_file[3580] <= 8'h00
            reg_file[3581] <= 8'h00
            reg_file[3582] <= 8'h00
            reg_file[3583] <= 8'h00
            reg_file[3584] <= 8'h10
            reg_file[3585] <= 8'h00
            reg_file[3586] <= 8'h00
            reg_file[3587] <= 8'h00
            reg_file[3588] <= 8'h7C
            reg_file[3589] <= 8'h00
            reg_file[3590] <= 8'h00
            reg_file[3591] <= 8'h00
            reg_file[3592] <= 8'h48
            reg_file[3593] <= 8'hFB
            reg_file[3594] <= 8'hFF
            reg_file[3595] <= 8'hFF
            reg_file[3596] <= 8'h08
            reg_file[3597] <= 8'h00
            reg_file[3598] <= 8'h00
            reg_file[3599] <= 8'h00
            reg_file[3600] <= 8'h00
            reg_file[3601] <= 8'h00
            reg_file[3602] <= 8'h00
            reg_file[3603] <= 8'h00
            reg_file[3604] <= 8'h10
            reg_file[3605] <= 8'h00
            reg_file[3606] <= 8'h00
            reg_file[3607] <= 8'h00
            reg_file[3608] <= 8'h90
            reg_file[3609] <= 8'h00
            reg_file[3610] <= 8'h00
            reg_file[3611] <= 8'h00
            reg_file[3612] <= 8'h3C
            reg_file[3613] <= 8'hFB
            reg_file[3614] <= 8'hFF
            reg_file[3615] <= 8'hFF
            reg_file[3616] <= 8'h08
            reg_file[3617] <= 8'h00
            reg_file[3618] <= 8'h00
            reg_file[3619] <= 8'h00
            reg_file[3620] <= 8'h00
            reg_file[3621] <= 8'h00
            reg_file[3622] <= 8'h00
            reg_file[3623] <= 8'h00
            reg_file[3624] <= 8'h10
            reg_file[3625] <= 8'h00
            reg_file[3626] <= 8'h00
            reg_file[3627] <= 8'h00
            reg_file[3628] <= 8'hA4
            reg_file[3629] <= 8'h00
            reg_file[3630] <= 8'h00
            reg_file[3631] <= 8'h00
            reg_file[3632] <= 8'h30
            reg_file[3633] <= 8'hFB
            reg_file[3634] <= 8'hFF
            reg_file[3635] <= 8'hFF
            reg_file[3636] <= 8'h08
            reg_file[3637] <= 8'h00
            reg_file[3638] <= 8'h00
            reg_file[3639] <= 8'h00
            reg_file[3640] <= 8'h00
            reg_file[3641] <= 8'h00
            reg_file[3642] <= 8'h00
            reg_file[3643] <= 8'h00
            reg_file[3644] <= 8'h10
            reg_file[3645] <= 8'h00
            reg_file[3646] <= 8'h00
            reg_file[3647] <= 8'h00
            reg_file[3648] <= 8'hB8
            reg_file[3649] <= 8'h00
            reg_file[3650] <= 8'h00
            reg_file[3651] <= 8'h00
            reg_file[3652] <= 8'h24
            reg_file[3653] <= 8'hFB
            reg_file[3654] <= 8'hFF
            reg_file[3655] <= 8'hFF
            reg_file[3656] <= 8'h08
            reg_file[3657] <= 8'h00
            reg_file[3658] <= 8'h00
            reg_file[3659] <= 8'h00
            reg_file[3660] <= 8'h00
            reg_file[3661] <= 8'h00
            reg_file[3662] <= 8'h00
            reg_file[3663] <= 8'h00
            reg_file[3664] <= 8'h10
            reg_file[3665] <= 8'h00
            reg_file[3666] <= 8'h00
            reg_file[3667] <= 8'h00
            reg_file[3668] <= 8'hCC
            reg_file[3669] <= 8'h00
            reg_file[3670] <= 8'h00
            reg_file[3671] <= 8'h00
            reg_file[3672] <= 8'h18
            reg_file[3673] <= 8'hFB
            reg_file[3674] <= 8'hFF
            reg_file[3675] <= 8'hFF
            reg_file[3676] <= 8'h08
            reg_file[3677] <= 8'h00
            reg_file[3678] <= 8'h00
            reg_file[3679] <= 8'h00
            reg_file[3680] <= 8'h00
            reg_file[3681] <= 8'h00
            reg_file[3682] <= 8'h00
            reg_file[3683] <= 8'h00
            reg_file[3684] <= 8'h10
            reg_file[3685] <= 8'h00
            reg_file[3686] <= 8'h00
            reg_file[3687] <= 8'h00
            reg_file[3688] <= 8'hE0
            reg_file[3689] <= 8'h00
            reg_file[3690] <= 8'h00
            reg_file[3691] <= 8'h00
            reg_file[3692] <= 8'h0C
            reg_file[3693] <= 8'hFB
            reg_file[3694] <= 8'hFF
            reg_file[3695] <= 8'hFF
            reg_file[3696] <= 8'h08
            reg_file[3697] <= 8'h00
            reg_file[3698] <= 8'h00
            reg_file[3699] <= 8'h00
            reg_file[3700] <= 8'h00
            reg_file[3701] <= 8'h00
            reg_file[3702] <= 8'h00
            reg_file[3703] <= 8'h00
            reg_file[3704] <= 8'h10
            reg_file[3705] <= 8'h00
            reg_file[3706] <= 8'h00
            reg_file[3707] <= 8'h00
            reg_file[3708] <= 8'hF4
            reg_file[3709] <= 8'h00
            reg_file[3710] <= 8'h00
            reg_file[3711] <= 8'h00
            reg_file[3712] <= 8'h00
            reg_file[3713] <= 8'hFB
            reg_file[3714] <= 8'hFF
            reg_file[3715] <= 8'hFF
            reg_file[3716] <= 8'h08
            reg_file[3717] <= 8'h00
            reg_file[3718] <= 8'h00
            reg_file[3719] <= 8'h00
            reg_file[3720] <= 8'h00
            reg_file[3721] <= 8'h00
            reg_file[3722] <= 8'h00
            reg_file[3723] <= 8'h00
            reg_file[3724] <= 8'h00
            reg_file[3725] <= 8'h00
            reg_file[3726] <= 8'h00
            reg_file[3727] <= 8'h00
            reg_file[3728] <= 8'h00
            reg_file[3729] <= 8'h00
            reg_file[3730] <= 8'h00
            reg_file[3731] <= 8'h00
            reg_file[3732] <= 8'h00
            reg_file[3733] <= 8'h00
            reg_file[3734] <= 8'h00
            reg_file[3735] <= 8'h00
            reg_file[3736] <= 8'h00
            reg_file[3737] <= 8'h00
            reg_file[3738] <= 8'h00
            reg_file[3739] <= 8'h00
            reg_file[3740] <= 8'h00
            reg_file[3741] <= 8'h00
            reg_file[3742] <= 8'h00
            reg_file[3743] <= 8'h00
            reg_file[3744] <= 8'h00
            reg_file[3745] <= 8'h00
            reg_file[3746] <= 8'h00
            reg_file[3747] <= 8'h00
            reg_file[3748] <= 8'h00
            reg_file[3749] <= 8'h00
            reg_file[3750] <= 8'h00
            reg_file[3751] <= 8'h00
            reg_file[3752] <= 8'h00
            reg_file[3753] <= 8'h00
            reg_file[3754] <= 8'h00
            reg_file[3755] <= 8'h00
            reg_file[3756] <= 8'h00
            reg_file[3757] <= 8'h00
            reg_file[3758] <= 8'h00
            reg_file[3759] <= 8'h00
            reg_file[3760] <= 8'h00
            reg_file[3761] <= 8'h00
            reg_file[3762] <= 8'h00
            reg_file[3763] <= 8'h00
            reg_file[3764] <= 8'h00
            reg_file[3765] <= 8'h00
            reg_file[3766] <= 8'h00
            reg_file[3767] <= 8'h00
            reg_file[3768] <= 8'h00
            reg_file[3769] <= 8'h00
            reg_file[3770] <= 8'h00
            reg_file[3771] <= 8'h00
            reg_file[3772] <= 8'h00
            reg_file[3773] <= 8'h00
            reg_file[3774] <= 8'h00
            reg_file[3775] <= 8'h00
            reg_file[3776] <= 8'h00
            reg_file[3777] <= 8'h00
            reg_file[3778] <= 8'h00
            reg_file[3779] <= 8'h00
            reg_file[3780] <= 8'h00
            reg_file[3781] <= 8'h00
            reg_file[3782] <= 8'h00
            reg_file[3783] <= 8'h00
            reg_file[3784] <= 8'h00
            reg_file[3785] <= 8'h00
            reg_file[3786] <= 8'h00
            reg_file[3787] <= 8'h00
            reg_file[3788] <= 8'h00
            reg_file[3789] <= 8'h00
            reg_file[3790] <= 8'h00
            reg_file[3791] <= 8'h00
            reg_file[3792] <= 8'h00
            reg_file[3793] <= 8'h00
            reg_file[3794] <= 8'h00
            reg_file[3795] <= 8'h00
            reg_file[3796] <= 8'h00
            reg_file[3797] <= 8'h00
            reg_file[3798] <= 8'h00
            reg_file[3799] <= 8'h00
            reg_file[3800] <= 8'h00
            reg_file[3801] <= 8'h00
            reg_file[3802] <= 8'h00
            reg_file[3803] <= 8'h00
            reg_file[3804] <= 8'h00
            reg_file[3805] <= 8'h00
            reg_file[3806] <= 8'h00
            reg_file[3807] <= 8'h00
            reg_file[3808] <= 8'h00
            reg_file[3809] <= 8'h00
            reg_file[3810] <= 8'h00
            reg_file[3811] <= 8'h00
            reg_file[3812] <= 8'h00
            reg_file[3813] <= 8'h00
            reg_file[3814] <= 8'h00
            reg_file[3815] <= 8'h00
            reg_file[3816] <= 8'h00
            reg_file[3817] <= 8'h00
            reg_file[3818] <= 8'h00
            reg_file[3819] <= 8'h00
            reg_file[3820] <= 8'h00
            reg_file[3821] <= 8'h00
            reg_file[3822] <= 8'h00
            reg_file[3823] <= 8'h00
            reg_file[3824] <= 8'h00
            reg_file[3825] <= 8'h00
            reg_file[3826] <= 8'h00
            reg_file[3827] <= 8'h00
            reg_file[3828] <= 8'h00
            reg_file[3829] <= 8'h00
            reg_file[3830] <= 8'h00
            reg_file[3831] <= 8'h00
            reg_file[3832] <= 8'h00
            reg_file[3833] <= 8'h00
            reg_file[3834] <= 8'h00
            reg_file[3835] <= 8'h00
            reg_file[3836] <= 8'h00
            reg_file[3837] <= 8'h00
            reg_file[3838] <= 8'h00
            reg_file[3839] <= 8'h00
            reg_file[3840] <= 8'h00
            reg_file[3841] <= 8'h00
            reg_file[3842] <= 8'h00
            reg_file[3843] <= 8'h00
            reg_file[3844] <= 8'h00
            reg_file[3845] <= 8'h00
            reg_file[3846] <= 8'h00
            reg_file[3847] <= 8'h00
            reg_file[3848] <= 8'h00
            reg_file[3849] <= 8'h00
            reg_file[3850] <= 8'h00
            reg_file[3851] <= 8'h00
            reg_file[3852] <= 8'h00
            reg_file[3853] <= 8'h00
            reg_file[3854] <= 8'h00
            reg_file[3855] <= 8'h00
            reg_file[3856] <= 8'h00
            reg_file[3857] <= 8'h00
            reg_file[3858] <= 8'h00
            reg_file[3859] <= 8'h00
            reg_file[3860] <= 8'h00
            reg_file[3861] <= 8'h00
            reg_file[3862] <= 8'h00
            reg_file[3863] <= 8'h00
            reg_file[3864] <= 8'h00
            reg_file[3865] <= 8'h00
            reg_file[3866] <= 8'h00
            reg_file[3867] <= 8'h00
            reg_file[3868] <= 8'h00
            reg_file[3869] <= 8'h00
            reg_file[3870] <= 8'h00
            reg_file[3871] <= 8'h00
            reg_file[3872] <= 8'h00
            reg_file[3873] <= 8'h00
            reg_file[3874] <= 8'h00
            reg_file[3875] <= 8'h00
            reg_file[3876] <= 8'h00
            reg_file[3877] <= 8'h00
            reg_file[3878] <= 8'h00
            reg_file[3879] <= 8'h00
            reg_file[3880] <= 8'h00
            reg_file[3881] <= 8'h00
            reg_file[3882] <= 8'h00
            reg_file[3883] <= 8'h00
            reg_file[3884] <= 8'h00
            reg_file[3885] <= 8'h00
            reg_file[3886] <= 8'h00
            reg_file[3887] <= 8'h00
            reg_file[3888] <= 8'h00
            reg_file[3889] <= 8'h00
            reg_file[3890] <= 8'h00
            reg_file[3891] <= 8'h00
            reg_file[3892] <= 8'h00
            reg_file[3893] <= 8'h00
            reg_file[3894] <= 8'h00
            reg_file[3895] <= 8'h00
            reg_file[3896] <= 8'h00
            reg_file[3897] <= 8'h00
            reg_file[3898] <= 8'h00
            reg_file[3899] <= 8'h00
            reg_file[3900] <= 8'h00
            reg_file[3901] <= 8'h00
            reg_file[3902] <= 8'h00
            reg_file[3903] <= 8'h00
            reg_file[3904] <= 8'h00
            reg_file[3905] <= 8'h00
            reg_file[3906] <= 8'h00
            reg_file[3907] <= 8'h00
            reg_file[3908] <= 8'h00
            reg_file[3909] <= 8'h00
            reg_file[3910] <= 8'h00
            reg_file[3911] <= 8'h00
            reg_file[3912] <= 8'h00
            reg_file[3913] <= 8'h00
            reg_file[3914] <= 8'h00
            reg_file[3915] <= 8'h00
            reg_file[3916] <= 8'h00
            reg_file[3917] <= 8'h00
            reg_file[3918] <= 8'h00
            reg_file[3919] <= 8'h00
            reg_file[3920] <= 8'h00
            reg_file[3921] <= 8'h00
            reg_file[3922] <= 8'h00
            reg_file[3923] <= 8'h00
            reg_file[3924] <= 8'h00
            reg_file[3925] <= 8'h00
            reg_file[3926] <= 8'h00
            reg_file[3927] <= 8'h00
            reg_file[3928] <= 8'h00
            reg_file[3929] <= 8'h00
            reg_file[3930] <= 8'h00
            reg_file[3931] <= 8'h00
            reg_file[3932] <= 8'h00
            reg_file[3933] <= 8'h00
            reg_file[3934] <= 8'h00
            reg_file[3935] <= 8'h00
            reg_file[3936] <= 8'h00
            reg_file[3937] <= 8'h00
            reg_file[3938] <= 8'h00
            reg_file[3939] <= 8'h00
            reg_file[3940] <= 8'h00
            reg_file[3941] <= 8'h00
            reg_file[3942] <= 8'h00
            reg_file[3943] <= 8'h00
            reg_file[3944] <= 8'h00
            reg_file[3945] <= 8'h00
            reg_file[3946] <= 8'h00
            reg_file[3947] <= 8'h00
            reg_file[3948] <= 8'h00
            reg_file[3949] <= 8'h00
            reg_file[3950] <= 8'h00
            reg_file[3951] <= 8'h00
            reg_file[3952] <= 8'h00
            reg_file[3953] <= 8'h00
            reg_file[3954] <= 8'h00
            reg_file[3955] <= 8'h00
            reg_file[3956] <= 8'h00
            reg_file[3957] <= 8'h00
            reg_file[3958] <= 8'h00
            reg_file[3959] <= 8'h00
            reg_file[3960] <= 8'h00
            reg_file[3961] <= 8'h00
            reg_file[3962] <= 8'h00
            reg_file[3963] <= 8'h00
            reg_file[3964] <= 8'h00
            reg_file[3965] <= 8'h00
            reg_file[3966] <= 8'h00
            reg_file[3967] <= 8'h00
            reg_file[3968] <= 8'h00
            reg_file[3969] <= 8'h00
            reg_file[3970] <= 8'h00
            reg_file[3971] <= 8'h00
            reg_file[3972] <= 8'h00
            reg_file[3973] <= 8'h00
            reg_file[3974] <= 8'h00
            reg_file[3975] <= 8'h00
            reg_file[3976] <= 8'h00
            reg_file[3977] <= 8'h00
            reg_file[3978] <= 8'h00
            reg_file[3979] <= 8'h00
            reg_file[3980] <= 8'h00
            reg_file[3981] <= 8'h00
            reg_file[3982] <= 8'h00
            reg_file[3983] <= 8'h00
            reg_file[3984] <= 8'h00
            reg_file[3985] <= 8'h00
            reg_file[3986] <= 8'h00
            reg_file[3987] <= 8'h00
            reg_file[3988] <= 8'h00
            reg_file[3989] <= 8'h00
            reg_file[3990] <= 8'h00
            reg_file[3991] <= 8'h00
            reg_file[3992] <= 8'h00
            reg_file[3993] <= 8'h00
            reg_file[3994] <= 8'h00
            reg_file[3995] <= 8'h00
            reg_file[3996] <= 8'h00
            reg_file[3997] <= 8'h00
            reg_file[3998] <= 8'h00
            reg_file[3999] <= 8'h00
            reg_file[4000] <= 8'h00
            reg_file[4001] <= 8'h00
            reg_file[4002] <= 8'h00
            reg_file[4003] <= 8'h00
            reg_file[4004] <= 8'h00
            reg_file[4005] <= 8'h00
            reg_file[4006] <= 8'h00
            reg_file[4007] <= 8'h00
            reg_file[4008] <= 8'h00
            reg_file[4009] <= 8'h00
            reg_file[4010] <= 8'h00
            reg_file[4011] <= 8'h00
            reg_file[4012] <= 8'h00
            reg_file[4013] <= 8'h00
            reg_file[4014] <= 8'h00
            reg_file[4015] <= 8'h00
            reg_file[4016] <= 8'h00
            reg_file[4017] <= 8'h00
            reg_file[4018] <= 8'h00
            reg_file[4019] <= 8'h00
            reg_file[4020] <= 8'h00
            reg_file[4021] <= 8'h00
            reg_file[4022] <= 8'h00
            reg_file[4023] <= 8'h00
            reg_file[4024] <= 8'h00
            reg_file[4025] <= 8'h00
            reg_file[4026] <= 8'h00
            reg_file[4027] <= 8'h00
            reg_file[4028] <= 8'h00
            reg_file[4029] <= 8'h00
            reg_file[4030] <= 8'h00
            reg_file[4031] <= 8'h00
            reg_file[4032] <= 8'h00
            reg_file[4033] <= 8'h00
            reg_file[4034] <= 8'h00
            reg_file[4035] <= 8'h00
            reg_file[4036] <= 8'h00
            reg_file[4037] <= 8'h00
            reg_file[4038] <= 8'h00
            reg_file[4039] <= 8'h00
            reg_file[4040] <= 8'h00
            reg_file[4041] <= 8'h00
            reg_file[4042] <= 8'h00
            reg_file[4043] <= 8'h00
            reg_file[4044] <= 8'h00
            reg_file[4045] <= 8'h00
            reg_file[4046] <= 8'h00
            reg_file[4047] <= 8'h00
            reg_file[4048] <= 8'h00
            reg_file[4049] <= 8'h00
            reg_file[4050] <= 8'h00
            reg_file[4051] <= 8'h00
            reg_file[4052] <= 8'h00
            reg_file[4053] <= 8'h00
            reg_file[4054] <= 8'h00
            reg_file[4055] <= 8'h00
            reg_file[4056] <= 8'h00
            reg_file[4057] <= 8'h00
            reg_file[4058] <= 8'h00
            reg_file[4059] <= 8'h00
            reg_file[4060] <= 8'h00
            reg_file[4061] <= 8'h00
            reg_file[4062] <= 8'h00
            reg_file[4063] <= 8'h00
            reg_file[4064] <= 8'h00
            reg_file[4065] <= 8'h00
            reg_file[4066] <= 8'h00
            reg_file[4067] <= 8'h00
            reg_file[4068] <= 8'h00
            reg_file[4069] <= 8'h00
            reg_file[4070] <= 8'h00
            reg_file[4071] <= 8'h00
            reg_file[4072] <= 8'h00
            reg_file[4073] <= 8'h00
            reg_file[4074] <= 8'h00
            reg_file[4075] <= 8'h00
            reg_file[4076] <= 8'h00
            reg_file[4077] <= 8'h00
            reg_file[4078] <= 8'h00
            reg_file[4079] <= 8'h00
            reg_file[4080] <= 8'h00
            reg_file[4081] <= 8'h00
            reg_file[4082] <= 8'h00
            reg_file[4083] <= 8'h00
            reg_file[4084] <= 8'h00
            reg_file[4085] <= 8'h00
            reg_file[4086] <= 8'h00
            reg_file[4087] <= 8'h00
            reg_file[4088] <= 8'h00
            reg_file[4089] <= 8'h00
            reg_file[4090] <= 8'h00
            reg_file[4091] <= 8'h00
            reg_file[4092] <= 8'h00
            reg_file[4093] <= 8'h00
            reg_file[4094] <= 8'h00
            reg_file[4095] <= 8'h00
            reg_file[4096] <= 8'h7C
            reg_file[4097] <= 8'h00
            reg_file[4098] <= 8'h00
            reg_file[4099] <= 8'h80
            reg_file[4100] <= 8'h00
            reg_file[4101] <= 8'h00
            reg_file[4102] <= 8'h00
            reg_file[4103] <= 8'h00
            reg_file[4104] <= 8'h00
            reg_file[4105] <= 8'h00
            reg_file[4106] <= 8'h00
            reg_file[4107] <= 8'h00
            reg_file[4108] <= 8'h00
            reg_file[4109] <= 8'h00
            reg_file[4110] <= 8'h00
            reg_file[4111] <= 8'h00
            reg_file[4112] <= 8'h00
            reg_file[4113] <= 8'h00
            reg_file[4114] <= 8'h00
            reg_file[4115] <= 8'h00
            reg_file[4116] <= 8'hFC
            reg_file[4117] <= 8'h12
            reg_file[4118] <= 8'h00
            reg_file[4119] <= 8'h80
            reg_file[4120] <= 8'h64
            reg_file[4121] <= 8'h13
            reg_file[4122] <= 8'h00
            reg_file[4123] <= 8'h80
            reg_file[4124] <= 8'hCC
            reg_file[4125] <= 8'h13
            reg_file[4126] <= 8'h00
            reg_file[4127] <= 8'h80
            reg_file[4128] <= 8'h00
            reg_file[4129] <= 8'h00
            reg_file[4130] <= 8'h00
            reg_file[4131] <= 8'h00
            reg_file[4132] <= 8'h00
            reg_file[4133] <= 8'h00
            reg_file[4134] <= 8'h00
            reg_file[4135] <= 8'h00
            reg_file[4136] <= 8'h00
            reg_file[4137] <= 8'h00
            reg_file[4138] <= 8'h00
            reg_file[4139] <= 8'h00
            reg_file[4140] <= 8'h00
            reg_file[4141] <= 8'h00
            reg_file[4142] <= 8'h00
            reg_file[4143] <= 8'h00
            reg_file[4144] <= 8'h00
            reg_file[4145] <= 8'h00
            reg_file[4146] <= 8'h00
            reg_file[4147] <= 8'h00
            reg_file[4148] <= 8'h00
            reg_file[4149] <= 8'h00
            reg_file[4150] <= 8'h00
            reg_file[4151] <= 8'h00
            reg_file[4152] <= 8'h00
            reg_file[4153] <= 8'h00
            reg_file[4154] <= 8'h00
            reg_file[4155] <= 8'h00
            reg_file[4156] <= 8'h00
            reg_file[4157] <= 8'h00
            reg_file[4158] <= 8'h00
            reg_file[4159] <= 8'h00
            reg_file[4160] <= 8'h00
            reg_file[4161] <= 8'h00
            reg_file[4162] <= 8'h00
            reg_file[4163] <= 8'h00
            reg_file[4164] <= 8'h00
            reg_file[4165] <= 8'h00
            reg_file[4166] <= 8'h00
            reg_file[4167] <= 8'h00
            reg_file[4168] <= 8'h00
            reg_file[4169] <= 8'h00
            reg_file[4170] <= 8'h00
            reg_file[4171] <= 8'h00
            reg_file[4172] <= 8'h00
            reg_file[4173] <= 8'h00
            reg_file[4174] <= 8'h00
            reg_file[4175] <= 8'h00
            reg_file[4176] <= 8'h00
            reg_file[4177] <= 8'h00
            reg_file[4178] <= 8'h00
            reg_file[4179] <= 8'h00
            reg_file[4180] <= 8'h00
            reg_file[4181] <= 8'h00
            reg_file[4182] <= 8'h00
            reg_file[4183] <= 8'h00
            reg_file[4184] <= 8'h00
            reg_file[4185] <= 8'h00
            reg_file[4186] <= 8'h00
            reg_file[4187] <= 8'h00
            reg_file[4188] <= 8'h00
            reg_file[4189] <= 8'h00
            reg_file[4190] <= 8'h00
            reg_file[4191] <= 8'h00
            reg_file[4192] <= 8'h00
            reg_file[4193] <= 8'h00
            reg_file[4194] <= 8'h00
            reg_file[4195] <= 8'h00
            reg_file[4196] <= 8'h00
            reg_file[4197] <= 8'h00
            reg_file[4198] <= 8'h00
            reg_file[4199] <= 8'h00
            reg_file[4200] <= 8'h00
            reg_file[4201] <= 8'h00
            reg_file[4202] <= 8'h00
            reg_file[4203] <= 8'h00
            reg_file[4204] <= 8'h00
            reg_file[4205] <= 8'h00
            reg_file[4206] <= 8'h00
            reg_file[4207] <= 8'h00
            reg_file[4208] <= 8'h00
            reg_file[4209] <= 8'h00
            reg_file[4210] <= 8'h00
            reg_file[4211] <= 8'h00
            reg_file[4212] <= 8'h00
            reg_file[4213] <= 8'h00
            reg_file[4214] <= 8'h00
            reg_file[4215] <= 8'h00
            reg_file[4216] <= 8'h00
            reg_file[4217] <= 8'h00
            reg_file[4218] <= 8'h00
            reg_file[4219] <= 8'h00
            reg_file[4220] <= 8'h00
            reg_file[4221] <= 8'h00
            reg_file[4222] <= 8'h00
            reg_file[4223] <= 8'h00
            reg_file[4224] <= 8'h00
            reg_file[4225] <= 8'h00
            reg_file[4226] <= 8'h00
            reg_file[4227] <= 8'h00
            reg_file[4228] <= 8'h00
            reg_file[4229] <= 8'h00
            reg_file[4230] <= 8'h00
            reg_file[4231] <= 8'h00
            reg_file[4232] <= 8'h00
            reg_file[4233] <= 8'h00
            reg_file[4234] <= 8'h00
            reg_file[4235] <= 8'h00
            reg_file[4236] <= 8'h00
            reg_file[4237] <= 8'h00
            reg_file[4238] <= 8'h00
            reg_file[4239] <= 8'h00
            reg_file[4240] <= 8'h00
            reg_file[4241] <= 8'h00
            reg_file[4242] <= 8'h00
            reg_file[4243] <= 8'h00
            reg_file[4244] <= 8'h00
            reg_file[4245] <= 8'h00
            reg_file[4246] <= 8'h00
            reg_file[4247] <= 8'h00
            reg_file[4248] <= 8'h00
            reg_file[4249] <= 8'h00
            reg_file[4250] <= 8'h00
            reg_file[4251] <= 8'h00
            reg_file[4252] <= 8'h00
            reg_file[4253] <= 8'h00
            reg_file[4254] <= 8'h00
            reg_file[4255] <= 8'h00
            reg_file[4256] <= 8'h00
            reg_file[4257] <= 8'h00
            reg_file[4258] <= 8'h00
            reg_file[4259] <= 8'h00
            reg_file[4260] <= 8'h00
            reg_file[4261] <= 8'h00
            reg_file[4262] <= 8'h00
            reg_file[4263] <= 8'h00
            reg_file[4264] <= 8'h00
            reg_file[4265] <= 8'h00
            reg_file[4266] <= 8'h00
            reg_file[4267] <= 8'h00
            reg_file[4268] <= 8'h00
            reg_file[4269] <= 8'h00
            reg_file[4270] <= 8'h00
            reg_file[4271] <= 8'h00
            reg_file[4272] <= 8'h00
            reg_file[4273] <= 8'h00
            reg_file[4274] <= 8'h00
            reg_file[4275] <= 8'h00
            reg_file[4276] <= 8'h00
            reg_file[4277] <= 8'h00
            reg_file[4278] <= 8'h00
            reg_file[4279] <= 8'h00
            reg_file[4280] <= 8'h01
            reg_file[4281] <= 8'h00
            reg_file[4282] <= 8'h00
            reg_file[4283] <= 8'h00
            reg_file[4284] <= 8'h00
            reg_file[4285] <= 8'h00
            reg_file[4286] <= 8'h00
            reg_file[4287] <= 8'h00
            reg_file[4288] <= 8'h0E
            reg_file[4289] <= 8'h33
            reg_file[4290] <= 8'hCD
            reg_file[4291] <= 8'hAB
            reg_file[4292] <= 8'h34
            reg_file[4293] <= 8'h12
            reg_file[4294] <= 8'h6D
            reg_file[4295] <= 8'hE6
            reg_file[4296] <= 8'hEC
            reg_file[4297] <= 8'hDE
            reg_file[4298] <= 8'h05
            reg_file[4299] <= 8'h00
            reg_file[4300] <= 8'h0B
            reg_file[4301] <= 8'h00
            reg_file[4302] <= 8'h00
            reg_file[4303] <= 8'h00
            reg_file[4304] <= 8'h00
            reg_file[4305] <= 8'h00
            reg_file[4306] <= 8'h00
            reg_file[4307] <= 8'h00
            reg_file[4308] <= 8'h00
            reg_file[4309] <= 8'h00
            reg_file[4310] <= 8'h00
            reg_file[4311] <= 8'h00
            reg_file[4312] <= 8'h00
            reg_file[4313] <= 8'h00
            reg_file[4314] <= 8'h00
            reg_file[4315] <= 8'h00
            reg_file[4316] <= 8'h00
            reg_file[4317] <= 8'h00
            reg_file[4318] <= 8'h00
            reg_file[4319] <= 8'h00
            reg_file[4320] <= 8'h00
            reg_file[4321] <= 8'h00
            reg_file[4322] <= 8'h00
            reg_file[4323] <= 8'h00
            reg_file[4324] <= 8'h00
            reg_file[4325] <= 8'h00
            reg_file[4326] <= 8'h00
            reg_file[4327] <= 8'h00
            reg_file[4328] <= 8'h00
            reg_file[4329] <= 8'h00
            reg_file[4330] <= 8'h00
            reg_file[4331] <= 8'h00
            reg_file[4332] <= 8'h00
            reg_file[4333] <= 8'h00
            reg_file[4334] <= 8'h00
            reg_file[4335] <= 8'h00
            reg_file[4336] <= 8'h00
            reg_file[4337] <= 8'h00
            reg_file[4338] <= 8'h00
            reg_file[4339] <= 8'h00
            reg_file[4340] <= 8'h00
            reg_file[4341] <= 8'h00
            reg_file[4342] <= 8'h00
            reg_file[4343] <= 8'h00
            reg_file[4344] <= 8'h00
            reg_file[4345] <= 8'h00
            reg_file[4346] <= 8'h00
            reg_file[4347] <= 8'h00
            reg_file[4348] <= 8'h00
            reg_file[4349] <= 8'h00
            reg_file[4350] <= 8'h00
            reg_file[4351] <= 8'h00
            reg_file[4352] <= 8'h00
            reg_file[4353] <= 8'h00
            reg_file[4354] <= 8'h00
            reg_file[4355] <= 8'h00
            reg_file[4356] <= 8'h00
            reg_file[4357] <= 8'h00
            reg_file[4358] <= 8'h00
            reg_file[4359] <= 8'h00
            reg_file[4360] <= 8'h00
            reg_file[4361] <= 8'h00
            reg_file[4362] <= 8'h00
            reg_file[4363] <= 8'h00
            reg_file[4364] <= 8'h00
            reg_file[4365] <= 8'h00
            reg_file[4366] <= 8'h00
            reg_file[4367] <= 8'h00
            reg_file[4368] <= 8'h00
            reg_file[4369] <= 8'h00
            reg_file[4370] <= 8'h00
            reg_file[4371] <= 8'h00
            reg_file[4372] <= 8'h00
            reg_file[4373] <= 8'h00
            reg_file[4374] <= 8'h00
            reg_file[4375] <= 8'h00
            reg_file[4376] <= 8'h00
            reg_file[4377] <= 8'h00
            reg_file[4378] <= 8'h00
            reg_file[4379] <= 8'h00
            reg_file[4380] <= 8'h00
            reg_file[4381] <= 8'h00
            reg_file[4382] <= 8'h00
            reg_file[4383] <= 8'h00
            reg_file[4384] <= 8'h00
            reg_file[4385] <= 8'h00
            reg_file[4386] <= 8'h00
            reg_file[4387] <= 8'h00
            reg_file[4388] <= 8'h00
            reg_file[4389] <= 8'h00
            reg_file[4390] <= 8'h00
            reg_file[4391] <= 8'h00
            reg_file[4392] <= 8'h00
            reg_file[4393] <= 8'h00
            reg_file[4394] <= 8'h00
            reg_file[4395] <= 8'h00
            reg_file[4396] <= 8'h00
            reg_file[4397] <= 8'h00
            reg_file[4398] <= 8'h00
            reg_file[4399] <= 8'h00
            reg_file[4400] <= 8'h00
            reg_file[4401] <= 8'h00
            reg_file[4402] <= 8'h00
            reg_file[4403] <= 8'h00
            reg_file[4404] <= 8'h00
            reg_file[4405] <= 8'h00
            reg_file[4406] <= 8'h00
            reg_file[4407] <= 8'h00
            reg_file[4408] <= 8'h00
            reg_file[4409] <= 8'h00
            reg_file[4410] <= 8'h00
            reg_file[4411] <= 8'h00
            reg_file[4412] <= 8'h00
            reg_file[4413] <= 8'h00
            reg_file[4414] <= 8'h00
            reg_file[4415] <= 8'h00
            reg_file[4416] <= 8'h00
            reg_file[4417] <= 8'h00
            reg_file[4418] <= 8'h00
            reg_file[4419] <= 8'h00
            reg_file[4420] <= 8'h00
            reg_file[4421] <= 8'h00
            reg_file[4422] <= 8'h00
            reg_file[4423] <= 8'h00
            reg_file[4424] <= 8'h00
            reg_file[4425] <= 8'h00
            reg_file[4426] <= 8'h00
            reg_file[4427] <= 8'h00
            reg_file[4428] <= 8'h00
            reg_file[4429] <= 8'h00
            reg_file[4430] <= 8'h00
            reg_file[4431] <= 8'h00
            reg_file[4432] <= 8'h00
            reg_file[4433] <= 8'h00
            reg_file[4434] <= 8'h00
            reg_file[4435] <= 8'h00
            reg_file[4436] <= 8'h00
            reg_file[4437] <= 8'h00
            reg_file[4438] <= 8'h00
            reg_file[4439] <= 8'h00
            reg_file[4440] <= 8'h00
            reg_file[4441] <= 8'h00
            reg_file[4442] <= 8'h00
            reg_file[4443] <= 8'h00
            reg_file[4444] <= 8'h00
            reg_file[4445] <= 8'h00
            reg_file[4446] <= 8'h00
            reg_file[4447] <= 8'h00
            reg_file[4448] <= 8'h00
            reg_file[4449] <= 8'h00
            reg_file[4450] <= 8'h00
            reg_file[4451] <= 8'h00
            reg_file[4452] <= 8'h00
            reg_file[4453] <= 8'h00
            reg_file[4454] <= 8'h00
            reg_file[4455] <= 8'h00
            reg_file[4456] <= 8'h00
            reg_file[4457] <= 8'h00
            reg_file[4458] <= 8'h00
            reg_file[4459] <= 8'h00
            reg_file[4460] <= 8'h00
            reg_file[4461] <= 8'h00
            reg_file[4462] <= 8'h00
            reg_file[4463] <= 8'h00
            reg_file[4464] <= 8'h00
            reg_file[4465] <= 8'h00
            reg_file[4466] <= 8'h00
            reg_file[4467] <= 8'h00
            reg_file[4468] <= 8'h00
            reg_file[4469] <= 8'h00
            reg_file[4470] <= 8'h00
            reg_file[4471] <= 8'h00
            reg_file[4472] <= 8'h00
            reg_file[4473] <= 8'h00
            reg_file[4474] <= 8'h00
            reg_file[4475] <= 8'h00
            reg_file[4476] <= 8'h00
            reg_file[4477] <= 8'h00
            reg_file[4478] <= 8'h00
            reg_file[4479] <= 8'h00
            reg_file[4480] <= 8'h00
            reg_file[4481] <= 8'h00
            reg_file[4482] <= 8'h00
            reg_file[4483] <= 8'h00
            reg_file[4484] <= 8'h00
            reg_file[4485] <= 8'h00
            reg_file[4486] <= 8'h00
            reg_file[4487] <= 8'h00
            reg_file[4488] <= 8'h00
            reg_file[4489] <= 8'h00
            reg_file[4490] <= 8'h00
            reg_file[4491] <= 8'h00
            reg_file[4492] <= 8'h00
            reg_file[4493] <= 8'h00
            reg_file[4494] <= 8'h00
            reg_file[4495] <= 8'h00
            reg_file[4496] <= 8'h00
            reg_file[4497] <= 8'h00
            reg_file[4498] <= 8'h00
            reg_file[4499] <= 8'h00
            reg_file[4500] <= 8'h00
            reg_file[4501] <= 8'h00
            reg_file[4502] <= 8'h00
            reg_file[4503] <= 8'h00
            reg_file[4504] <= 8'h00
            reg_file[4505] <= 8'h00
            reg_file[4506] <= 8'h00
            reg_file[4507] <= 8'h00
            reg_file[4508] <= 8'h00
            reg_file[4509] <= 8'h00
            reg_file[4510] <= 8'h00
            reg_file[4511] <= 8'h00
            reg_file[4512] <= 8'h00
            reg_file[4513] <= 8'h00
            reg_file[4514] <= 8'h00
            reg_file[4515] <= 8'h00
            reg_file[4516] <= 8'h00
            reg_file[4517] <= 8'h00
            reg_file[4518] <= 8'h00
            reg_file[4519] <= 8'h00
            reg_file[4520] <= 8'h00
            reg_file[4521] <= 8'h00
            reg_file[4522] <= 8'h00
            reg_file[4523] <= 8'h00
            reg_file[4524] <= 8'h00
            reg_file[4525] <= 8'h00
            reg_file[4526] <= 8'h00
            reg_file[4527] <= 8'h00
            reg_file[4528] <= 8'h00
            reg_file[4529] <= 8'h00
            reg_file[4530] <= 8'h00
            reg_file[4531] <= 8'h00
            reg_file[4532] <= 8'h00
            reg_file[4533] <= 8'h00
            reg_file[4534] <= 8'h00
            reg_file[4535] <= 8'h00
            reg_file[4536] <= 8'h00
            reg_file[4537] <= 8'h00
            reg_file[4538] <= 8'h00
            reg_file[4539] <= 8'h00
            reg_file[4540] <= 8'h00
            reg_file[4541] <= 8'h00
            reg_file[4542] <= 8'h00
            reg_file[4543] <= 8'h00
            reg_file[4544] <= 8'h00
            reg_file[4545] <= 8'h00
            reg_file[4546] <= 8'h00
            reg_file[4547] <= 8'h00
            reg_file[4548] <= 8'h00
            reg_file[4549] <= 8'h00
            reg_file[4550] <= 8'h00
            reg_file[4551] <= 8'h00
            reg_file[4552] <= 8'h00
            reg_file[4553] <= 8'h00
            reg_file[4554] <= 8'h00
            reg_file[4555] <= 8'h00
            reg_file[4556] <= 8'h00
            reg_file[4557] <= 8'h00
            reg_file[4558] <= 8'h00
            reg_file[4559] <= 8'h00
            reg_file[4560] <= 8'h00
            reg_file[4561] <= 8'h00
            reg_file[4562] <= 8'h00
            reg_file[4563] <= 8'h00
            reg_file[4564] <= 8'h00
            reg_file[4565] <= 8'h00
            reg_file[4566] <= 8'h00
            reg_file[4567] <= 8'h00
            reg_file[4568] <= 8'h00
            reg_file[4569] <= 8'h00
            reg_file[4570] <= 8'h00
            reg_file[4571] <= 8'h00
            reg_file[4572] <= 8'h00
            reg_file[4573] <= 8'h00
            reg_file[4574] <= 8'h00
            reg_file[4575] <= 8'h00
            reg_file[4576] <= 8'h00
            reg_file[4577] <= 8'h00
            reg_file[4578] <= 8'h00
            reg_file[4579] <= 8'h00
            reg_file[4580] <= 8'h00
            reg_file[4581] <= 8'h00
            reg_file[4582] <= 8'h00
            reg_file[4583] <= 8'h00
            reg_file[4584] <= 8'h00
            reg_file[4585] <= 8'h00
            reg_file[4586] <= 8'h00
            reg_file[4587] <= 8'h00
            reg_file[4588] <= 8'h00
            reg_file[4589] <= 8'h00
            reg_file[4590] <= 8'h00
            reg_file[4591] <= 8'h00
            reg_file[4592] <= 8'h00
            reg_file[4593] <= 8'h00
            reg_file[4594] <= 8'h00
            reg_file[4595] <= 8'h00
            reg_file[4596] <= 8'h00
            reg_file[4597] <= 8'h00
            reg_file[4598] <= 8'h00
            reg_file[4599] <= 8'h00
            reg_file[4600] <= 8'h00
            reg_file[4601] <= 8'h00
            reg_file[4602] <= 8'h00
            reg_file[4603] <= 8'h00
            reg_file[4604] <= 8'h00
            reg_file[4605] <= 8'h00
            reg_file[4606] <= 8'h00
            reg_file[4607] <= 8'h00
            reg_file[4608] <= 8'h00
            reg_file[4609] <= 8'h00
            reg_file[4610] <= 8'h00
            reg_file[4611] <= 8'h00
            reg_file[4612] <= 8'h00
            reg_file[4613] <= 8'h00
            reg_file[4614] <= 8'h00
            reg_file[4615] <= 8'h00
            reg_file[4616] <= 8'h00
            reg_file[4617] <= 8'h00
            reg_file[4618] <= 8'h00
            reg_file[4619] <= 8'h00
            reg_file[4620] <= 8'h00
            reg_file[4621] <= 8'h00
            reg_file[4622] <= 8'h00
            reg_file[4623] <= 8'h00
            reg_file[4624] <= 8'h00
            reg_file[4625] <= 8'h00
            reg_file[4626] <= 8'h00
            reg_file[4627] <= 8'h00
            reg_file[4628] <= 8'h00
            reg_file[4629] <= 8'h00
            reg_file[4630] <= 8'h00
            reg_file[4631] <= 8'h00
            reg_file[4632] <= 8'h00
            reg_file[4633] <= 8'h00
            reg_file[4634] <= 8'h00
            reg_file[4635] <= 8'h00
            reg_file[4636] <= 8'h00
            reg_file[4637] <= 8'h00
            reg_file[4638] <= 8'h00
            reg_file[4639] <= 8'h00
            reg_file[4640] <= 8'h00
            reg_file[4641] <= 8'h00
            reg_file[4642] <= 8'h00
            reg_file[4643] <= 8'h00
            reg_file[4644] <= 8'h00
            reg_file[4645] <= 8'h00
            reg_file[4646] <= 8'h00
            reg_file[4647] <= 8'h00
            reg_file[4648] <= 8'h00
            reg_file[4649] <= 8'h00
            reg_file[4650] <= 8'h00
            reg_file[4651] <= 8'h00
            reg_file[4652] <= 8'h00
            reg_file[4653] <= 8'h00
            reg_file[4654] <= 8'h00
            reg_file[4655] <= 8'h00
            reg_file[4656] <= 8'h00
            reg_file[4657] <= 8'h00
            reg_file[4658] <= 8'h00
            reg_file[4659] <= 8'h00
            reg_file[4660] <= 8'h00
            reg_file[4661] <= 8'h00
            reg_file[4662] <= 8'h00
            reg_file[4663] <= 8'h00
            reg_file[4664] <= 8'h00
            reg_file[4665] <= 8'h00
            reg_file[4666] <= 8'h00
            reg_file[4667] <= 8'h00
            reg_file[4668] <= 8'h00
            reg_file[4669] <= 8'h00
            reg_file[4670] <= 8'h00
            reg_file[4671] <= 8'h00
            reg_file[4672] <= 8'h00
            reg_file[4673] <= 8'h00
            reg_file[4674] <= 8'h00
            reg_file[4675] <= 8'h00
            reg_file[4676] <= 8'h00
            reg_file[4677] <= 8'h00
            reg_file[4678] <= 8'h00
            reg_file[4679] <= 8'h00
            reg_file[4680] <= 8'h00
            reg_file[4681] <= 8'h00
            reg_file[4682] <= 8'h00
            reg_file[4683] <= 8'h00
            reg_file[4684] <= 8'h00
            reg_file[4685] <= 8'h00
            reg_file[4686] <= 8'h00
            reg_file[4687] <= 8'h00
            reg_file[4688] <= 8'h00
            reg_file[4689] <= 8'h00
            reg_file[4690] <= 8'h00
            reg_file[4691] <= 8'h00
            reg_file[4692] <= 8'h00
            reg_file[4693] <= 8'h00
            reg_file[4694] <= 8'h00
            reg_file[4695] <= 8'h00
            reg_file[4696] <= 8'h00
            reg_file[4697] <= 8'h00
            reg_file[4698] <= 8'h00
            reg_file[4699] <= 8'h00
            reg_file[4700] <= 8'h00
            reg_file[4701] <= 8'h00
            reg_file[4702] <= 8'h00
            reg_file[4703] <= 8'h00
            reg_file[4704] <= 8'h00
            reg_file[4705] <= 8'h00
            reg_file[4706] <= 8'h00
            reg_file[4707] <= 8'h00
            reg_file[4708] <= 8'h00
            reg_file[4709] <= 8'h00
            reg_file[4710] <= 8'h00
            reg_file[4711] <= 8'h00
            reg_file[4712] <= 8'h00
            reg_file[4713] <= 8'h00
            reg_file[4714] <= 8'h00
            reg_file[4715] <= 8'h00
            reg_file[4716] <= 8'h00
            reg_file[4717] <= 8'h00
            reg_file[4718] <= 8'h00
            reg_file[4719] <= 8'h00
            reg_file[4720] <= 8'h00
            reg_file[4721] <= 8'h00
            reg_file[4722] <= 8'h00
            reg_file[4723] <= 8'h00
            reg_file[4724] <= 8'h00
            reg_file[4725] <= 8'h00
            reg_file[4726] <= 8'h00
            reg_file[4727] <= 8'h00
            reg_file[4728] <= 8'h00
            reg_file[4729] <= 8'h00
            reg_file[4730] <= 8'h00
            reg_file[4731] <= 8'h00
            reg_file[4732] <= 8'h00
            reg_file[4733] <= 8'h00
            reg_file[4734] <= 8'h00
            reg_file[4735] <= 8'h00
            reg_file[4736] <= 8'h00
            reg_file[4737] <= 8'h00
            reg_file[4738] <= 8'h00
            reg_file[4739] <= 8'h00
            reg_file[4740] <= 8'h00
            reg_file[4741] <= 8'h00
            reg_file[4742] <= 8'h00
            reg_file[4743] <= 8'h00
            reg_file[4744] <= 8'h00
            reg_file[4745] <= 8'h00
            reg_file[4746] <= 8'h00
            reg_file[4747] <= 8'h00
            reg_file[4748] <= 8'h00
            reg_file[4749] <= 8'h00
            reg_file[4750] <= 8'h00
            reg_file[4751] <= 8'h00
            reg_file[4752] <= 8'h00
            reg_file[4753] <= 8'h00
            reg_file[4754] <= 8'h00
            reg_file[4755] <= 8'h00
            reg_file[4756] <= 8'h00
            reg_file[4757] <= 8'h00
            reg_file[4758] <= 8'h00
            reg_file[4759] <= 8'h00
            reg_file[4760] <= 8'h00
            reg_file[4761] <= 8'h00
            reg_file[4762] <= 8'h00
            reg_file[4763] <= 8'h00
            reg_file[4764] <= 8'h00
            reg_file[4765] <= 8'h00
            reg_file[4766] <= 8'h00
            reg_file[4767] <= 8'h00
            reg_file[4768] <= 8'h00
            reg_file[4769] <= 8'h00
            reg_file[4770] <= 8'h00
            reg_file[4771] <= 8'h00
            reg_file[4772] <= 8'h00
            reg_file[4773] <= 8'h00
            reg_file[4774] <= 8'h00
            reg_file[4775] <= 8'h00
            reg_file[4776] <= 8'h00
            reg_file[4777] <= 8'h00
            reg_file[4778] <= 8'h00
            reg_file[4779] <= 8'h00
            reg_file[4780] <= 8'h00
            reg_file[4781] <= 8'h00
            reg_file[4782] <= 8'h00
            reg_file[4783] <= 8'h00
            reg_file[4784] <= 8'h00
            reg_file[4785] <= 8'h00
            reg_file[4786] <= 8'h00
            reg_file[4787] <= 8'h00
            reg_file[4788] <= 8'h00
            reg_file[4789] <= 8'h00
            reg_file[4790] <= 8'h00
            reg_file[4791] <= 8'h00
            reg_file[4792] <= 8'h00
            reg_file[4793] <= 8'h00
            reg_file[4794] <= 8'h00
            reg_file[4795] <= 8'h00
            reg_file[4796] <= 8'h00
            reg_file[4797] <= 8'h00
            reg_file[4798] <= 8'h00
            reg_file[4799] <= 8'h00
            reg_file[4800] <= 8'h00
            reg_file[4801] <= 8'h00
            reg_file[4802] <= 8'h00
            reg_file[4803] <= 8'h00
            reg_file[4804] <= 8'h00
            reg_file[4805] <= 8'h00
            reg_file[4806] <= 8'h00
            reg_file[4807] <= 8'h00
            reg_file[4808] <= 8'h00
            reg_file[4809] <= 8'h00
            reg_file[4810] <= 8'h00
            reg_file[4811] <= 8'h00
            reg_file[4812] <= 8'h00
            reg_file[4813] <= 8'h00
            reg_file[4814] <= 8'h00
            reg_file[4815] <= 8'h00
            reg_file[4816] <= 8'h00
            reg_file[4817] <= 8'h00
            reg_file[4818] <= 8'h00
            reg_file[4819] <= 8'h00
            reg_file[4820] <= 8'h00
            reg_file[4821] <= 8'h00
            reg_file[4822] <= 8'h00
            reg_file[4823] <= 8'h00
            reg_file[4824] <= 8'h00
            reg_file[4825] <= 8'h00
            reg_file[4826] <= 8'h00
            reg_file[4827] <= 8'h00
            reg_file[4828] <= 8'h00
            reg_file[4829] <= 8'h00
            reg_file[4830] <= 8'h00
            reg_file[4831] <= 8'h00
            reg_file[4832] <= 8'h00
            reg_file[4833] <= 8'h00
            reg_file[4834] <= 8'h00
            reg_file[4835] <= 8'h00
            reg_file[4836] <= 8'h00
            reg_file[4837] <= 8'h00
            reg_file[4838] <= 8'h00
            reg_file[4839] <= 8'h00
            reg_file[4840] <= 8'h00
            reg_file[4841] <= 8'h00
            reg_file[4842] <= 8'h00
            reg_file[4843] <= 8'h00
            reg_file[4844] <= 8'h00
            reg_file[4845] <= 8'h00
            reg_file[4846] <= 8'h00
            reg_file[4847] <= 8'h00
            reg_file[4848] <= 8'h00
            reg_file[4849] <= 8'h00
            reg_file[4850] <= 8'h00
            reg_file[4851] <= 8'h00
            reg_file[4852] <= 8'h00
            reg_file[4853] <= 8'h00
            reg_file[4854] <= 8'h00
            reg_file[4855] <= 8'h00
            reg_file[4856] <= 8'h00
            reg_file[4857] <= 8'h00
            reg_file[4858] <= 8'h00
            reg_file[4859] <= 8'h00
            reg_file[4860] <= 8'h00
            reg_file[4861] <= 8'h00
            reg_file[4862] <= 8'h00
            reg_file[4863] <= 8'h00
            reg_file[4864] <= 8'h00
            reg_file[4865] <= 8'h00
            reg_file[4866] <= 8'h00
            reg_file[4867] <= 8'h00
            reg_file[4868] <= 8'h00
            reg_file[4869] <= 8'h00
            reg_file[4870] <= 8'h00
            reg_file[4871] <= 8'h00
            reg_file[4872] <= 8'h00
            reg_file[4873] <= 8'h00
            reg_file[4874] <= 8'h00
            reg_file[4875] <= 8'h00
            reg_file[4876] <= 8'h00
            reg_file[4877] <= 8'h00
            reg_file[4878] <= 8'h00
            reg_file[4879] <= 8'h00
            reg_file[4880] <= 8'h00
            reg_file[4881] <= 8'h00
            reg_file[4882] <= 8'h00
            reg_file[4883] <= 8'h00
            reg_file[4884] <= 8'h00
            reg_file[4885] <= 8'h00
            reg_file[4886] <= 8'h00
            reg_file[4887] <= 8'h00
            reg_file[4888] <= 8'h00
            reg_file[4889] <= 8'h00
            reg_file[4890] <= 8'h00
            reg_file[4891] <= 8'h00
            reg_file[4892] <= 8'h00
            reg_file[4893] <= 8'h00
            reg_file[4894] <= 8'h00
            reg_file[4895] <= 8'h00
            reg_file[4896] <= 8'h00
            reg_file[4897] <= 8'h00
            reg_file[4898] <= 8'h00
            reg_file[4899] <= 8'h00
            reg_file[4900] <= 8'h00
            reg_file[4901] <= 8'h00
            reg_file[4902] <= 8'h00
            reg_file[4903] <= 8'h00
            reg_file[4904] <= 8'h00
            reg_file[4905] <= 8'h00
            reg_file[4906] <= 8'h00
            reg_file[4907] <= 8'h00
            reg_file[4908] <= 8'h00
            reg_file[4909] <= 8'h00
            reg_file[4910] <= 8'h00
            reg_file[4911] <= 8'h00
            reg_file[4912] <= 8'h00
            reg_file[4913] <= 8'h00
            reg_file[4914] <= 8'h00
            reg_file[4915] <= 8'h00
            reg_file[4916] <= 8'h00
            reg_file[4917] <= 8'h00
            reg_file[4918] <= 8'h00
            reg_file[4919] <= 8'h00
            reg_file[4920] <= 8'h00
            reg_file[4921] <= 8'h00
            reg_file[4922] <= 8'h00
            reg_file[4923] <= 8'h00
            reg_file[4924] <= 8'h00
            reg_file[4925] <= 8'h00
            reg_file[4926] <= 8'h00
            reg_file[4927] <= 8'h00
            reg_file[4928] <= 8'h00
            reg_file[4929] <= 8'h00
            reg_file[4930] <= 8'h00
            reg_file[4931] <= 8'h00
            reg_file[4932] <= 8'h00
            reg_file[4933] <= 8'h00
            reg_file[4934] <= 8'h00
            reg_file[4935] <= 8'h00
            reg_file[4936] <= 8'h00
            reg_file[4937] <= 8'h00
            reg_file[4938] <= 8'h00
            reg_file[4939] <= 8'h00
            reg_file[4940] <= 8'h00
            reg_file[4941] <= 8'h00
            reg_file[4942] <= 8'h00
            reg_file[4943] <= 8'h00
            reg_file[4944] <= 8'h00
            reg_file[4945] <= 8'h00
            reg_file[4946] <= 8'h00
            reg_file[4947] <= 8'h00
            reg_file[4948] <= 8'h00
            reg_file[4949] <= 8'h00
            reg_file[4950] <= 8'h00
            reg_file[4951] <= 8'h00
            reg_file[4952] <= 8'h00
            reg_file[4953] <= 8'h00
            reg_file[4954] <= 8'h00
            reg_file[4955] <= 8'h00
            reg_file[4956] <= 8'h00
            reg_file[4957] <= 8'h00
            reg_file[4958] <= 8'h00
            reg_file[4959] <= 8'h00
            reg_file[4960] <= 8'h00
            reg_file[4961] <= 8'h00
            reg_file[4962] <= 8'h00
            reg_file[4963] <= 8'h00
            reg_file[4964] <= 8'h00
            reg_file[4965] <= 8'h00
            reg_file[4966] <= 8'h00
            reg_file[4967] <= 8'h00
            reg_file[4968] <= 8'h00
            reg_file[4969] <= 8'h00
            reg_file[4970] <= 8'h00
            reg_file[4971] <= 8'h00
            reg_file[4972] <= 8'h00
            reg_file[4973] <= 8'h00
            reg_file[4974] <= 8'h00
            reg_file[4975] <= 8'h00
            reg_file[4976] <= 8'h00
            reg_file[4977] <= 8'h00
            reg_file[4978] <= 8'h00
            reg_file[4979] <= 8'h00
            reg_file[4980] <= 8'h00
            reg_file[4981] <= 8'h00
            reg_file[4982] <= 8'h00
            reg_file[4983] <= 8'h00
            reg_file[4984] <= 8'h00
            reg_file[4985] <= 8'h00
            reg_file[4986] <= 8'h00
            reg_file[4987] <= 8'h00
            reg_file[4988] <= 8'h00
            reg_file[4989] <= 8'h00
            reg_file[4990] <= 8'h00
            reg_file[4991] <= 8'h00
            reg_file[4992] <= 8'h00
            reg_file[4993] <= 8'h00
            reg_file[4994] <= 8'h00
            reg_file[4995] <= 8'h00
            reg_file[4996] <= 8'h00
            reg_file[4997] <= 8'h00
            reg_file[4998] <= 8'h00
            reg_file[4999] <= 8'h00
            reg_file[5000] <= 8'h00
            reg_file[5001] <= 8'h00
            reg_file[5002] <= 8'h00
            reg_file[5003] <= 8'h00
            reg_file[5004] <= 8'h00
            reg_file[5005] <= 8'h00
            reg_file[5006] <= 8'h00
            reg_file[5007] <= 8'h00
            reg_file[5008] <= 8'h00
            reg_file[5009] <= 8'h00
            reg_file[5010] <= 8'h00
            reg_file[5011] <= 8'h00
            reg_file[5012] <= 8'h00
            reg_file[5013] <= 8'h00
            reg_file[5014] <= 8'h00
            reg_file[5015] <= 8'h00
            reg_file[5016] <= 8'h00
            reg_file[5017] <= 8'h00
            reg_file[5018] <= 8'h00
            reg_file[5019] <= 8'h00
            reg_file[5020] <= 8'h00
            reg_file[5021] <= 8'h00
            reg_file[5022] <= 8'h00
            reg_file[5023] <= 8'h00
            reg_file[5024] <= 8'h00
            reg_file[5025] <= 8'h00
            reg_file[5026] <= 8'h00
            reg_file[5027] <= 8'h00
            reg_file[5028] <= 8'h00
            reg_file[5029] <= 8'h00
            reg_file[5030] <= 8'h00
            reg_file[5031] <= 8'h00
            reg_file[5032] <= 8'h00
            reg_file[5033] <= 8'h00
            reg_file[5034] <= 8'h00
            reg_file[5035] <= 8'h00
            reg_file[5036] <= 8'h00
            reg_file[5037] <= 8'h00
            reg_file[5038] <= 8'h00
            reg_file[5039] <= 8'h00
            reg_file[5040] <= 8'h00
            reg_file[5041] <= 8'h00
            reg_file[5042] <= 8'h00
            reg_file[5043] <= 8'h00
            reg_file[5044] <= 8'h00
            reg_file[5045] <= 8'h00
            reg_file[5046] <= 8'h00
            reg_file[5047] <= 8'h00
            reg_file[5048] <= 8'h00
            reg_file[5049] <= 8'h00
            reg_file[5050] <= 8'h00
            reg_file[5051] <= 8'h00
            reg_file[5052] <= 8'h00
            reg_file[5053] <= 8'h00
            reg_file[5054] <= 8'h00
            reg_file[5055] <= 8'h00
            reg_file[5056] <= 8'h00
            reg_file[5057] <= 8'h00
            reg_file[5058] <= 8'h00
            reg_file[5059] <= 8'h00
            reg_file[5060] <= 8'h00
            reg_file[5061] <= 8'h00
            reg_file[5062] <= 8'h00
            reg_file[5063] <= 8'h00
            reg_file[5064] <= 8'h00
            reg_file[5065] <= 8'h00
            reg_file[5066] <= 8'h00
            reg_file[5067] <= 8'h00
            reg_file[5068] <= 8'h00
            reg_file[5069] <= 8'h00
            reg_file[5070] <= 8'h00
            reg_file[5071] <= 8'h00
            reg_file[5072] <= 8'h00
            reg_file[5073] <= 8'h00
            reg_file[5074] <= 8'h00
            reg_file[5075] <= 8'h00
            reg_file[5076] <= 8'h00
            reg_file[5077] <= 8'h00
            reg_file[5078] <= 8'h00
            reg_file[5079] <= 8'h00
            reg_file[5080] <= 8'h00
            reg_file[5081] <= 8'h00
            reg_file[5082] <= 8'h00
            reg_file[5083] <= 8'h00
            reg_file[5084] <= 8'h00
            reg_file[5085] <= 8'h00
            reg_file[5086] <= 8'h00
            reg_file[5087] <= 8'h00
            reg_file[5088] <= 8'h00
            reg_file[5089] <= 8'h00
            reg_file[5090] <= 8'h00
            reg_file[5091] <= 8'h00
            reg_file[5092] <= 8'h00
            reg_file[5093] <= 8'h00
            reg_file[5094] <= 8'h00
            reg_file[5095] <= 8'h00
            reg_file[5096] <= 8'h00
            reg_file[5097] <= 8'h00
            reg_file[5098] <= 8'h00
            reg_file[5099] <= 8'h00
            reg_file[5100] <= 8'h00
            reg_file[5101] <= 8'h00
            reg_file[5102] <= 8'h00
            reg_file[5103] <= 8'h00
            reg_file[5104] <= 8'h00
            reg_file[5105] <= 8'h00
            reg_file[5106] <= 8'h00
            reg_file[5107] <= 8'h00
            reg_file[5108] <= 8'h00
            reg_file[5109] <= 8'h00
            reg_file[5110] <= 8'h00
            reg_file[5111] <= 8'h00
            reg_file[5112] <= 8'h00
            reg_file[5113] <= 8'h00
            reg_file[5114] <= 8'h00
            reg_file[5115] <= 8'h00
            reg_file[5116] <= 8'h00
            reg_file[5117] <= 8'h00
            reg_file[5118] <= 8'h00
            reg_file[5119] <= 8'h00
            reg_file[5120] <= 8'h00
            reg_file[5121] <= 8'h00
            reg_file[5122] <= 8'h00
            reg_file[5123] <= 8'h00
            reg_file[5124] <= 8'h00
            reg_file[5125] <= 8'h00
            reg_file[5126] <= 8'h00
            reg_file[5127] <= 8'h00
            reg_file[5128] <= 8'h00
            reg_file[5129] <= 8'h00
            reg_file[5130] <= 8'h00
            reg_file[5131] <= 8'h00
            reg_file[5132] <= 8'h00
            reg_file[5133] <= 8'h00
            reg_file[5134] <= 8'h00
            reg_file[5135] <= 8'h00
            reg_file[5136] <= 8'h00
            reg_file[5137] <= 8'h00
            reg_file[5138] <= 8'h00
            reg_file[5139] <= 8'h00
            reg_file[5140] <= 8'h00
            reg_file[5141] <= 8'h00
            reg_file[5142] <= 8'h00
            reg_file[5143] <= 8'h00
            reg_file[5144] <= 8'h00
            reg_file[5145] <= 8'h00
            reg_file[5146] <= 8'h00
            reg_file[5147] <= 8'h00
            reg_file[5148] <= 8'h00
            reg_file[5149] <= 8'h00
            reg_file[5150] <= 8'h00
            reg_file[5151] <= 8'h00
            reg_file[5152] <= 8'h00
            reg_file[5153] <= 8'h00
            reg_file[5154] <= 8'h00
            reg_file[5155] <= 8'h00
            reg_file[5156] <= 8'h00
            reg_file[5157] <= 8'h00
            reg_file[5158] <= 8'h00
            reg_file[5159] <= 8'h00
            reg_file[5160] <= 8'h00
            reg_file[5161] <= 8'h00
            reg_file[5162] <= 8'h00
            reg_file[5163] <= 8'h00
            reg_file[5164] <= 8'h00
            reg_file[5165] <= 8'h00
            reg_file[5166] <= 8'h00
            reg_file[5167] <= 8'h00
            reg_file[5168] <= 8'h00
            reg_file[5169] <= 8'h00
            reg_file[5170] <= 8'h00
            reg_file[5171] <= 8'h00
            reg_file[5172] <= 8'h00
            reg_file[5173] <= 8'h00
            reg_file[5174] <= 8'h00
            reg_file[5175] <= 8'h00
            reg_file[5176] <= 8'h10
            reg_file[5177] <= 8'h10
            reg_file[5178] <= 8'h00
            reg_file[5179] <= 8'h80
            reg_file[5180] <= 8'h10
            reg_file[5181] <= 8'h10
            reg_file[5182] <= 8'h00
            reg_file[5183] <= 8'h80
            reg_file[5184] <= 8'h00
            reg_file[5185] <= 8'h00
            reg_file[5186] <= 8'h00
            reg_file[5187] <= 8'h00
            reg_file[5188] <= 8'h00
            reg_file[5189] <= 8'h00
            reg_file[5190] <= 8'h00
            reg_file[5191] <= 8'h00
            reg_file[5192] <= 8'h00
            reg_file[5193] <= 8'h00
            reg_file[5194] <= 8'h00
            reg_file[5195] <= 8'h00
            reg_file[5196] <= 8'h00
            reg_file[5197] <= 8'h00
            reg_file[5198] <= 8'h00
            reg_file[5199] <= 8'h00
            reg_file[5200] <= 8'h00
            reg_file[5201] <= 8'h00
            reg_file[5202] <= 8'h00
            reg_file[5203] <= 8'h00
            reg_file[5204] <= 8'h00
            reg_file[5205] <= 8'h00
            reg_file[5206] <= 8'h00
            reg_file[5207] <= 8'h00
            reg_file[5208] <= 8'h00
            reg_file[5209] <= 8'h00
            reg_file[5210] <= 8'h00
            reg_file[5211] <= 8'h00
            reg_file[5212] <= 8'h00
            reg_file[5213] <= 8'h00
            reg_file[5214] <= 8'h00
            reg_file[5215] <= 8'h00
            reg_file[5216] <= 8'h00
            reg_file[5217] <= 8'h00
            reg_file[5218] <= 8'h00
            reg_file[5219] <= 8'h00
            reg_file[5220] <= 8'h00
            reg_file[5221] <= 8'h00
            reg_file[5222] <= 8'h00
            reg_file[5223] <= 8'h00
            reg_file[5224] <= 8'h00
            reg_file[5225] <= 8'h00
            reg_file[5226] <= 8'h00
            reg_file[5227] <= 8'h00
            reg_file[5228] <= 8'h00
            reg_file[5229] <= 8'h00
            reg_file[5230] <= 8'h00
            reg_file[5231] <= 8'h00
            reg_file[5232] <= 8'h00
            reg_file[5233] <= 8'h00
            reg_file[5234] <= 8'h00
            reg_file[5235] <= 8'h00
            reg_file[5236] <= 8'h00
            reg_file[5237] <= 8'h00
            reg_file[5238] <= 8'h00
            reg_file[5239] <= 8'h00
            reg_file[5240] <= 8'h00
            reg_file[5241] <= 8'h00
            reg_file[5242] <= 8'h00
            reg_file[5243] <= 8'h00
            reg_file[5244] <= 8'h00
            reg_file[5245] <= 8'h00
            reg_file[5246] <= 8'h00
            reg_file[5247] <= 8'h00
            reg_file[5248] <= 8'h00
            reg_file[5249] <= 8'h00
            reg_file[5250] <= 8'h00
            reg_file[5251] <= 8'h00
            reg_file[5252] <= 8'h00
            reg_file[5253] <= 8'h00
            reg_file[5254] <= 8'h00
            reg_file[5255] <= 8'h00
            reg_file[5256] <= 8'h00
            reg_file[5257] <= 8'h00
            reg_file[5258] <= 8'h00
            reg_file[5259] <= 8'h00
            reg_file[5260] <= 8'h00
            reg_file[5261] <= 8'h00
            reg_file[5262] <= 8'h00
            reg_file[5263] <= 8'h00
            reg_file[5264] <= 8'h00
            reg_file[5265] <= 8'h00
            reg_file[5266] <= 8'h00
            reg_file[5267] <= 8'h00
            reg_file[5268] <= 8'h00
            reg_file[5269] <= 8'h00
            reg_file[5270] <= 8'h00
            reg_file[5271] <= 8'h00
            reg_file[5272] <= 8'h00
            reg_file[5273] <= 8'h00
            reg_file[5274] <= 8'h00
            reg_file[5275] <= 8'h00
            reg_file[5276] <= 8'h00
            reg_file[5277] <= 8'h00
            reg_file[5278] <= 8'h00
            reg_file[5279] <= 8'h00
            reg_file[5280] <= 8'h00
            reg_file[5281] <= 8'h00
            reg_file[5282] <= 8'h00
            reg_file[5283] <= 8'h00
            reg_file[5284] <= 8'h00
            reg_file[5285] <= 8'h00
            reg_file[5286] <= 8'h00
            reg_file[5287] <= 8'h00
            reg_file[5288] <= 8'h00
            reg_file[5289] <= 8'h00
            reg_file[5290] <= 8'h00
            reg_file[5291] <= 8'h00
            reg_file[5292] <= 8'h00
            reg_file[5293] <= 8'h00
            reg_file[5294] <= 8'h00
            reg_file[5295] <= 8'h00
            reg_file[5296] <= 8'h00
            reg_file[5297] <= 8'h00
            reg_file[5298] <= 8'h00
            reg_file[5299] <= 8'h00
            reg_file[5300] <= 8'h00
            reg_file[5301] <= 8'h00
            reg_file[5302] <= 8'h00
            reg_file[5303] <= 8'h00
            reg_file[5304] <= 8'h00
            reg_file[5305] <= 8'h00
            reg_file[5306] <= 8'h00
            reg_file[5307] <= 8'h00
            reg_file[5308] <= 8'h00
            reg_file[5309] <= 8'h00
            reg_file[5310] <= 8'h00
            reg_file[5311] <= 8'h00
            reg_file[5312] <= 8'h00
            reg_file[5313] <= 8'h00
            reg_file[5314] <= 8'h00
            reg_file[5315] <= 8'h00
            reg_file[5316] <= 8'h00
            reg_file[5317] <= 8'h00
            reg_file[5318] <= 8'h00
            reg_file[5319] <= 8'h00
            reg_file[5320] <= 8'h00
            reg_file[5321] <= 8'h00
            reg_file[5322] <= 8'h00
            reg_file[5323] <= 8'h00
            reg_file[5324] <= 8'h00
            reg_file[5325] <= 8'h00
            reg_file[5326] <= 8'h00
            reg_file[5327] <= 8'h00
            reg_file[5328] <= 8'h00
            reg_file[5329] <= 8'h00
            reg_file[5330] <= 8'h00
            reg_file[5331] <= 8'h00
            reg_file[5332] <= 8'h00
            reg_file[5333] <= 8'h00
            reg_file[5334] <= 8'h00
            reg_file[5335] <= 8'h00
            reg_file[5336] <= 8'h00
            reg_file[5337] <= 8'h00
            reg_file[5338] <= 8'h00
            reg_file[5339] <= 8'h00
            reg_file[5340] <= 8'h00
            reg_file[5341] <= 8'h00
            reg_file[5342] <= 8'h00
            reg_file[5343] <= 8'h00
            reg_file[5344] <= 8'h00
            reg_file[5345] <= 8'h00
            reg_file[5346] <= 8'h00
            reg_file[5347] <= 8'h00
            reg_file[5348] <= 8'h00
            reg_file[5349] <= 8'h00
            reg_file[5350] <= 8'h00
            reg_file[5351] <= 8'h00
            reg_file[5352] <= 8'h00
            reg_file[5353] <= 8'h00
            reg_file[5354] <= 8'h00
            reg_file[5355] <= 8'h00
            reg_file[5356] <= 8'h00
            reg_file[5357] <= 8'h00
            reg_file[5358] <= 8'h00
            reg_file[5359] <= 8'h00
            reg_file[5360] <= 8'h00
            reg_file[5361] <= 8'h00
            reg_file[5362] <= 8'h00
            reg_file[5363] <= 8'h00
            reg_file[5364] <= 8'h00
            reg_file[5365] <= 8'h00
            reg_file[5366] <= 8'h00
            reg_file[5367] <= 8'h00
            reg_file[5368] <= 8'h00
            reg_file[5369] <= 8'h00
            reg_file[5370] <= 8'h00
            reg_file[5371] <= 8'h00
            reg_file[5372] <= 8'h00
            reg_file[5373] <= 8'h00
            reg_file[5374] <= 8'h00
            reg_file[5375] <= 8'h00
            reg_file[5376] <= 8'h00
            reg_file[5377] <= 8'h00
            reg_file[5378] <= 8'h00
            reg_file[5379] <= 8'h00
            reg_file[5380] <= 8'h00
            reg_file[5381] <= 8'h00
            reg_file[5382] <= 8'h00
            reg_file[5383] <= 8'h00
            reg_file[5384] <= 8'h00
            reg_file[5385] <= 8'h00
            reg_file[5386] <= 8'h00
            reg_file[5387] <= 8'h00
            reg_file[5388] <= 8'h00
            reg_file[5389] <= 8'h00
            reg_file[5390] <= 8'h00
            reg_file[5391] <= 8'h00
            reg_file[5392] <= 8'h00
            reg_file[5393] <= 8'h00
            reg_file[5394] <= 8'h00
            reg_file[5395] <= 8'h00
            reg_file[5396] <= 8'h00
            reg_file[5397] <= 8'h00
            reg_file[5398] <= 8'h00
            reg_file[5399] <= 8'h00
            reg_file[5400] <= 8'h00
            reg_file[5401] <= 8'h00
            reg_file[5402] <= 8'h00
            reg_file[5403] <= 8'h00
            reg_file[5404] <= 8'h00
            reg_file[5405] <= 8'h00
            reg_file[5406] <= 8'h00
            reg_file[5407] <= 8'h00
            reg_file[5408] <= 8'h00
            reg_file[5409] <= 8'h00
            reg_file[5410] <= 8'h00
            reg_file[5411] <= 8'h00
            reg_file[5412] <= 8'h00
            reg_file[5413] <= 8'h00
            reg_file[5414] <= 8'h00
            reg_file[5415] <= 8'h00
            reg_file[5416] <= 8'h00
            reg_file[5417] <= 8'h00
            reg_file[5418] <= 8'h00
            reg_file[5419] <= 8'h00
            reg_file[5420] <= 8'h00
            reg_file[5421] <= 8'h00
            reg_file[5422] <= 8'h00
            reg_file[5423] <= 8'h00
            reg_file[5424] <= 8'h00
            reg_file[5425] <= 8'h00
            reg_file[5426] <= 8'h00
            reg_file[5427] <= 8'h00
            reg_file[5428] <= 8'h00
            reg_file[5429] <= 8'h00
            reg_file[5430] <= 8'h00
            reg_file[5431] <= 8'h00
            reg_file[5432] <= 8'h00
            reg_file[5433] <= 8'h00
            reg_file[5434] <= 8'h00
            reg_file[5435] <= 8'h00
            reg_file[5436] <= 8'h00
            reg_file[5437] <= 8'h00
            reg_file[5438] <= 8'h00
            reg_file[5439] <= 8'h00
            reg_file[5440] <= 8'h00
            reg_file[5441] <= 8'h00
            reg_file[5442] <= 8'h00
            reg_file[5443] <= 8'h00
            reg_file[5444] <= 8'h00
            reg_file[5445] <= 8'h00
            reg_file[5446] <= 8'h00
            reg_file[5447] <= 8'h00
            reg_file[5448] <= 8'h00
            reg_file[5449] <= 8'h00
            reg_file[5450] <= 8'h00
            reg_file[5451] <= 8'h00
            reg_file[5452] <= 8'h00
            reg_file[5453] <= 8'h00
            reg_file[5454] <= 8'h00
            reg_file[5455] <= 8'h00
            reg_file[5456] <= 8'h00
            reg_file[5457] <= 8'h00
            reg_file[5458] <= 8'h00
            reg_file[5459] <= 8'h00
            reg_file[5460] <= 8'h00
            reg_file[5461] <= 8'h00
            reg_file[5462] <= 8'h00
            reg_file[5463] <= 8'h00
            reg_file[5464] <= 8'h00
            reg_file[5465] <= 8'h00
            reg_file[5466] <= 8'h00
            reg_file[5467] <= 8'h00
            reg_file[5468] <= 8'h00
            reg_file[5469] <= 8'h00
            reg_file[5470] <= 8'h00
            reg_file[5471] <= 8'h00
            reg_file[5472] <= 8'h00
            reg_file[5473] <= 8'h00
            reg_file[5474] <= 8'h00
            reg_file[5475] <= 8'h00
            reg_file[5476] <= 8'h00
            reg_file[5477] <= 8'h00
            reg_file[5478] <= 8'h00
            reg_file[5479] <= 8'h00
            reg_file[5480] <= 8'h00
            reg_file[5481] <= 8'h00
            reg_file[5482] <= 8'h00
            reg_file[5483] <= 8'h00
            reg_file[5484] <= 8'h00
            reg_file[5485] <= 8'h00
            reg_file[5486] <= 8'h00
            reg_file[5487] <= 8'h00
            reg_file[5488] <= 8'h00
            reg_file[5489] <= 8'h00
            reg_file[5490] <= 8'h00
            reg_file[5491] <= 8'h00
            reg_file[5492] <= 8'h00
            reg_file[5493] <= 8'h00
            reg_file[5494] <= 8'h00
            reg_file[5495] <= 8'h00
            reg_file[5496] <= 8'h00
            reg_file[5497] <= 8'h00
            reg_file[5498] <= 8'h00
            reg_file[5499] <= 8'h00
            reg_file[5500] <= 8'h00
            reg_file[5501] <= 8'h00
            reg_file[5502] <= 8'h00
            reg_file[5503] <= 8'h00
            reg_file[5504] <= 8'h00
            reg_file[5505] <= 8'h00
            reg_file[5506] <= 8'h00
            reg_file[5507] <= 8'h00
            reg_file[5508] <= 8'h00
            reg_file[5509] <= 8'h00
            reg_file[5510] <= 8'h00
            reg_file[5511] <= 8'h00
            reg_file[5512] <= 8'h00
            reg_file[5513] <= 8'h00
            reg_file[5514] <= 8'h00
            reg_file[5515] <= 8'h00
            reg_file[5516] <= 8'h00
            reg_file[5517] <= 8'h00
            reg_file[5518] <= 8'h00
            reg_file[5519] <= 8'h00
            reg_file[5520] <= 8'h00
            reg_file[5521] <= 8'h00
            reg_file[5522] <= 8'h00
            reg_file[5523] <= 8'h00
            reg_file[5524] <= 8'h00
            reg_file[5525] <= 8'h00
            reg_file[5526] <= 8'h00
            reg_file[5527] <= 8'h00
            reg_file[5528] <= 8'h00
            reg_file[5529] <= 8'h00
            reg_file[5530] <= 8'h00
            reg_file[5531] <= 8'h00
            reg_file[5532] <= 8'h00
            reg_file[5533] <= 8'h00
            reg_file[5534] <= 8'h00
            reg_file[5535] <= 8'h00
            reg_file[5536] <= 8'h00
            reg_file[5537] <= 8'h00
            reg_file[5538] <= 8'h00
            reg_file[5539] <= 8'h00
            reg_file[5540] <= 8'h00
            reg_file[5541] <= 8'h00
            reg_file[5542] <= 8'h00
            reg_file[5543] <= 8'h00
            reg_file[5544] <= 8'h00
            reg_file[5545] <= 8'h00
            reg_file[5546] <= 8'h00
            reg_file[5547] <= 8'h00
            reg_file[5548] <= 8'h00
            reg_file[5549] <= 8'h00
            reg_file[5550] <= 8'h00
            reg_file[5551] <= 8'h00
            reg_file[5552] <= 8'h00
            reg_file[5553] <= 8'h00
            reg_file[5554] <= 8'h00
            reg_file[5555] <= 8'h00
            reg_file[5556] <= 8'h00
            reg_file[5557] <= 8'h00
            reg_file[5558] <= 8'h00
            reg_file[5559] <= 8'h00
            reg_file[5560] <= 8'h00
            reg_file[5561] <= 8'h00
            reg_file[5562] <= 8'h00
            reg_file[5563] <= 8'h00
            reg_file[5564] <= 8'h00
            reg_file[5565] <= 8'h00
            reg_file[5566] <= 8'h00
            reg_file[5567] <= 8'h00
            reg_file[5568] <= 8'h00
            reg_file[5569] <= 8'h00
            reg_file[5570] <= 8'h00
            reg_file[5571] <= 8'h00
            reg_file[5572] <= 8'h00
            reg_file[5573] <= 8'h00
            reg_file[5574] <= 8'h00
            reg_file[5575] <= 8'h00
            reg_file[5576] <= 8'h00
            reg_file[5577] <= 8'h00
            reg_file[5578] <= 8'h00
            reg_file[5579] <= 8'h00
            reg_file[5580] <= 8'h00
            reg_file[5581] <= 8'h00
            reg_file[5582] <= 8'h00
            reg_file[5583] <= 8'h00
            reg_file[5584] <= 8'h00
            reg_file[5585] <= 8'h00
            reg_file[5586] <= 8'h00
            reg_file[5587] <= 8'h00
            reg_file[5588] <= 8'h00
            reg_file[5589] <= 8'h00
            reg_file[5590] <= 8'h00
            reg_file[5591] <= 8'h00
            reg_file[5592] <= 8'h00
            reg_file[5593] <= 8'h00
            reg_file[5594] <= 8'h00
            reg_file[5595] <= 8'h00
            reg_file[5596] <= 8'h00
            reg_file[5597] <= 8'h00
            reg_file[5598] <= 8'h00
            reg_file[5599] <= 8'h00
            reg_file[5600] <= 8'h00
            reg_file[5601] <= 8'h00
            reg_file[5602] <= 8'h00
            reg_file[5603] <= 8'h00
            reg_file[5604] <= 8'h00
            reg_file[5605] <= 8'h00
            reg_file[5606] <= 8'h00
            reg_file[5607] <= 8'h00
            reg_file[5608] <= 8'h00
            reg_file[5609] <= 8'h00
            reg_file[5610] <= 8'h00
            reg_file[5611] <= 8'h00
            reg_file[5612] <= 8'h00
            reg_file[5613] <= 8'h00
            reg_file[5614] <= 8'h00
            reg_file[5615] <= 8'h00
            reg_file[5616] <= 8'h00
            reg_file[5617] <= 8'h00
            reg_file[5618] <= 8'h00
            reg_file[5619] <= 8'h00
            reg_file[5620] <= 8'h00
            reg_file[5621] <= 8'h00
            reg_file[5622] <= 8'h00
            reg_file[5623] <= 8'h00
            reg_file[5624] <= 8'h00
            reg_file[5625] <= 8'h00
            reg_file[5626] <= 8'h00
            reg_file[5627] <= 8'h00
            reg_file[5628] <= 8'h00
            reg_file[5629] <= 8'h00
            reg_file[5630] <= 8'h00
            reg_file[5631] <= 8'h00
            reg_file[5632] <= 8'h00
            reg_file[5633] <= 8'h00
            reg_file[5634] <= 8'h00
            reg_file[5635] <= 8'h00
            reg_file[5636] <= 8'h00
            reg_file[5637] <= 8'h00
            reg_file[5638] <= 8'h00
            reg_file[5639] <= 8'h00
            reg_file[5640] <= 8'h00
            reg_file[5641] <= 8'h00
            reg_file[5642] <= 8'h00
            reg_file[5643] <= 8'h00
            reg_file[5644] <= 8'h00
            reg_file[5645] <= 8'h00
            reg_file[5646] <= 8'h00
            reg_file[5647] <= 8'h00
            reg_file[5648] <= 8'h00
            reg_file[5649] <= 8'h00
            reg_file[5650] <= 8'h00
            reg_file[5651] <= 8'h00
            reg_file[5652] <= 8'h00
            reg_file[5653] <= 8'h00
            reg_file[5654] <= 8'h00
            reg_file[5655] <= 8'h00
            reg_file[5656] <= 8'h00
            reg_file[5657] <= 8'h00
            reg_file[5658] <= 8'h00
            reg_file[5659] <= 8'h00
            reg_file[5660] <= 8'h00
            reg_file[5661] <= 8'h00
            reg_file[5662] <= 8'h00
            reg_file[5663] <= 8'h00
            reg_file[5664] <= 8'h00
            reg_file[5665] <= 8'h00
            reg_file[5666] <= 8'h00
            reg_file[5667] <= 8'h00
            reg_file[5668] <= 8'h00
            reg_file[5669] <= 8'h00
            reg_file[5670] <= 8'h00
            reg_file[5671] <= 8'h00
            reg_file[5672] <= 8'h00
            reg_file[5673] <= 8'h00
            reg_file[5674] <= 8'h00
            reg_file[5675] <= 8'h00
            reg_file[5676] <= 8'h00
            reg_file[5677] <= 8'h00
            reg_file[5678] <= 8'h00
            reg_file[5679] <= 8'h00
            reg_file[5680] <= 8'h00
            reg_file[5681] <= 8'h00
            reg_file[5682] <= 8'h00
            reg_file[5683] <= 8'h00
            reg_file[5684] <= 8'h00
            reg_file[5685] <= 8'h00
            reg_file[5686] <= 8'h00
            reg_file[5687] <= 8'h00
            reg_file[5688] <= 8'h00
            reg_file[5689] <= 8'h00
            reg_file[5690] <= 8'h00
            reg_file[5691] <= 8'h00
            reg_file[5692] <= 8'h00
            reg_file[5693] <= 8'h00
            reg_file[5694] <= 8'h00
            reg_file[5695] <= 8'h00
            reg_file[5696] <= 8'h00
            reg_file[5697] <= 8'h00
            reg_file[5698] <= 8'h00
            reg_file[5699] <= 8'h00
            reg_file[5700] <= 8'h00
            reg_file[5701] <= 8'h00
            reg_file[5702] <= 8'h00
            reg_file[5703] <= 8'h00
            reg_file[5704] <= 8'h00
            reg_file[5705] <= 8'h00
            reg_file[5706] <= 8'h00
            reg_file[5707] <= 8'h00
            reg_file[5708] <= 8'h00
            reg_file[5709] <= 8'h00
            reg_file[5710] <= 8'h00
            reg_file[5711] <= 8'h00
            reg_file[5712] <= 8'h00
            reg_file[5713] <= 8'h00
            reg_file[5714] <= 8'h00
            reg_file[5715] <= 8'h00
            reg_file[5716] <= 8'h00
            reg_file[5717] <= 8'h00
            reg_file[5718] <= 8'h00
            reg_file[5719] <= 8'h00
            reg_file[5720] <= 8'h00
            reg_file[5721] <= 8'h00
            reg_file[5722] <= 8'h00
            reg_file[5723] <= 8'h00
            reg_file[5724] <= 8'h00
            reg_file[5725] <= 8'h00
            reg_file[5726] <= 8'h00
            reg_file[5727] <= 8'h00
            reg_file[5728] <= 8'h00
            reg_file[5729] <= 8'h00
            reg_file[5730] <= 8'h00
            reg_file[5731] <= 8'h00
            reg_file[5732] <= 8'h00
            reg_file[5733] <= 8'h00
            reg_file[5734] <= 8'h00
            reg_file[5735] <= 8'h00
            reg_file[5736] <= 8'h00
            reg_file[5737] <= 8'h00
            reg_file[5738] <= 8'h00
            reg_file[5739] <= 8'h00
            reg_file[5740] <= 8'h00
            reg_file[5741] <= 8'h00
            reg_file[5742] <= 8'h00
            reg_file[5743] <= 8'h00
            reg_file[5744] <= 8'h00
            reg_file[5745] <= 8'h00
            reg_file[5746] <= 8'h00
            reg_file[5747] <= 8'h00
            reg_file[5748] <= 8'h00
            reg_file[5749] <= 8'h00
            reg_file[5750] <= 8'h00
            reg_file[5751] <= 8'h00
            reg_file[5752] <= 8'h00
            reg_file[5753] <= 8'h00
            reg_file[5754] <= 8'h00
            reg_file[5755] <= 8'h00
            reg_file[5756] <= 8'h00
            reg_file[5757] <= 8'h00
            reg_file[5758] <= 8'h00
            reg_file[5759] <= 8'h00
            reg_file[5760] <= 8'h00
            reg_file[5761] <= 8'h00
            reg_file[5762] <= 8'h00
            reg_file[5763] <= 8'h00
            reg_file[5764] <= 8'h00
            reg_file[5765] <= 8'h00
            reg_file[5766] <= 8'h00
            reg_file[5767] <= 8'h00
            reg_file[5768] <= 8'h00
            reg_file[5769] <= 8'h00
            reg_file[5770] <= 8'h00
            reg_file[5771] <= 8'h00
            reg_file[5772] <= 8'h00
            reg_file[5773] <= 8'h00
            reg_file[5774] <= 8'h00
            reg_file[5775] <= 8'h00
            reg_file[5776] <= 8'h00
            reg_file[5777] <= 8'h00
            reg_file[5778] <= 8'h00
            reg_file[5779] <= 8'h00
            reg_file[5780] <= 8'h00
            reg_file[5781] <= 8'h00
            reg_file[5782] <= 8'h00
            reg_file[5783] <= 8'h00
            reg_file[5784] <= 8'h00
            reg_file[5785] <= 8'h00
            reg_file[5786] <= 8'h00
            reg_file[5787] <= 8'h00
            reg_file[5788] <= 8'h00
            reg_file[5789] <= 8'h00
            reg_file[5790] <= 8'h00
            reg_file[5791] <= 8'h00
            reg_file[5792] <= 8'h00
            reg_file[5793] <= 8'h00
            reg_file[5794] <= 8'h00
            reg_file[5795] <= 8'h00
            reg_file[5796] <= 8'h00
            reg_file[5797] <= 8'h00
            reg_file[5798] <= 8'h00
            reg_file[5799] <= 8'h00
            reg_file[5800] <= 8'h00
            reg_file[5801] <= 8'h00
            reg_file[5802] <= 8'h00
            reg_file[5803] <= 8'h00
            reg_file[5804] <= 8'h00
            reg_file[5805] <= 8'h00
            reg_file[5806] <= 8'h00
            reg_file[5807] <= 8'h00
            reg_file[5808] <= 8'h00
            reg_file[5809] <= 8'h00
            reg_file[5810] <= 8'h00
            reg_file[5811] <= 8'h00
            reg_file[5812] <= 8'h00
            reg_file[5813] <= 8'h00
            reg_file[5814] <= 8'h00
            reg_file[5815] <= 8'h00
            reg_file[5816] <= 8'h00
            reg_file[5817] <= 8'h00
            reg_file[5818] <= 8'h00
            reg_file[5819] <= 8'h00
            reg_file[5820] <= 8'h00
            reg_file[5821] <= 8'h00
            reg_file[5822] <= 8'h00
            reg_file[5823] <= 8'h00
            reg_file[5824] <= 8'h00
            reg_file[5825] <= 8'h00
            reg_file[5826] <= 8'h00
            reg_file[5827] <= 8'h00
            reg_file[5828] <= 8'h00
            reg_file[5829] <= 8'h00
            reg_file[5830] <= 8'h00
            reg_file[5831] <= 8'h00
            reg_file[5832] <= 8'h00
            reg_file[5833] <= 8'h00
            reg_file[5834] <= 8'h00
            reg_file[5835] <= 8'h00
            reg_file[5836] <= 8'h00
            reg_file[5837] <= 8'h00
            reg_file[5838] <= 8'h00
            reg_file[5839] <= 8'h00
            reg_file[5840] <= 8'h00
            reg_file[5841] <= 8'h00
            reg_file[5842] <= 8'h00
            reg_file[5843] <= 8'h00
            reg_file[5844] <= 8'h00
            reg_file[5845] <= 8'h00
            reg_file[5846] <= 8'h00
            reg_file[5847] <= 8'h00
            reg_file[5848] <= 8'h00
            reg_file[5849] <= 8'h00
            reg_file[5850] <= 8'h00
            reg_file[5851] <= 8'h00
            reg_file[5852] <= 8'h00
            reg_file[5853] <= 8'h00
            reg_file[5854] <= 8'h00
            reg_file[5855] <= 8'h00
            reg_file[5856] <= 8'h00
            reg_file[5857] <= 8'h00
            reg_file[5858] <= 8'h00
            reg_file[5859] <= 8'h00
            reg_file[5860] <= 8'h00
            reg_file[5861] <= 8'h00
            reg_file[5862] <= 8'h00
            reg_file[5863] <= 8'h00
            reg_file[5864] <= 8'h00
            reg_file[5865] <= 8'h00
            reg_file[5866] <= 8'h00
            reg_file[5867] <= 8'h00
            reg_file[5868] <= 8'h00
            reg_file[5869] <= 8'h00
            reg_file[5870] <= 8'h00
            reg_file[5871] <= 8'h00
            reg_file[5872] <= 8'h00
            reg_file[5873] <= 8'h00
            reg_file[5874] <= 8'h00
            reg_file[5875] <= 8'h00
            reg_file[5876] <= 8'h00
            reg_file[5877] <= 8'h00
            reg_file[5878] <= 8'h00
            reg_file[5879] <= 8'h00
            reg_file[5880] <= 8'h00
            reg_file[5881] <= 8'h00
            reg_file[5882] <= 8'h00
            reg_file[5883] <= 8'h00
            reg_file[5884] <= 8'h00
            reg_file[5885] <= 8'h00
            reg_file[5886] <= 8'h00
            reg_file[5887] <= 8'h00
            reg_file[5888] <= 8'h00
            reg_file[5889] <= 8'h00
            reg_file[5890] <= 8'h00
            reg_file[5891] <= 8'h00
            reg_file[5892] <= 8'h00
            reg_file[5893] <= 8'h00
            reg_file[5894] <= 8'h00
            reg_file[5895] <= 8'h00
            reg_file[5896] <= 8'h00
            reg_file[5897] <= 8'h00
            reg_file[5898] <= 8'h00
            reg_file[5899] <= 8'h00
            reg_file[5900] <= 8'h00
            reg_file[5901] <= 8'h00
            reg_file[5902] <= 8'h00
            reg_file[5903] <= 8'h00
            reg_file[5904] <= 8'h00
            reg_file[5905] <= 8'h00
            reg_file[5906] <= 8'h00
            reg_file[5907] <= 8'h00
            reg_file[5908] <= 8'h00
            reg_file[5909] <= 8'h00
            reg_file[5910] <= 8'h00
            reg_file[5911] <= 8'h00
            reg_file[5912] <= 8'h00
            reg_file[5913] <= 8'h00
            reg_file[5914] <= 8'h00
            reg_file[5915] <= 8'h00
            reg_file[5916] <= 8'h00
            reg_file[5917] <= 8'h00
            reg_file[5918] <= 8'h00
            reg_file[5919] <= 8'h00
            reg_file[5920] <= 8'h00
            reg_file[5921] <= 8'h00
            reg_file[5922] <= 8'h00
            reg_file[5923] <= 8'h00
            reg_file[5924] <= 8'h00
            reg_file[5925] <= 8'h00
            reg_file[5926] <= 8'h00
            reg_file[5927] <= 8'h00
            reg_file[5928] <= 8'h00
            reg_file[5929] <= 8'h00
            reg_file[5930] <= 8'h00
            reg_file[5931] <= 8'h00
            reg_file[5932] <= 8'h00
            reg_file[5933] <= 8'h00
            reg_file[5934] <= 8'h00
            reg_file[5935] <= 8'h00
            reg_file[5936] <= 8'h00
            reg_file[5937] <= 8'h00
            reg_file[5938] <= 8'h00
            reg_file[5939] <= 8'h00
            reg_file[5940] <= 8'h00
            reg_file[5941] <= 8'h00
            reg_file[5942] <= 8'h00
            reg_file[5943] <= 8'h00
            reg_file[5944] <= 8'h00
            reg_file[5945] <= 8'h00
            reg_file[5946] <= 8'h00
            reg_file[5947] <= 8'h00
            reg_file[5948] <= 8'h00
            reg_file[5949] <= 8'h00
            reg_file[5950] <= 8'h00
            reg_file[5951] <= 8'h00
            reg_file[5952] <= 8'h00
            reg_file[5953] <= 8'h00
            reg_file[5954] <= 8'h00
            reg_file[5955] <= 8'h00
            reg_file[5956] <= 8'h00
            reg_file[5957] <= 8'h00
            reg_file[5958] <= 8'h00
            reg_file[5959] <= 8'h00
            reg_file[5960] <= 8'h00
            reg_file[5961] <= 8'h00
            reg_file[5962] <= 8'h00
            reg_file[5963] <= 8'h00
            reg_file[5964] <= 8'h00
            reg_file[5965] <= 8'h00
            reg_file[5966] <= 8'h00
            reg_file[5967] <= 8'h00
            reg_file[5968] <= 8'h00
            reg_file[5969] <= 8'h00
            reg_file[5970] <= 8'h00
            reg_file[5971] <= 8'h00
            reg_file[5972] <= 8'h00
            reg_file[5973] <= 8'h00
            reg_file[5974] <= 8'h00
            reg_file[5975] <= 8'h00
            reg_file[5976] <= 8'h00
            reg_file[5977] <= 8'h00
            reg_file[5978] <= 8'h00
            reg_file[5979] <= 8'h00
            reg_file[5980] <= 8'h00
            reg_file[5981] <= 8'h00
            reg_file[5982] <= 8'h00
            reg_file[5983] <= 8'h00
            reg_file[5984] <= 8'h00
            reg_file[5985] <= 8'h00
            reg_file[5986] <= 8'h00
            reg_file[5987] <= 8'h00
            reg_file[5988] <= 8'h00
            reg_file[5989] <= 8'h00
            reg_file[5990] <= 8'h00
            reg_file[5991] <= 8'h00
            reg_file[5992] <= 8'h00
            reg_file[5993] <= 8'h00
            reg_file[5994] <= 8'h00
            reg_file[5995] <= 8'h00
            reg_file[5996] <= 8'h00
            reg_file[5997] <= 8'h00
            reg_file[5998] <= 8'h00
            reg_file[5999] <= 8'h00
            reg_file[6000] <= 8'h00
            reg_file[6001] <= 8'h00
            reg_file[6002] <= 8'h00
            reg_file[6003] <= 8'h00
            reg_file[6004] <= 8'h00
            reg_file[6005] <= 8'h00
            reg_file[6006] <= 8'h00
            reg_file[6007] <= 8'h00
            reg_file[6008] <= 8'h00
            reg_file[6009] <= 8'h00
            reg_file[6010] <= 8'h00
            reg_file[6011] <= 8'h00
            reg_file[6012] <= 8'h00
            reg_file[6013] <= 8'h00
            reg_file[6014] <= 8'h00
            reg_file[6015] <= 8'h00
            reg_file[6016] <= 8'h00
            reg_file[6017] <= 8'h00
            reg_file[6018] <= 8'h00
            reg_file[6019] <= 8'h00
            reg_file[6020] <= 8'h00
            reg_file[6021] <= 8'h00
            reg_file[6022] <= 8'h00
            reg_file[6023] <= 8'h00
            reg_file[6024] <= 8'h00
            reg_file[6025] <= 8'h00
            reg_file[6026] <= 8'h00
            reg_file[6027] <= 8'h00
            reg_file[6028] <= 8'h00
            reg_file[6029] <= 8'h00
            reg_file[6030] <= 8'h00
            reg_file[6031] <= 8'h00
            reg_file[6032] <= 8'h00
            reg_file[6033] <= 8'h00
            reg_file[6034] <= 8'h00
            reg_file[6035] <= 8'h00
            reg_file[6036] <= 8'h00
            reg_file[6037] <= 8'h00
            reg_file[6038] <= 8'h00
            reg_file[6039] <= 8'h00
            reg_file[6040] <= 8'h00
            reg_file[6041] <= 8'h00
            reg_file[6042] <= 8'h00
            reg_file[6043] <= 8'h00
            reg_file[6044] <= 8'h00
            reg_file[6045] <= 8'h00
            reg_file[6046] <= 8'h00
            reg_file[6047] <= 8'h00
            reg_file[6048] <= 8'h00
            reg_file[6049] <= 8'h00
            reg_file[6050] <= 8'h00
            reg_file[6051] <= 8'h00
            reg_file[6052] <= 8'h00
            reg_file[6053] <= 8'h00
            reg_file[6054] <= 8'h00
            reg_file[6055] <= 8'h00
            reg_file[6056] <= 8'h00
            reg_file[6057] <= 8'h00
            reg_file[6058] <= 8'h00
            reg_file[6059] <= 8'h00
            reg_file[6060] <= 8'h00
            reg_file[6061] <= 8'h00
            reg_file[6062] <= 8'h00
            reg_file[6063] <= 8'h00
            reg_file[6064] <= 8'h00
            reg_file[6065] <= 8'h00
            reg_file[6066] <= 8'h00
            reg_file[6067] <= 8'h00
            reg_file[6068] <= 8'h00
            reg_file[6069] <= 8'h00
            reg_file[6070] <= 8'h00
            reg_file[6071] <= 8'h00
            reg_file[6072] <= 8'h00
            reg_file[6073] <= 8'h00
            reg_file[6074] <= 8'h00
            reg_file[6075] <= 8'h00
            reg_file[6076] <= 8'h00
            reg_file[6077] <= 8'h00
            reg_file[6078] <= 8'h00
            reg_file[6079] <= 8'h00
            reg_file[6080] <= 8'h00
            reg_file[6081] <= 8'h00
            reg_file[6082] <= 8'h00
            reg_file[6083] <= 8'h00
            reg_file[6084] <= 8'h00
            reg_file[6085] <= 8'h00
            reg_file[6086] <= 8'h00
            reg_file[6087] <= 8'h00
            reg_file[6088] <= 8'h00
            reg_file[6089] <= 8'h00
            reg_file[6090] <= 8'h00
            reg_file[6091] <= 8'h00
            reg_file[6092] <= 8'h00
            reg_file[6093] <= 8'h00
            reg_file[6094] <= 8'h00
            reg_file[6095] <= 8'h00
            reg_file[6096] <= 8'h00
            reg_file[6097] <= 8'h00
            reg_file[6098] <= 8'h00
            reg_file[6099] <= 8'h00
            reg_file[6100] <= 8'h00
            reg_file[6101] <= 8'h00
            reg_file[6102] <= 8'h00
            reg_file[6103] <= 8'h00
            reg_file[6104] <= 8'h00
            reg_file[6105] <= 8'h00
            reg_file[6106] <= 8'h00
            reg_file[6107] <= 8'h00
            reg_file[6108] <= 8'h00
            reg_file[6109] <= 8'h00
            reg_file[6110] <= 8'h00
            reg_file[6111] <= 8'h00
            reg_file[6112] <= 8'h00
            reg_file[6113] <= 8'h00
            reg_file[6114] <= 8'h00
            reg_file[6115] <= 8'h00
            reg_file[6116] <= 8'h00
            reg_file[6117] <= 8'h00
            reg_file[6118] <= 8'h00
            reg_file[6119] <= 8'h00
            reg_file[6120] <= 8'h00
            reg_file[6121] <= 8'h00
            reg_file[6122] <= 8'h00
            reg_file[6123] <= 8'h00
            reg_file[6124] <= 8'h00
            reg_file[6125] <= 8'h00
            reg_file[6126] <= 8'h00
            reg_file[6127] <= 8'h00
            reg_file[6128] <= 8'h00
            reg_file[6129] <= 8'h00
            reg_file[6130] <= 8'h00
            reg_file[6131] <= 8'h00
            reg_file[6132] <= 8'h00
            reg_file[6133] <= 8'h00
            reg_file[6134] <= 8'h00
            reg_file[6135] <= 8'h00
            reg_file[6136] <= 8'h00
            reg_file[6137] <= 8'h00
            reg_file[6138] <= 8'h00
            reg_file[6139] <= 8'h00
            reg_file[6140] <= 8'h00
            reg_file[6141] <= 8'h00
            reg_file[6142] <= 8'h00
            reg_file[6143] <= 8'h00
            reg_file[6144] <= 8'h00
            reg_file[6145] <= 8'h00
            reg_file[6146] <= 8'h00
            reg_file[6147] <= 8'h00
            reg_file[6148] <= 8'h00
            reg_file[6149] <= 8'h00
            reg_file[6150] <= 8'h00
            reg_file[6151] <= 8'h00
            reg_file[6152] <= 8'h00
            reg_file[6153] <= 8'h00
            reg_file[6154] <= 8'h00
            reg_file[6155] <= 8'h00
            reg_file[6156] <= 8'h00
            reg_file[6157] <= 8'h00
            reg_file[6158] <= 8'h00
            reg_file[6159] <= 8'h00
            reg_file[6160] <= 8'h00
            reg_file[6161] <= 8'h00
            reg_file[6162] <= 8'h00
            reg_file[6163] <= 8'h00
            reg_file[6164] <= 8'h00
            reg_file[6165] <= 8'h00
            reg_file[6166] <= 8'h00
            reg_file[6167] <= 8'h00
            reg_file[6168] <= 8'h00
            reg_file[6169] <= 8'h00
            reg_file[6170] <= 8'h00
            reg_file[6171] <= 8'h00
            reg_file[6172] <= 8'h00
            reg_file[6173] <= 8'h00
            reg_file[6174] <= 8'h00
            reg_file[6175] <= 8'h00
            reg_file[6176] <= 8'h00
            reg_file[6177] <= 8'h00
            reg_file[6178] <= 8'h00
            reg_file[6179] <= 8'h00
            reg_file[6180] <= 8'h00
            reg_file[6181] <= 8'h00
            reg_file[6182] <= 8'h00
            reg_file[6183] <= 8'h00
            reg_file[6184] <= 8'h00
            reg_file[6185] <= 8'h00
            reg_file[6186] <= 8'h00
            reg_file[6187] <= 8'h00
            reg_file[6188] <= 8'h00
            reg_file[6189] <= 8'h00
            reg_file[6190] <= 8'h00
            reg_file[6191] <= 8'h00
            reg_file[6192] <= 8'h00
            reg_file[6193] <= 8'h00
            reg_file[6194] <= 8'h00
            reg_file[6195] <= 8'h00
            reg_file[6196] <= 8'h00
            reg_file[6197] <= 8'h00
            reg_file[6198] <= 8'h00
            reg_file[6199] <= 8'h00
            reg_file[6200] <= 8'h00
            reg_file[6201] <= 8'h00
            reg_file[6202] <= 8'h00
            reg_file[6203] <= 8'h00
            reg_file[6204] <= 8'h00
            reg_file[6205] <= 8'h00
            reg_file[6206] <= 8'h00
            reg_file[6207] <= 8'h00
            reg_file[6208] <= 8'h00
            reg_file[6209] <= 8'h00
            reg_file[6210] <= 8'h00
            reg_file[6211] <= 8'h00
            reg_file[6212] <= 8'h00
            reg_file[6213] <= 8'h00
            reg_file[6214] <= 8'h00
            reg_file[6215] <= 8'h00
            reg_file[6216] <= 8'h00
            reg_file[6217] <= 8'h00
            reg_file[6218] <= 8'h00
            reg_file[6219] <= 8'h00
            reg_file[6220] <= 8'h00
            reg_file[6221] <= 8'h00
            reg_file[6222] <= 8'h00
            reg_file[6223] <= 8'h00
            reg_file[6224] <= 8'h00
            reg_file[6225] <= 8'h00
            reg_file[6226] <= 8'h00
            reg_file[6227] <= 8'h00
            reg_file[6228] <= 8'h00
            reg_file[6229] <= 8'h00
            reg_file[6230] <= 8'h00
            reg_file[6231] <= 8'h00
            reg_file[6232] <= 8'h00
            reg_file[6233] <= 8'h00
            reg_file[6234] <= 8'h00
            reg_file[6235] <= 8'h00
            reg_file[6236] <= 8'h00
            reg_file[6237] <= 8'h00
            reg_file[6238] <= 8'h00
            reg_file[6239] <= 8'h00
            reg_file[6240] <= 8'h00
            reg_file[6241] <= 8'h00
            reg_file[6242] <= 8'h00
            reg_file[6243] <= 8'h00
            reg_file[6244] <= 8'h00
            reg_file[6245] <= 8'h00
            reg_file[6246] <= 8'h00
            reg_file[6247] <= 8'h00
            reg_file[6248] <= 8'h00
            reg_file[6249] <= 8'h00
            reg_file[6250] <= 8'h00
            reg_file[6251] <= 8'h00
            reg_file[6252] <= 8'h00
            reg_file[6253] <= 8'h00
            reg_file[6254] <= 8'h00
            reg_file[6255] <= 8'h00
            reg_file[6256] <= 8'h00
            reg_file[6257] <= 8'h00
            reg_file[6258] <= 8'h00
            reg_file[6259] <= 8'h00
            reg_file[6260] <= 8'h00
            reg_file[6261] <= 8'h00
            reg_file[6262] <= 8'h00
            reg_file[6263] <= 8'h00
            reg_file[6264] <= 8'h00
            reg_file[6265] <= 8'h00
            reg_file[6266] <= 8'h00
            reg_file[6267] <= 8'h00
            reg_file[6268] <= 8'h00
            reg_file[6269] <= 8'h00
            reg_file[6270] <= 8'h00
            reg_file[6271] <= 8'h00
            reg_file[6272] <= 8'h00
            reg_file[6273] <= 8'h00
            reg_file[6274] <= 8'h00
            reg_file[6275] <= 8'h00
            reg_file[6276] <= 8'h00
            reg_file[6277] <= 8'h00
            reg_file[6278] <= 8'h00
            reg_file[6279] <= 8'h00
            reg_file[6280] <= 8'h00
            reg_file[6281] <= 8'h00
            reg_file[6282] <= 8'h00
            reg_file[6283] <= 8'h00
            reg_file[6284] <= 8'h00
            reg_file[6285] <= 8'h00
            reg_file[6286] <= 8'h00
            reg_file[6287] <= 8'h00
            reg_file[6288] <= 8'h00
            reg_file[6289] <= 8'h00
            reg_file[6290] <= 8'h00
            reg_file[6291] <= 8'h00
            reg_file[6292] <= 8'h00
            reg_file[6293] <= 8'h00
            reg_file[6294] <= 8'h00
            reg_file[6295] <= 8'h00
            reg_file[6296] <= 8'h00
            reg_file[6297] <= 8'h00
            reg_file[6298] <= 8'h00
            reg_file[6299] <= 8'h00
            reg_file[6300] <= 8'h00
            reg_file[6301] <= 8'h00
            reg_file[6302] <= 8'h00
            reg_file[6303] <= 8'h00
            reg_file[6304] <= 8'h00
            reg_file[6305] <= 8'h00
            reg_file[6306] <= 8'h00
            reg_file[6307] <= 8'h00
            reg_file[6308] <= 8'h00
            reg_file[6309] <= 8'h00
            reg_file[6310] <= 8'h00
            reg_file[6311] <= 8'h00
            reg_file[6312] <= 8'h00
            reg_file[6313] <= 8'h00
            reg_file[6314] <= 8'h00
            reg_file[6315] <= 8'h00
            reg_file[6316] <= 8'h00
            reg_file[6317] <= 8'h00
            reg_file[6318] <= 8'h00
            reg_file[6319] <= 8'h00
            reg_file[6320] <= 8'h00
            reg_file[6321] <= 8'h00
            reg_file[6322] <= 8'h00
            reg_file[6323] <= 8'h00
            reg_file[6324] <= 8'h00
            reg_file[6325] <= 8'h00
            reg_file[6326] <= 8'h00
            reg_file[6327] <= 8'h00
            reg_file[6328] <= 8'h00
            reg_file[6329] <= 8'h00
            reg_file[6330] <= 8'h00
            reg_file[6331] <= 8'h00
            reg_file[6332] <= 8'h00
            reg_file[6333] <= 8'h00
            reg_file[6334] <= 8'h00
            reg_file[6335] <= 8'h00
            reg_file[6336] <= 8'h00
            reg_file[6337] <= 8'h00
            reg_file[6338] <= 8'h00
            reg_file[6339] <= 8'h00
            reg_file[6340] <= 8'h00
            reg_file[6341] <= 8'h00
            reg_file[6342] <= 8'h00
            reg_file[6343] <= 8'h00
            reg_file[6344] <= 8'h00
            reg_file[6345] <= 8'h00
            reg_file[6346] <= 8'h00
            reg_file[6347] <= 8'h00
            reg_file[6348] <= 8'h00
            reg_file[6349] <= 8'h00
            reg_file[6350] <= 8'h00
            reg_file[6351] <= 8'h00
            reg_file[6352] <= 8'h00
            reg_file[6353] <= 8'h00
            reg_file[6354] <= 8'h00
            reg_file[6355] <= 8'h00
            reg_file[6356] <= 8'h00
            reg_file[6357] <= 8'h00
            reg_file[6358] <= 8'h00
            reg_file[6359] <= 8'h00
            reg_file[6360] <= 8'h00
            reg_file[6361] <= 8'h00
            reg_file[6362] <= 8'h00
            reg_file[6363] <= 8'h00
            reg_file[6364] <= 8'h00
            reg_file[6365] <= 8'h00
            reg_file[6366] <= 8'h00
            reg_file[6367] <= 8'h00
            reg_file[6368] <= 8'h00
            reg_file[6369] <= 8'h00
            reg_file[6370] <= 8'h00
            reg_file[6371] <= 8'h00
            reg_file[6372] <= 8'h00
            reg_file[6373] <= 8'h00
            reg_file[6374] <= 8'h00
            reg_file[6375] <= 8'h00
            reg_file[6376] <= 8'h00
            reg_file[6377] <= 8'h00
            reg_file[6378] <= 8'h00
            reg_file[6379] <= 8'h00
            reg_file[6380] <= 8'h00
            reg_file[6381] <= 8'h00
            reg_file[6382] <= 8'h00
            reg_file[6383] <= 8'h00
            reg_file[6384] <= 8'h00
            reg_file[6385] <= 8'h00
            reg_file[6386] <= 8'h00
            reg_file[6387] <= 8'h00
            reg_file[6388] <= 8'h00
            reg_file[6389] <= 8'h00
            reg_file[6390] <= 8'h00
            reg_file[6391] <= 8'h00
            reg_file[6392] <= 8'h00
            reg_file[6393] <= 8'h00
            reg_file[6394] <= 8'h00
            reg_file[6395] <= 8'h00
            reg_file[6396] <= 8'h00
            reg_file[6397] <= 8'h00
            reg_file[6398] <= 8'h00
            reg_file[6399] <= 8'h00
            reg_file[6400] <= 8'h00
            reg_file[6401] <= 8'h00
            reg_file[6402] <= 8'h00
            reg_file[6403] <= 8'h00
            reg_file[6404] <= 8'h00
            reg_file[6405] <= 8'h00
            reg_file[6406] <= 8'h00
            reg_file[6407] <= 8'h00
            reg_file[6408] <= 8'h00
            reg_file[6409] <= 8'h00
            reg_file[6410] <= 8'h00
            reg_file[6411] <= 8'h00
            reg_file[6412] <= 8'h00
            reg_file[6413] <= 8'h00
            reg_file[6414] <= 8'h00
            reg_file[6415] <= 8'h00
            reg_file[6416] <= 8'h00
            reg_file[6417] <= 8'h00
            reg_file[6418] <= 8'h00
            reg_file[6419] <= 8'h00
            reg_file[6420] <= 8'h00
            reg_file[6421] <= 8'h00
            reg_file[6422] <= 8'h00
            reg_file[6423] <= 8'h00
            reg_file[6424] <= 8'h00
            reg_file[6425] <= 8'h00
            reg_file[6426] <= 8'h00
            reg_file[6427] <= 8'h00
            reg_file[6428] <= 8'h00
            reg_file[6429] <= 8'h00
            reg_file[6430] <= 8'h00
            reg_file[6431] <= 8'h00
            reg_file[6432] <= 8'h00
            reg_file[6433] <= 8'h00
            reg_file[6434] <= 8'h00
            reg_file[6435] <= 8'h00
            reg_file[6436] <= 8'h00
            reg_file[6437] <= 8'h00
            reg_file[6438] <= 8'h00
            reg_file[6439] <= 8'h00
            reg_file[6440] <= 8'h00
            reg_file[6441] <= 8'h00
            reg_file[6442] <= 8'h00
            reg_file[6443] <= 8'h00
            reg_file[6444] <= 8'h00
            reg_file[6445] <= 8'h00
            reg_file[6446] <= 8'h00
            reg_file[6447] <= 8'h00
            reg_file[6448] <= 8'h00
            reg_file[6449] <= 8'h00
            reg_file[6450] <= 8'h00
            reg_file[6451] <= 8'h00
            reg_file[6452] <= 8'h00
            reg_file[6453] <= 8'h00
            reg_file[6454] <= 8'h00
            reg_file[6455] <= 8'h00
            reg_file[6456] <= 8'h00
            reg_file[6457] <= 8'h00
            reg_file[6458] <= 8'h00
            reg_file[6459] <= 8'h00
            reg_file[6460] <= 8'h00
            reg_file[6461] <= 8'h00
            reg_file[6462] <= 8'h00
            reg_file[6463] <= 8'h00
            reg_file[6464] <= 8'h00
            reg_file[6465] <= 8'h00
            reg_file[6466] <= 8'h00
            reg_file[6467] <= 8'h00
            reg_file[6468] <= 8'h00
            reg_file[6469] <= 8'h00
            reg_file[6470] <= 8'h00
            reg_file[6471] <= 8'h00
            reg_file[6472] <= 8'h00
            reg_file[6473] <= 8'h00
            reg_file[6474] <= 8'h00
            reg_file[6475] <= 8'h00
            reg_file[6476] <= 8'h00
            reg_file[6477] <= 8'h00
            reg_file[6478] <= 8'h00
            reg_file[6479] <= 8'h00
            reg_file[6480] <= 8'h00
            reg_file[6481] <= 8'h00
            reg_file[6482] <= 8'h00
            reg_file[6483] <= 8'h00
            reg_file[6484] <= 8'h00
            reg_file[6485] <= 8'h00
            reg_file[6486] <= 8'h00
            reg_file[6487] <= 8'h00
            reg_file[6488] <= 8'h00
            reg_file[6489] <= 8'h00
            reg_file[6490] <= 8'h00
            reg_file[6491] <= 8'h00
            reg_file[6492] <= 8'h00
            reg_file[6493] <= 8'h00
            reg_file[6494] <= 8'h00
            reg_file[6495] <= 8'h00
            reg_file[6496] <= 8'h00
            reg_file[6497] <= 8'h00
            reg_file[6498] <= 8'h00
            reg_file[6499] <= 8'h00
            reg_file[6500] <= 8'h00
            reg_file[6501] <= 8'h00
            reg_file[6502] <= 8'h00
            reg_file[6503] <= 8'h00
            reg_file[6504] <= 8'h00
            reg_file[6505] <= 8'h00
            reg_file[6506] <= 8'h00
            reg_file[6507] <= 8'h00
            reg_file[6508] <= 8'h00
            reg_file[6509] <= 8'h00
            reg_file[6510] <= 8'h00
            reg_file[6511] <= 8'h00
            reg_file[6512] <= 8'h00
            reg_file[6513] <= 8'h00
            reg_file[6514] <= 8'h00
            reg_file[6515] <= 8'h00
            reg_file[6516] <= 8'h00
            reg_file[6517] <= 8'h00
            reg_file[6518] <= 8'h00
            reg_file[6519] <= 8'h00
            reg_file[6520] <= 8'h00
            reg_file[6521] <= 8'h00
            reg_file[6522] <= 8'h00
            reg_file[6523] <= 8'h00
            reg_file[6524] <= 8'h00
            reg_file[6525] <= 8'h00
            reg_file[6526] <= 8'h00
            reg_file[6527] <= 8'h00
            reg_file[6528] <= 8'h00
            reg_file[6529] <= 8'h00
            reg_file[6530] <= 8'h00
            reg_file[6531] <= 8'h00
            reg_file[6532] <= 8'h00
            reg_file[6533] <= 8'h00
            reg_file[6534] <= 8'h00
            reg_file[6535] <= 8'h00
            reg_file[6536] <= 8'h00
            reg_file[6537] <= 8'h00
            reg_file[6538] <= 8'h00
            reg_file[6539] <= 8'h00
            reg_file[6540] <= 8'h00
            reg_file[6541] <= 8'h00
            reg_file[6542] <= 8'h00
            reg_file[6543] <= 8'h00
            reg_file[6544] <= 8'h00
            reg_file[6545] <= 8'h00
            reg_file[6546] <= 8'h00
            reg_file[6547] <= 8'h00
            reg_file[6548] <= 8'h00
            reg_file[6549] <= 8'h00
            reg_file[6550] <= 8'h00
            reg_file[6551] <= 8'h00
            reg_file[6552] <= 8'h00
            reg_file[6553] <= 8'h00
            reg_file[6554] <= 8'h00
            reg_file[6555] <= 8'h00
            reg_file[6556] <= 8'h00
            reg_file[6557] <= 8'h00
            reg_file[6558] <= 8'h00
            reg_file[6559] <= 8'h00
            reg_file[6560] <= 8'h00
            reg_file[6561] <= 8'h00
            reg_file[6562] <= 8'h00
            reg_file[6563] <= 8'h00
            reg_file[6564] <= 8'h00
            reg_file[6565] <= 8'h00
            reg_file[6566] <= 8'h00
            reg_file[6567] <= 8'h00
            reg_file[6568] <= 8'h00
            reg_file[6569] <= 8'h00
            reg_file[6570] <= 8'h00
            reg_file[6571] <= 8'h00
            reg_file[6572] <= 8'h00
            reg_file[6573] <= 8'h00
            reg_file[6574] <= 8'h00
            reg_file[6575] <= 8'h00
            reg_file[6576] <= 8'h00
            reg_file[6577] <= 8'h00
            reg_file[6578] <= 8'h00
            reg_file[6579] <= 8'h00
            reg_file[6580] <= 8'h00
            reg_file[6581] <= 8'h00
            reg_file[6582] <= 8'h00
            reg_file[6583] <= 8'h00
            reg_file[6584] <= 8'h00
            reg_file[6585] <= 8'h00
            reg_file[6586] <= 8'h00
            reg_file[6587] <= 8'h00
            reg_file[6588] <= 8'h00
            reg_file[6589] <= 8'h00
            reg_file[6590] <= 8'h00
            reg_file[6591] <= 8'h00
            reg_file[6592] <= 8'h00
            reg_file[6593] <= 8'h00
            reg_file[6594] <= 8'h00
            reg_file[6595] <= 8'h00
            reg_file[6596] <= 8'h00
            reg_file[6597] <= 8'h00
            reg_file[6598] <= 8'h00
            reg_file[6599] <= 8'h00
            reg_file[6600] <= 8'h00
            reg_file[6601] <= 8'h00
            reg_file[6602] <= 8'h00
            reg_file[6603] <= 8'h00
            reg_file[6604] <= 8'h00
            reg_file[6605] <= 8'h00
            reg_file[6606] <= 8'h00
            reg_file[6607] <= 8'h00
            reg_file[6608] <= 8'h00
            reg_file[6609] <= 8'h00
            reg_file[6610] <= 8'h00
            reg_file[6611] <= 8'h00
            reg_file[6612] <= 8'h00
            reg_file[6613] <= 8'h00
            reg_file[6614] <= 8'h00
            reg_file[6615] <= 8'h00
            reg_file[6616] <= 8'h00
            reg_file[6617] <= 8'h00
            reg_file[6618] <= 8'h00
            reg_file[6619] <= 8'h00
            reg_file[6620] <= 8'h00
            reg_file[6621] <= 8'h00
            reg_file[6622] <= 8'h00
            reg_file[6623] <= 8'h00
            reg_file[6624] <= 8'h00
            reg_file[6625] <= 8'h00
            reg_file[6626] <= 8'h00
            reg_file[6627] <= 8'h00
            reg_file[6628] <= 8'h00
            reg_file[6629] <= 8'h00
            reg_file[6630] <= 8'h00
            reg_file[6631] <= 8'h00
            reg_file[6632] <= 8'h00
            reg_file[6633] <= 8'h00
            reg_file[6634] <= 8'h00
            reg_file[6635] <= 8'h00
            reg_file[6636] <= 8'h00
            reg_file[6637] <= 8'h00
            reg_file[6638] <= 8'h00
            reg_file[6639] <= 8'h00
            reg_file[6640] <= 8'h00
            reg_file[6641] <= 8'h00
            reg_file[6642] <= 8'h00
            reg_file[6643] <= 8'h00
            reg_file[6644] <= 8'h00
            reg_file[6645] <= 8'h00
            reg_file[6646] <= 8'h00
            reg_file[6647] <= 8'h00
            reg_file[6648] <= 8'h00
            reg_file[6649] <= 8'h00
            reg_file[6650] <= 8'h00
            reg_file[6651] <= 8'h00
            reg_file[6652] <= 8'h00
            reg_file[6653] <= 8'h00
            reg_file[6654] <= 8'h00
            reg_file[6655] <= 8'h00
            reg_file[6656] <= 8'h00
            reg_file[6657] <= 8'h00
            reg_file[6658] <= 8'h00
            reg_file[6659] <= 8'h00
            reg_file[6660] <= 8'h00
            reg_file[6661] <= 8'h00
            reg_file[6662] <= 8'h00
            reg_file[6663] <= 8'h00
            reg_file[6664] <= 8'h00
            reg_file[6665] <= 8'h00
            reg_file[6666] <= 8'h00
            reg_file[6667] <= 8'h00
            reg_file[6668] <= 8'h00
            reg_file[6669] <= 8'h00
            reg_file[6670] <= 8'h00
            reg_file[6671] <= 8'h00
            reg_file[6672] <= 8'h00
            reg_file[6673] <= 8'h00
            reg_file[6674] <= 8'h00
            reg_file[6675] <= 8'h00
            reg_file[6676] <= 8'h00
            reg_file[6677] <= 8'h00
            reg_file[6678] <= 8'h00
            reg_file[6679] <= 8'h00
            reg_file[6680] <= 8'h00
            reg_file[6681] <= 8'h00
            reg_file[6682] <= 8'h00
            reg_file[6683] <= 8'h00
            reg_file[6684] <= 8'h00
            reg_file[6685] <= 8'h00
            reg_file[6686] <= 8'h00
            reg_file[6687] <= 8'h00
            reg_file[6688] <= 8'h00
            reg_file[6689] <= 8'h00
            reg_file[6690] <= 8'h00
            reg_file[6691] <= 8'h00
            reg_file[6692] <= 8'h00
            reg_file[6693] <= 8'h00
            reg_file[6694] <= 8'h00
            reg_file[6695] <= 8'h00
            reg_file[6696] <= 8'h00
            reg_file[6697] <= 8'h00
            reg_file[6698] <= 8'h00
            reg_file[6699] <= 8'h00
            reg_file[6700] <= 8'h00
            reg_file[6701] <= 8'h00
            reg_file[6702] <= 8'h00
            reg_file[6703] <= 8'h00
            reg_file[6704] <= 8'h00
            reg_file[6705] <= 8'h00
            reg_file[6706] <= 8'h00
            reg_file[6707] <= 8'h00
            reg_file[6708] <= 8'h00
            reg_file[6709] <= 8'h00
            reg_file[6710] <= 8'h00
            reg_file[6711] <= 8'h00
            reg_file[6712] <= 8'h00
            reg_file[6713] <= 8'h00
            reg_file[6714] <= 8'h00
            reg_file[6715] <= 8'h00
            reg_file[6716] <= 8'h00
            reg_file[6717] <= 8'h00
            reg_file[6718] <= 8'h00
            reg_file[6719] <= 8'h00
            reg_file[6720] <= 8'h00
            reg_file[6721] <= 8'h00
            reg_file[6722] <= 8'h00
            reg_file[6723] <= 8'h00
            reg_file[6724] <= 8'h00
            reg_file[6725] <= 8'h00
            reg_file[6726] <= 8'h00
            reg_file[6727] <= 8'h00
            reg_file[6728] <= 8'h00
            reg_file[6729] <= 8'h00
            reg_file[6730] <= 8'h00
            reg_file[6731] <= 8'h00
            reg_file[6732] <= 8'h00
            reg_file[6733] <= 8'h00
            reg_file[6734] <= 8'h00
            reg_file[6735] <= 8'h00
            reg_file[6736] <= 8'h00
            reg_file[6737] <= 8'h00
            reg_file[6738] <= 8'h00
            reg_file[6739] <= 8'h00
            reg_file[6740] <= 8'h00
            reg_file[6741] <= 8'h00
            reg_file[6742] <= 8'h00
            reg_file[6743] <= 8'h00
            reg_file[6744] <= 8'h00
            reg_file[6745] <= 8'h00
            reg_file[6746] <= 8'h00
            reg_file[6747] <= 8'h00
            reg_file[6748] <= 8'h00
            reg_file[6749] <= 8'h00
            reg_file[6750] <= 8'h00
            reg_file[6751] <= 8'h00
            reg_file[6752] <= 8'h00
            reg_file[6753] <= 8'h00
            reg_file[6754] <= 8'h00
            reg_file[6755] <= 8'h00
            reg_file[6756] <= 8'h00
            reg_file[6757] <= 8'h00
            reg_file[6758] <= 8'h00
            reg_file[6759] <= 8'h00
            reg_file[6760] <= 8'h00
            reg_file[6761] <= 8'h00
            reg_file[6762] <= 8'h00
            reg_file[6763] <= 8'h00
            reg_file[6764] <= 8'h00
            reg_file[6765] <= 8'h00
            reg_file[6766] <= 8'h00
            reg_file[6767] <= 8'h00
            reg_file[6768] <= 8'h00
            reg_file[6769] <= 8'h00
            reg_file[6770] <= 8'h00
            reg_file[6771] <= 8'h00
            reg_file[6772] <= 8'h00
            reg_file[6773] <= 8'h00
            reg_file[6774] <= 8'h00
            reg_file[6775] <= 8'h00
            reg_file[6776] <= 8'h00
            reg_file[6777] <= 8'h00
            reg_file[6778] <= 8'h00
            reg_file[6779] <= 8'h00
            reg_file[6780] <= 8'h00
            reg_file[6781] <= 8'h00
            reg_file[6782] <= 8'h00
            reg_file[6783] <= 8'h00
            reg_file[6784] <= 8'h00
            reg_file[6785] <= 8'h00
            reg_file[6786] <= 8'h00
            reg_file[6787] <= 8'h00
            reg_file[6788] <= 8'h00
            reg_file[6789] <= 8'h00
            reg_file[6790] <= 8'h00
            reg_file[6791] <= 8'h00
            reg_file[6792] <= 8'h00
            reg_file[6793] <= 8'h00
            reg_file[6794] <= 8'h00
            reg_file[6795] <= 8'h00
            reg_file[6796] <= 8'h00
            reg_file[6797] <= 8'h00
            reg_file[6798] <= 8'h00
            reg_file[6799] <= 8'h00
            reg_file[6800] <= 8'h00
            reg_file[6801] <= 8'h00
            reg_file[6802] <= 8'h00
            reg_file[6803] <= 8'h00
            reg_file[6804] <= 8'h00
            reg_file[6805] <= 8'h00
            reg_file[6806] <= 8'h00
            reg_file[6807] <= 8'h00
            reg_file[6808] <= 8'h00
            reg_file[6809] <= 8'h00
            reg_file[6810] <= 8'h00
            reg_file[6811] <= 8'h00
            reg_file[6812] <= 8'h00
            reg_file[6813] <= 8'h00
            reg_file[6814] <= 8'h00
            reg_file[6815] <= 8'h00
            reg_file[6816] <= 8'h00
            reg_file[6817] <= 8'h00
            reg_file[6818] <= 8'h00
            reg_file[6819] <= 8'h00
            reg_file[6820] <= 8'h00
            reg_file[6821] <= 8'h00
            reg_file[6822] <= 8'h00
            reg_file[6823] <= 8'h00
            reg_file[6824] <= 8'h00
            reg_file[6825] <= 8'h00
            reg_file[6826] <= 8'h00
            reg_file[6827] <= 8'h00
            reg_file[6828] <= 8'h00
            reg_file[6829] <= 8'h00
            reg_file[6830] <= 8'h00
            reg_file[6831] <= 8'h00
            reg_file[6832] <= 8'h00
            reg_file[6833] <= 8'h00
            reg_file[6834] <= 8'h00
            reg_file[6835] <= 8'h00
            reg_file[6836] <= 8'h00
            reg_file[6837] <= 8'h00
            reg_file[6838] <= 8'h00
            reg_file[6839] <= 8'h00
            reg_file[6840] <= 8'h00
            reg_file[6841] <= 8'h00
            reg_file[6842] <= 8'h00
            reg_file[6843] <= 8'h00
            reg_file[6844] <= 8'h00
            reg_file[6845] <= 8'h00
            reg_file[6846] <= 8'h00
            reg_file[6847] <= 8'h00
            reg_file[6848] <= 8'h00
            reg_file[6849] <= 8'h00
            reg_file[6850] <= 8'h00
            reg_file[6851] <= 8'h00
            reg_file[6852] <= 8'h00
            reg_file[6853] <= 8'h00
            reg_file[6854] <= 8'h00
            reg_file[6855] <= 8'h00
            reg_file[6856] <= 8'h00
            reg_file[6857] <= 8'h00
            reg_file[6858] <= 8'h00
            reg_file[6859] <= 8'h00
            reg_file[6860] <= 8'h00
            reg_file[6861] <= 8'h00
            reg_file[6862] <= 8'h00
            reg_file[6863] <= 8'h00
            reg_file[6864] <= 8'h00
            reg_file[6865] <= 8'h00
            reg_file[6866] <= 8'h00
            reg_file[6867] <= 8'h00
            reg_file[6868] <= 8'h00
            reg_file[6869] <= 8'h00
            reg_file[6870] <= 8'h00
            reg_file[6871] <= 8'h00
            reg_file[6872] <= 8'h00
            reg_file[6873] <= 8'h00
            reg_file[6874] <= 8'h00
            reg_file[6875] <= 8'h00
            reg_file[6876] <= 8'h00
            reg_file[6877] <= 8'h00
            reg_file[6878] <= 8'h00
            reg_file[6879] <= 8'h00
            reg_file[6880] <= 8'h00
            reg_file[6881] <= 8'h00
            reg_file[6882] <= 8'h00
            reg_file[6883] <= 8'h00
            reg_file[6884] <= 8'h00
            reg_file[6885] <= 8'h00
            reg_file[6886] <= 8'h00
            reg_file[6887] <= 8'h00
            reg_file[6888] <= 8'h00
            reg_file[6889] <= 8'h00
            reg_file[6890] <= 8'h00
            reg_file[6891] <= 8'h00
            reg_file[6892] <= 8'h00
            reg_file[6893] <= 8'h00
            reg_file[6894] <= 8'h00
            reg_file[6895] <= 8'h00
            reg_file[6896] <= 8'h00
            reg_file[6897] <= 8'h00
            reg_file[6898] <= 8'h00
            reg_file[6899] <= 8'h00
            reg_file[6900] <= 8'h00
            reg_file[6901] <= 8'h00
            reg_file[6902] <= 8'h00
            reg_file[6903] <= 8'h00
            reg_file[6904] <= 8'h00
            reg_file[6905] <= 8'h00
            reg_file[6906] <= 8'h00
            reg_file[6907] <= 8'h00
            reg_file[6908] <= 8'h00
            reg_file[6909] <= 8'h00
            reg_file[6910] <= 8'h00
            reg_file[6911] <= 8'h00
            reg_file[6912] <= 8'h00
            reg_file[6913] <= 8'h00
            reg_file[6914] <= 8'h00
            reg_file[6915] <= 8'h00
            reg_file[6916] <= 8'h00
            reg_file[6917] <= 8'h00
            reg_file[6918] <= 8'h00
            reg_file[6919] <= 8'h00
            reg_file[6920] <= 8'h00
            reg_file[6921] <= 8'h00
            reg_file[6922] <= 8'h00
            reg_file[6923] <= 8'h00
            reg_file[6924] <= 8'h00
            reg_file[6925] <= 8'h00
            reg_file[6926] <= 8'h00
            reg_file[6927] <= 8'h00
            reg_file[6928] <= 8'h00
            reg_file[6929] <= 8'h00
            reg_file[6930] <= 8'h00
            reg_file[6931] <= 8'h00
            reg_file[6932] <= 8'h00
            reg_file[6933] <= 8'h00
            reg_file[6934] <= 8'h00
            reg_file[6935] <= 8'h00
            reg_file[6936] <= 8'h00
            reg_file[6937] <= 8'h00
            reg_file[6938] <= 8'h00
            reg_file[6939] <= 8'h00
            reg_file[6940] <= 8'h00
            reg_file[6941] <= 8'h00
            reg_file[6942] <= 8'h00
            reg_file[6943] <= 8'h00
            reg_file[6944] <= 8'h00
            reg_file[6945] <= 8'h00
            reg_file[6946] <= 8'h00
            reg_file[6947] <= 8'h00
            reg_file[6948] <= 8'h00
            reg_file[6949] <= 8'h00
            reg_file[6950] <= 8'h00
            reg_file[6951] <= 8'h00
            reg_file[6952] <= 8'h00
            reg_file[6953] <= 8'h00
            reg_file[6954] <= 8'h00
            reg_file[6955] <= 8'h00
            reg_file[6956] <= 8'h00
            reg_file[6957] <= 8'h00
            reg_file[6958] <= 8'h00
            reg_file[6959] <= 8'h00
            reg_file[6960] <= 8'h00
            reg_file[6961] <= 8'h00
            reg_file[6962] <= 8'h00
            reg_file[6963] <= 8'h00
            reg_file[6964] <= 8'h00
            reg_file[6965] <= 8'h00
            reg_file[6966] <= 8'h00
            reg_file[6967] <= 8'h00
            reg_file[6968] <= 8'h00
            reg_file[6969] <= 8'h00
            reg_file[6970] <= 8'h00
            reg_file[6971] <= 8'h00
            reg_file[6972] <= 8'h00
            reg_file[6973] <= 8'h00
            reg_file[6974] <= 8'h00
            reg_file[6975] <= 8'h00
            reg_file[6976] <= 8'h00
            reg_file[6977] <= 8'h00
            reg_file[6978] <= 8'h00
            reg_file[6979] <= 8'h00
            reg_file[6980] <= 8'h00
            reg_file[6981] <= 8'h00
            reg_file[6982] <= 8'h00
            reg_file[6983] <= 8'h00
            reg_file[6984] <= 8'h00
            reg_file[6985] <= 8'h00
            reg_file[6986] <= 8'h00
            reg_file[6987] <= 8'h00
            reg_file[6988] <= 8'h00
            reg_file[6989] <= 8'h00
            reg_file[6990] <= 8'h00
            reg_file[6991] <= 8'h00
            reg_file[6992] <= 8'h00
            reg_file[6993] <= 8'h00
            reg_file[6994] <= 8'h00
            reg_file[6995] <= 8'h00
            reg_file[6996] <= 8'h00
            reg_file[6997] <= 8'h00
            reg_file[6998] <= 8'h00
            reg_file[6999] <= 8'h00
            reg_file[7000] <= 8'h00
            reg_file[7001] <= 8'h00
            reg_file[7002] <= 8'h00
            reg_file[7003] <= 8'h00
            reg_file[7004] <= 8'h00
            reg_file[7005] <= 8'h00
            reg_file[7006] <= 8'h00
            reg_file[7007] <= 8'h00
            reg_file[7008] <= 8'h00
            reg_file[7009] <= 8'h00
            reg_file[7010] <= 8'h00
            reg_file[7011] <= 8'h00
            reg_file[7012] <= 8'h00
            reg_file[7013] <= 8'h00
            reg_file[7014] <= 8'h00
            reg_file[7015] <= 8'h00
            reg_file[7016] <= 8'h00
            reg_file[7017] <= 8'h00
            reg_file[7018] <= 8'h00
            reg_file[7019] <= 8'h00
            reg_file[7020] <= 8'h00
            reg_file[7021] <= 8'h00
            reg_file[7022] <= 8'h00
            reg_file[7023] <= 8'h00
            reg_file[7024] <= 8'h00
            reg_file[7025] <= 8'h00
            reg_file[7026] <= 8'h00
            reg_file[7027] <= 8'h00
            reg_file[7028] <= 8'h00
            reg_file[7029] <= 8'h00
            reg_file[7030] <= 8'h00
            reg_file[7031] <= 8'h00
            reg_file[7032] <= 8'h00
            reg_file[7033] <= 8'h00
            reg_file[7034] <= 8'h00
            reg_file[7035] <= 8'h00
            reg_file[7036] <= 8'h00
            reg_file[7037] <= 8'h00
            reg_file[7038] <= 8'h00
            reg_file[7039] <= 8'h00
            reg_file[7040] <= 8'h00
            reg_file[7041] <= 8'h00
            reg_file[7042] <= 8'h00
            reg_file[7043] <= 8'h00
            reg_file[7044] <= 8'h00
            reg_file[7045] <= 8'h00
            reg_file[7046] <= 8'h00
            reg_file[7047] <= 8'h00
            reg_file[7048] <= 8'h00
            reg_file[7049] <= 8'h00
            reg_file[7050] <= 8'h00
            reg_file[7051] <= 8'h00
            reg_file[7052] <= 8'h00
            reg_file[7053] <= 8'h00
            reg_file[7054] <= 8'h00
            reg_file[7055] <= 8'h00
            reg_file[7056] <= 8'h00
            reg_file[7057] <= 8'h00
            reg_file[7058] <= 8'h00
            reg_file[7059] <= 8'h00
            reg_file[7060] <= 8'h00
            reg_file[7061] <= 8'h00
            reg_file[7062] <= 8'h00
            reg_file[7063] <= 8'h00
            reg_file[7064] <= 8'h00
            reg_file[7065] <= 8'h00
            reg_file[7066] <= 8'h00
            reg_file[7067] <= 8'h00
            reg_file[7068] <= 8'h00
            reg_file[7069] <= 8'h00
            reg_file[7070] <= 8'h00
            reg_file[7071] <= 8'h00
            reg_file[7072] <= 8'h00
            reg_file[7073] <= 8'h00
            reg_file[7074] <= 8'h00
            reg_file[7075] <= 8'h00
            reg_file[7076] <= 8'h00
            reg_file[7077] <= 8'h00
            reg_file[7078] <= 8'h00
            reg_file[7079] <= 8'h00
            reg_file[7080] <= 8'h00
            reg_file[7081] <= 8'h00
            reg_file[7082] <= 8'h00
            reg_file[7083] <= 8'h00
            reg_file[7084] <= 8'h00
            reg_file[7085] <= 8'h00
            reg_file[7086] <= 8'h00
            reg_file[7087] <= 8'h00
            reg_file[7088] <= 8'h00
            reg_file[7089] <= 8'h00
            reg_file[7090] <= 8'h00
            reg_file[7091] <= 8'h00
            reg_file[7092] <= 8'h00
            reg_file[7093] <= 8'h00
            reg_file[7094] <= 8'h00
            reg_file[7095] <= 8'h00
            reg_file[7096] <= 8'h00
            reg_file[7097] <= 8'h00
            reg_file[7098] <= 8'h00
            reg_file[7099] <= 8'h00
            reg_file[7100] <= 8'h00
            reg_file[7101] <= 8'h00
            reg_file[7102] <= 8'h00
            reg_file[7103] <= 8'h00
            reg_file[7104] <= 8'h00
            reg_file[7105] <= 8'h00
            reg_file[7106] <= 8'h00
            reg_file[7107] <= 8'h00
            reg_file[7108] <= 8'h00
            reg_file[7109] <= 8'h00
            reg_file[7110] <= 8'h00
            reg_file[7111] <= 8'h00
            reg_file[7112] <= 8'h00
            reg_file[7113] <= 8'h00
            reg_file[7114] <= 8'h00
            reg_file[7115] <= 8'h00
            reg_file[7116] <= 8'h00
            reg_file[7117] <= 8'h00
            reg_file[7118] <= 8'h00
            reg_file[7119] <= 8'h00
            reg_file[7120] <= 8'h00
            reg_file[7121] <= 8'h00
            reg_file[7122] <= 8'h00
            reg_file[7123] <= 8'h00
            reg_file[7124] <= 8'h00
            reg_file[7125] <= 8'h00
            reg_file[7126] <= 8'h00
            reg_file[7127] <= 8'h00
            reg_file[7128] <= 8'h00
            reg_file[7129] <= 8'h00
            reg_file[7130] <= 8'h00
            reg_file[7131] <= 8'h00
            reg_file[7132] <= 8'h00
            reg_file[7133] <= 8'h00
            reg_file[7134] <= 8'h00
            reg_file[7135] <= 8'h00
            reg_file[7136] <= 8'h00
            reg_file[7137] <= 8'h00
            reg_file[7138] <= 8'h00
            reg_file[7139] <= 8'h00
            reg_file[7140] <= 8'h00
            reg_file[7141] <= 8'h00
            reg_file[7142] <= 8'h00
            reg_file[7143] <= 8'h00
            reg_file[7144] <= 8'h00
            reg_file[7145] <= 8'h00
            reg_file[7146] <= 8'h00
            reg_file[7147] <= 8'h00
            reg_file[7148] <= 8'h00
            reg_file[7149] <= 8'h00
            reg_file[7150] <= 8'h00
            reg_file[7151] <= 8'h00
            reg_file[7152] <= 8'h00
            reg_file[7153] <= 8'h00
            reg_file[7154] <= 8'h00
            reg_file[7155] <= 8'h00
            reg_file[7156] <= 8'h00
            reg_file[7157] <= 8'h00
            reg_file[7158] <= 8'h00
            reg_file[7159] <= 8'h00
            reg_file[7160] <= 8'h00
            reg_file[7161] <= 8'h00
            reg_file[7162] <= 8'h00
            reg_file[7163] <= 8'h00
            reg_file[7164] <= 8'h00
            reg_file[7165] <= 8'h00
            reg_file[7166] <= 8'h00
            reg_file[7167] <= 8'h00
            reg_file[7168] <= 8'h00
            reg_file[7169] <= 8'h00
            reg_file[7170] <= 8'h00
            reg_file[7171] <= 8'h00
            reg_file[7172] <= 8'h00
            reg_file[7173] <= 8'h00
            reg_file[7174] <= 8'h00
            reg_file[7175] <= 8'h00
            reg_file[7176] <= 8'h00
            reg_file[7177] <= 8'h00
            reg_file[7178] <= 8'h00
            reg_file[7179] <= 8'h00
            reg_file[7180] <= 8'h00
            reg_file[7181] <= 8'h00
            reg_file[7182] <= 8'h00
            reg_file[7183] <= 8'h00
            reg_file[7184] <= 8'h00
            reg_file[7185] <= 8'h00
            reg_file[7186] <= 8'h00
            reg_file[7187] <= 8'h00
            reg_file[7188] <= 8'h00
            reg_file[7189] <= 8'h00
            reg_file[7190] <= 8'h00
            reg_file[7191] <= 8'h00
            reg_file[7192] <= 8'h00
            reg_file[7193] <= 8'h00
            reg_file[7194] <= 8'h00
            reg_file[7195] <= 8'h00
            reg_file[7196] <= 8'h00
            reg_file[7197] <= 8'h00
            reg_file[7198] <= 8'h00
            reg_file[7199] <= 8'h00
            reg_file[7200] <= 8'h00
            reg_file[7201] <= 8'h00
            reg_file[7202] <= 8'h00
            reg_file[7203] <= 8'h00
            reg_file[7204] <= 8'h00
            reg_file[7205] <= 8'h00
            reg_file[7206] <= 8'h00
            reg_file[7207] <= 8'h00
            reg_file[7208] <= 8'h00
            reg_file[7209] <= 8'h00
            reg_file[7210] <= 8'h00
            reg_file[7211] <= 8'h00
            reg_file[7212] <= 8'h00
            reg_file[7213] <= 8'h00
            reg_file[7214] <= 8'h00
            reg_file[7215] <= 8'h00
            reg_file[7216] <= 8'h00
            reg_file[7217] <= 8'h00
            reg_file[7218] <= 8'h00
            reg_file[7219] <= 8'h00
            reg_file[7220] <= 8'h00
            reg_file[7221] <= 8'h00
            reg_file[7222] <= 8'h00
            reg_file[7223] <= 8'h00
            reg_file[7224] <= 8'h00
            reg_file[7225] <= 8'h00
            reg_file[7226] <= 8'h00
            reg_file[7227] <= 8'h00
            reg_file[7228] <= 8'h00
            reg_file[7229] <= 8'h00
            reg_file[7230] <= 8'h00
            reg_file[7231] <= 8'h00
            reg_file[7232] <= 8'h00
            reg_file[7233] <= 8'h00
            reg_file[7234] <= 8'h00
            reg_file[7235] <= 8'h00
            reg_file[7236] <= 8'h00
            reg_file[7237] <= 8'h00
            reg_file[7238] <= 8'h00
            reg_file[7239] <= 8'h00
            reg_file[7240] <= 8'h00
            reg_file[7241] <= 8'h00
            reg_file[7242] <= 8'h00
            reg_file[7243] <= 8'h00
            reg_file[7244] <= 8'h00
            reg_file[7245] <= 8'h00
            reg_file[7246] <= 8'h00
            reg_file[7247] <= 8'h00
            reg_file[7248] <= 8'h00
            reg_file[7249] <= 8'h00
            reg_file[7250] <= 8'h00
            reg_file[7251] <= 8'h00
            reg_file[7252] <= 8'h00
            reg_file[7253] <= 8'h00
            reg_file[7254] <= 8'h00
            reg_file[7255] <= 8'h00
            reg_file[7256] <= 8'h00
            reg_file[7257] <= 8'h00
            reg_file[7258] <= 8'h00
            reg_file[7259] <= 8'h00
            reg_file[7260] <= 8'h00
            reg_file[7261] <= 8'h00
            reg_file[7262] <= 8'h00
            reg_file[7263] <= 8'h00
            reg_file[7264] <= 8'h00
            reg_file[7265] <= 8'h00
            reg_file[7266] <= 8'h00
            reg_file[7267] <= 8'h00
            reg_file[7268] <= 8'h00
            reg_file[7269] <= 8'h00
            reg_file[7270] <= 8'h00
            reg_file[7271] <= 8'h00
            reg_file[7272] <= 8'h00
            reg_file[7273] <= 8'h00
            reg_file[7274] <= 8'h00
            reg_file[7275] <= 8'h00
            reg_file[7276] <= 8'h00
            reg_file[7277] <= 8'h00
            reg_file[7278] <= 8'h00
            reg_file[7279] <= 8'h00
            reg_file[7280] <= 8'h00
            reg_file[7281] <= 8'h00
            reg_file[7282] <= 8'h00
            reg_file[7283] <= 8'h00
            reg_file[7284] <= 8'h00
            reg_file[7285] <= 8'h00
            reg_file[7286] <= 8'h00
            reg_file[7287] <= 8'h00
            reg_file[7288] <= 8'h00
            reg_file[7289] <= 8'h00
            reg_file[7290] <= 8'h00
            reg_file[7291] <= 8'h00
            reg_file[7292] <= 8'h00
            reg_file[7293] <= 8'h00
            reg_file[7294] <= 8'h00
            reg_file[7295] <= 8'h00
            reg_file[7296] <= 8'h00
            reg_file[7297] <= 8'h00
            reg_file[7298] <= 8'h00
            reg_file[7299] <= 8'h00
            reg_file[7300] <= 8'h00
            reg_file[7301] <= 8'h00
            reg_file[7302] <= 8'h00
            reg_file[7303] <= 8'h00
            reg_file[7304] <= 8'h00
            reg_file[7305] <= 8'h00
            reg_file[7306] <= 8'h00
            reg_file[7307] <= 8'h00
            reg_file[7308] <= 8'h00
            reg_file[7309] <= 8'h00
            reg_file[7310] <= 8'h00
            reg_file[7311] <= 8'h00
            reg_file[7312] <= 8'h00
            reg_file[7313] <= 8'h00
            reg_file[7314] <= 8'h00
            reg_file[7315] <= 8'h00
            reg_file[7316] <= 8'h00
            reg_file[7317] <= 8'h00
            reg_file[7318] <= 8'h00
            reg_file[7319] <= 8'h00
            reg_file[7320] <= 8'h00
            reg_file[7321] <= 8'h00
            reg_file[7322] <= 8'h00
            reg_file[7323] <= 8'h00
            reg_file[7324] <= 8'h00
            reg_file[7325] <= 8'h00
            reg_file[7326] <= 8'h00
            reg_file[7327] <= 8'h00
            reg_file[7328] <= 8'h00
            reg_file[7329] <= 8'h00
            reg_file[7330] <= 8'h00
            reg_file[7331] <= 8'h00
            reg_file[7332] <= 8'h00
            reg_file[7333] <= 8'h00
            reg_file[7334] <= 8'h00
            reg_file[7335] <= 8'h00
            reg_file[7336] <= 8'h00
            reg_file[7337] <= 8'h00
            reg_file[7338] <= 8'h00
            reg_file[7339] <= 8'h00
            reg_file[7340] <= 8'h00
            reg_file[7341] <= 8'h00
            reg_file[7342] <= 8'h00
            reg_file[7343] <= 8'h00
            reg_file[7344] <= 8'h00
            reg_file[7345] <= 8'h00
            reg_file[7346] <= 8'h00
            reg_file[7347] <= 8'h00
            reg_file[7348] <= 8'h00
            reg_file[7349] <= 8'h00
            reg_file[7350] <= 8'h00
            reg_file[7351] <= 8'h00
            reg_file[7352] <= 8'h00
            reg_file[7353] <= 8'h00
            reg_file[7354] <= 8'h00
            reg_file[7355] <= 8'h00
            reg_file[7356] <= 8'h00
            reg_file[7357] <= 8'h00
            reg_file[7358] <= 8'h00
            reg_file[7359] <= 8'h00
            reg_file[7360] <= 8'h00
            reg_file[7361] <= 8'h00
            reg_file[7362] <= 8'h00
            reg_file[7363] <= 8'h00
            reg_file[7364] <= 8'h00
            reg_file[7365] <= 8'h00
            reg_file[7366] <= 8'h00
            reg_file[7367] <= 8'h00
            reg_file[7368] <= 8'h00
            reg_file[7369] <= 8'h00
            reg_file[7370] <= 8'h00
            reg_file[7371] <= 8'h00
            reg_file[7372] <= 8'h00
            reg_file[7373] <= 8'h00
            reg_file[7374] <= 8'h00
            reg_file[7375] <= 8'h00
            reg_file[7376] <= 8'h00
            reg_file[7377] <= 8'h00
            reg_file[7378] <= 8'h00
            reg_file[7379] <= 8'h00
            reg_file[7380] <= 8'h00
            reg_file[7381] <= 8'h00
            reg_file[7382] <= 8'h00
            reg_file[7383] <= 8'h00
            reg_file[7384] <= 8'h00
            reg_file[7385] <= 8'h00
            reg_file[7386] <= 8'h00
            reg_file[7387] <= 8'h00
            reg_file[7388] <= 8'h00
            reg_file[7389] <= 8'h00
            reg_file[7390] <= 8'h00
            reg_file[7391] <= 8'h00
            reg_file[7392] <= 8'h00
            reg_file[7393] <= 8'h00
            reg_file[7394] <= 8'h00
            reg_file[7395] <= 8'h00
            reg_file[7396] <= 8'h00
            reg_file[7397] <= 8'h00
            reg_file[7398] <= 8'h00
            reg_file[7399] <= 8'h00
            reg_file[7400] <= 8'h00
            reg_file[7401] <= 8'h00
            reg_file[7402] <= 8'h00
            reg_file[7403] <= 8'h00
            reg_file[7404] <= 8'h00
            reg_file[7405] <= 8'h00
            reg_file[7406] <= 8'h00
            reg_file[7407] <= 8'h00
            reg_file[7408] <= 8'h00
            reg_file[7409] <= 8'h00
            reg_file[7410] <= 8'h00
            reg_file[7411] <= 8'h00
            reg_file[7412] <= 8'h00
            reg_file[7413] <= 8'h00
            reg_file[7414] <= 8'h00
            reg_file[7415] <= 8'h00
            reg_file[7416] <= 8'h00
            reg_file[7417] <= 8'h00
            reg_file[7418] <= 8'h00
            reg_file[7419] <= 8'h00
            reg_file[7420] <= 8'h00
            reg_file[7421] <= 8'h00
            reg_file[7422] <= 8'h00
            reg_file[7423] <= 8'h00
            reg_file[7424] <= 8'h00
            reg_file[7425] <= 8'h00
            reg_file[7426] <= 8'h00
            reg_file[7427] <= 8'h00
            reg_file[7428] <= 8'h00
            reg_file[7429] <= 8'h00
            reg_file[7430] <= 8'h00
            reg_file[7431] <= 8'h00
            reg_file[7432] <= 8'h00
            reg_file[7433] <= 8'h00
            reg_file[7434] <= 8'h00
            reg_file[7435] <= 8'h00
            reg_file[7436] <= 8'h00
            reg_file[7437] <= 8'h00
            reg_file[7438] <= 8'h00
            reg_file[7439] <= 8'h00
            reg_file[7440] <= 8'h00
            reg_file[7441] <= 8'h00
            reg_file[7442] <= 8'h00
            reg_file[7443] <= 8'h00
            reg_file[7444] <= 8'h00
            reg_file[7445] <= 8'h00
            reg_file[7446] <= 8'h00
            reg_file[7447] <= 8'h00
            reg_file[7448] <= 8'h00
            reg_file[7449] <= 8'h00
            reg_file[7450] <= 8'h00
            reg_file[7451] <= 8'h00
            reg_file[7452] <= 8'h00
            reg_file[7453] <= 8'h00
            reg_file[7454] <= 8'h00
            reg_file[7455] <= 8'h00
            reg_file[7456] <= 8'h00
            reg_file[7457] <= 8'h00
            reg_file[7458] <= 8'h00
            reg_file[7459] <= 8'h00
            reg_file[7460] <= 8'h00
            reg_file[7461] <= 8'h00
            reg_file[7462] <= 8'h00
            reg_file[7463] <= 8'h00
            reg_file[7464] <= 8'h00
            reg_file[7465] <= 8'h00
            reg_file[7466] <= 8'h00
            reg_file[7467] <= 8'h00
            reg_file[7468] <= 8'h00
            reg_file[7469] <= 8'h00
            reg_file[7470] <= 8'h00
            reg_file[7471] <= 8'h00
            reg_file[7472] <= 8'h00
            reg_file[7473] <= 8'h00
            reg_file[7474] <= 8'h00
            reg_file[7475] <= 8'h00
            reg_file[7476] <= 8'h00
            reg_file[7477] <= 8'h00
            reg_file[7478] <= 8'h00
            reg_file[7479] <= 8'h00
            reg_file[7480] <= 8'h00
            reg_file[7481] <= 8'h00
            reg_file[7482] <= 8'h00
            reg_file[7483] <= 8'h00
            reg_file[7484] <= 8'h00
            reg_file[7485] <= 8'h00
            reg_file[7486] <= 8'h00
            reg_file[7487] <= 8'h00
            reg_file[7488] <= 8'h00
            reg_file[7489] <= 8'h00
            reg_file[7490] <= 8'h00
            reg_file[7491] <= 8'h00
            reg_file[7492] <= 8'h00
            reg_file[7493] <= 8'h00
            reg_file[7494] <= 8'h00
            reg_file[7495] <= 8'h00
            reg_file[7496] <= 8'h00
            reg_file[7497] <= 8'h00
            reg_file[7498] <= 8'h00
            reg_file[7499] <= 8'h00
            reg_file[7500] <= 8'h00
            reg_file[7501] <= 8'h00
            reg_file[7502] <= 8'h00
            reg_file[7503] <= 8'h00
            reg_file[7504] <= 8'h00
            reg_file[7505] <= 8'h00
            reg_file[7506] <= 8'h00
            reg_file[7507] <= 8'h00
            reg_file[7508] <= 8'h00
            reg_file[7509] <= 8'h00
            reg_file[7510] <= 8'h00
            reg_file[7511] <= 8'h00
            reg_file[7512] <= 8'h00
            reg_file[7513] <= 8'h00
            reg_file[7514] <= 8'h00
            reg_file[7515] <= 8'h00
            reg_file[7516] <= 8'h00
            reg_file[7517] <= 8'h00
            reg_file[7518] <= 8'h00
            reg_file[7519] <= 8'h00
            reg_file[7520] <= 8'h00
            reg_file[7521] <= 8'h00
            reg_file[7522] <= 8'h00
            reg_file[7523] <= 8'h00
            reg_file[7524] <= 8'h00
            reg_file[7525] <= 8'h00
            reg_file[7526] <= 8'h00
            reg_file[7527] <= 8'h00
            reg_file[7528] <= 8'h00
            reg_file[7529] <= 8'h00
            reg_file[7530] <= 8'h00
            reg_file[7531] <= 8'h00
            reg_file[7532] <= 8'h00
            reg_file[7533] <= 8'h00
            reg_file[7534] <= 8'h00
            reg_file[7535] <= 8'h00
            reg_file[7536] <= 8'h00
            reg_file[7537] <= 8'h00
            reg_file[7538] <= 8'h00
            reg_file[7539] <= 8'h00
            reg_file[7540] <= 8'h00
            reg_file[7541] <= 8'h00
            reg_file[7542] <= 8'h00
            reg_file[7543] <= 8'h00
            reg_file[7544] <= 8'h00
            reg_file[7545] <= 8'h00
            reg_file[7546] <= 8'h00
            reg_file[7547] <= 8'h00
            reg_file[7548] <= 8'h00
            reg_file[7549] <= 8'h00
            reg_file[7550] <= 8'h00
            reg_file[7551] <= 8'h00
            reg_file[7552] <= 8'h00
            reg_file[7553] <= 8'h00
            reg_file[7554] <= 8'h00
            reg_file[7555] <= 8'h00
            reg_file[7556] <= 8'h00
            reg_file[7557] <= 8'h00
            reg_file[7558] <= 8'h00
            reg_file[7559] <= 8'h00
            reg_file[7560] <= 8'h00
            reg_file[7561] <= 8'h00
            reg_file[7562] <= 8'h00
            reg_file[7563] <= 8'h00
            reg_file[7564] <= 8'h00
            reg_file[7565] <= 8'h00
            reg_file[7566] <= 8'h00
            reg_file[7567] <= 8'h00
            reg_file[7568] <= 8'h00
            reg_file[7569] <= 8'h00
            reg_file[7570] <= 8'h00
            reg_file[7571] <= 8'h00
            reg_file[7572] <= 8'h00
            reg_file[7573] <= 8'h00
            reg_file[7574] <= 8'h00
            reg_file[7575] <= 8'h00
            reg_file[7576] <= 8'h00
            reg_file[7577] <= 8'h00
            reg_file[7578] <= 8'h00
            reg_file[7579] <= 8'h00
            reg_file[7580] <= 8'h00
            reg_file[7581] <= 8'h00
            reg_file[7582] <= 8'h00
            reg_file[7583] <= 8'h00
            reg_file[7584] <= 8'h00
            reg_file[7585] <= 8'h00
            reg_file[7586] <= 8'h00
            reg_file[7587] <= 8'h00
            reg_file[7588] <= 8'h00
            reg_file[7589] <= 8'h00
            reg_file[7590] <= 8'h00
            reg_file[7591] <= 8'h00
            reg_file[7592] <= 8'h00
            reg_file[7593] <= 8'h00
            reg_file[7594] <= 8'h00
            reg_file[7595] <= 8'h00
            reg_file[7596] <= 8'h00
            reg_file[7597] <= 8'h00
            reg_file[7598] <= 8'h00
            reg_file[7599] <= 8'h00
            reg_file[7600] <= 8'h00
            reg_file[7601] <= 8'h00
            reg_file[7602] <= 8'h00
            reg_file[7603] <= 8'h00
            reg_file[7604] <= 8'h00
            reg_file[7605] <= 8'h00
            reg_file[7606] <= 8'h00
            reg_file[7607] <= 8'h00
            reg_file[7608] <= 8'h00
            reg_file[7609] <= 8'h00
            reg_file[7610] <= 8'h00
            reg_file[7611] <= 8'h00
            reg_file[7612] <= 8'h00
            reg_file[7613] <= 8'h00
            reg_file[7614] <= 8'h00
            reg_file[7615] <= 8'h00
            reg_file[7616] <= 8'h00
            reg_file[7617] <= 8'h00
            reg_file[7618] <= 8'h00
            reg_file[7619] <= 8'h00
            reg_file[7620] <= 8'h00
            reg_file[7621] <= 8'h00
            reg_file[7622] <= 8'h00
            reg_file[7623] <= 8'h00
            reg_file[7624] <= 8'h00
            reg_file[7625] <= 8'h00
            reg_file[7626] <= 8'h00
            reg_file[7627] <= 8'h00
            reg_file[7628] <= 8'h00
            reg_file[7629] <= 8'h00
            reg_file[7630] <= 8'h00
            reg_file[7631] <= 8'h00
            reg_file[7632] <= 8'h00
            reg_file[7633] <= 8'h00
            reg_file[7634] <= 8'h00
            reg_file[7635] <= 8'h00
            reg_file[7636] <= 8'h00
            reg_file[7637] <= 8'h00
            reg_file[7638] <= 8'h00
            reg_file[7639] <= 8'h00
            reg_file[7640] <= 8'h00
            reg_file[7641] <= 8'h00
            reg_file[7642] <= 8'h00
            reg_file[7643] <= 8'h00
            reg_file[7644] <= 8'h00
            reg_file[7645] <= 8'h00
            reg_file[7646] <= 8'h00
            reg_file[7647] <= 8'h00
            reg_file[7648] <= 8'h00
            reg_file[7649] <= 8'h00
            reg_file[7650] <= 8'h00
            reg_file[7651] <= 8'h00
            reg_file[7652] <= 8'h00
            reg_file[7653] <= 8'h00
            reg_file[7654] <= 8'h00
            reg_file[7655] <= 8'h00
            reg_file[7656] <= 8'h00
            reg_file[7657] <= 8'h00
            reg_file[7658] <= 8'h00
            reg_file[7659] <= 8'h00
            reg_file[7660] <= 8'h00
            reg_file[7661] <= 8'h00
            reg_file[7662] <= 8'h00
            reg_file[7663] <= 8'h00
            reg_file[7664] <= 8'h00
            reg_file[7665] <= 8'h00
            reg_file[7666] <= 8'h00
            reg_file[7667] <= 8'h00
            reg_file[7668] <= 8'h00
            reg_file[7669] <= 8'h00
            reg_file[7670] <= 8'h00
            reg_file[7671] <= 8'h00
            reg_file[7672] <= 8'h00
            reg_file[7673] <= 8'h00
            reg_file[7674] <= 8'h00
            reg_file[7675] <= 8'h00
            reg_file[7676] <= 8'h00
            reg_file[7677] <= 8'h00
            reg_file[7678] <= 8'h00
            reg_file[7679] <= 8'h00
            reg_file[7680] <= 8'h00
            reg_file[7681] <= 8'h00
            reg_file[7682] <= 8'h00
            reg_file[7683] <= 8'h00
            reg_file[7684] <= 8'h00
            reg_file[7685] <= 8'h00
            reg_file[7686] <= 8'h00
            reg_file[7687] <= 8'h00
            reg_file[7688] <= 8'h00
            reg_file[7689] <= 8'h00
            reg_file[7690] <= 8'h00
            reg_file[7691] <= 8'h00
            reg_file[7692] <= 8'h00
            reg_file[7693] <= 8'h00
            reg_file[7694] <= 8'h00
            reg_file[7695] <= 8'h00
            reg_file[7696] <= 8'h00
            reg_file[7697] <= 8'h00
            reg_file[7698] <= 8'h00
            reg_file[7699] <= 8'h00
            reg_file[7700] <= 8'h00
            reg_file[7701] <= 8'h00
            reg_file[7702] <= 8'h00
            reg_file[7703] <= 8'h00
            reg_file[7704] <= 8'h00
            reg_file[7705] <= 8'h00
            reg_file[7706] <= 8'h00
            reg_file[7707] <= 8'h00
            reg_file[7708] <= 8'h00
            reg_file[7709] <= 8'h00
            reg_file[7710] <= 8'h00
            reg_file[7711] <= 8'h00
            reg_file[7712] <= 8'h00
            reg_file[7713] <= 8'h00
            reg_file[7714] <= 8'h00
            reg_file[7715] <= 8'h00
            reg_file[7716] <= 8'h00
            reg_file[7717] <= 8'h00
            reg_file[7718] <= 8'h00
            reg_file[7719] <= 8'h00
            reg_file[7720] <= 8'h00
            reg_file[7721] <= 8'h00
            reg_file[7722] <= 8'h00
            reg_file[7723] <= 8'h00
            reg_file[7724] <= 8'h00
            reg_file[7725] <= 8'h00
            reg_file[7726] <= 8'h00
            reg_file[7727] <= 8'h00
            reg_file[7728] <= 8'h00
            reg_file[7729] <= 8'h00
            reg_file[7730] <= 8'h00
            reg_file[7731] <= 8'h00
            reg_file[7732] <= 8'h00
            reg_file[7733] <= 8'h00
            reg_file[7734] <= 8'h00
            reg_file[7735] <= 8'h00
            reg_file[7736] <= 8'h00
            reg_file[7737] <= 8'h00
            reg_file[7738] <= 8'h00
            reg_file[7739] <= 8'h00
            reg_file[7740] <= 8'h00
            reg_file[7741] <= 8'h00
            reg_file[7742] <= 8'h00
            reg_file[7743] <= 8'h00
            reg_file[7744] <= 8'h00
            reg_file[7745] <= 8'h00
            reg_file[7746] <= 8'h00
            reg_file[7747] <= 8'h00
            reg_file[7748] <= 8'h00
            reg_file[7749] <= 8'h00
            reg_file[7750] <= 8'h00
            reg_file[7751] <= 8'h00
            reg_file[7752] <= 8'h00
            reg_file[7753] <= 8'h00
            reg_file[7754] <= 8'h00
            reg_file[7755] <= 8'h00
            reg_file[7756] <= 8'h00
            reg_file[7757] <= 8'h00
            reg_file[7758] <= 8'h00
            reg_file[7759] <= 8'h00
            reg_file[7760] <= 8'h00
            reg_file[7761] <= 8'h00
            reg_file[7762] <= 8'h00
            reg_file[7763] <= 8'h00
            reg_file[7764] <= 8'h00
            reg_file[7765] <= 8'h00
            reg_file[7766] <= 8'h00
            reg_file[7767] <= 8'h00
            reg_file[7768] <= 8'h00
            reg_file[7769] <= 8'h00
            reg_file[7770] <= 8'h00
            reg_file[7771] <= 8'h00
            reg_file[7772] <= 8'h00
            reg_file[7773] <= 8'h00
            reg_file[7774] <= 8'h00
            reg_file[7775] <= 8'h00
            reg_file[7776] <= 8'h00
            reg_file[7777] <= 8'h00
            reg_file[7778] <= 8'h00
            reg_file[7779] <= 8'h00
            reg_file[7780] <= 8'h00
            reg_file[7781] <= 8'h00
            reg_file[7782] <= 8'h00
            reg_file[7783] <= 8'h00
            reg_file[7784] <= 8'h00
            reg_file[7785] <= 8'h00
            reg_file[7786] <= 8'h00
            reg_file[7787] <= 8'h00
            reg_file[7788] <= 8'h00
            reg_file[7789] <= 8'h00
            reg_file[7790] <= 8'h00
            reg_file[7791] <= 8'h00
            reg_file[7792] <= 8'h00
            reg_file[7793] <= 8'h00
            reg_file[7794] <= 8'h00
            reg_file[7795] <= 8'h00
            reg_file[7796] <= 8'h00
            reg_file[7797] <= 8'h00
            reg_file[7798] <= 8'h00
            reg_file[7799] <= 8'h00
            reg_file[7800] <= 8'h00
            reg_file[7801] <= 8'h00
            reg_file[7802] <= 8'h00
            reg_file[7803] <= 8'h00
            reg_file[7804] <= 8'h00
            reg_file[7805] <= 8'h00
            reg_file[7806] <= 8'h00
            reg_file[7807] <= 8'h00
            reg_file[7808] <= 8'h00
            reg_file[7809] <= 8'h00
            reg_file[7810] <= 8'h00
            reg_file[7811] <= 8'h00
            reg_file[7812] <= 8'h00
            reg_file[7813] <= 8'h00
            reg_file[7814] <= 8'h00
            reg_file[7815] <= 8'h00
            reg_file[7816] <= 8'h00
            reg_file[7817] <= 8'h00
            reg_file[7818] <= 8'h00
            reg_file[7819] <= 8'h00
            reg_file[7820] <= 8'h00
            reg_file[7821] <= 8'h00
            reg_file[7822] <= 8'h00
            reg_file[7823] <= 8'h00
            reg_file[7824] <= 8'h00
            reg_file[7825] <= 8'h00
            reg_file[7826] <= 8'h00
            reg_file[7827] <= 8'h00
            reg_file[7828] <= 8'h00
            reg_file[7829] <= 8'h00
            reg_file[7830] <= 8'h00
            reg_file[7831] <= 8'h00
            reg_file[7832] <= 8'h00
            reg_file[7833] <= 8'h00
            reg_file[7834] <= 8'h00
            reg_file[7835] <= 8'h00
            reg_file[7836] <= 8'h00
            reg_file[7837] <= 8'h00
            reg_file[7838] <= 8'h00
            reg_file[7839] <= 8'h00
            reg_file[7840] <= 8'h00
            reg_file[7841] <= 8'h00
            reg_file[7842] <= 8'h00
            reg_file[7843] <= 8'h00
            reg_file[7844] <= 8'h00
            reg_file[7845] <= 8'h00
            reg_file[7846] <= 8'h00
            reg_file[7847] <= 8'h00
            reg_file[7848] <= 8'h00
            reg_file[7849] <= 8'h00
            reg_file[7850] <= 8'h00
            reg_file[7851] <= 8'h00
            reg_file[7852] <= 8'h00
            reg_file[7853] <= 8'h00
            reg_file[7854] <= 8'h00
            reg_file[7855] <= 8'h00
            reg_file[7856] <= 8'h00
            reg_file[7857] <= 8'h00
            reg_file[7858] <= 8'h00
            reg_file[7859] <= 8'h00
            reg_file[7860] <= 8'h00
            reg_file[7861] <= 8'h00
            reg_file[7862] <= 8'h00
            reg_file[7863] <= 8'h00
            reg_file[7864] <= 8'h00
            reg_file[7865] <= 8'h00
            reg_file[7866] <= 8'h00
            reg_file[7867] <= 8'h00
            reg_file[7868] <= 8'h00
            reg_file[7869] <= 8'h00
            reg_file[7870] <= 8'h00
            reg_file[7871] <= 8'h00
            reg_file[7872] <= 8'h00
            reg_file[7873] <= 8'h00
            reg_file[7874] <= 8'h00
            reg_file[7875] <= 8'h00
            reg_file[7876] <= 8'h00
            reg_file[7877] <= 8'h00
            reg_file[7878] <= 8'h00
            reg_file[7879] <= 8'h00
            reg_file[7880] <= 8'h00
            reg_file[7881] <= 8'h00
            reg_file[7882] <= 8'h00
            reg_file[7883] <= 8'h00
            reg_file[7884] <= 8'h00
            reg_file[7885] <= 8'h00
            reg_file[7886] <= 8'h00
            reg_file[7887] <= 8'h00
            reg_file[7888] <= 8'h00
            reg_file[7889] <= 8'h00
            reg_file[7890] <= 8'h00
            reg_file[7891] <= 8'h00
            reg_file[7892] <= 8'h00
            reg_file[7893] <= 8'h00
            reg_file[7894] <= 8'h00
            reg_file[7895] <= 8'h00
            reg_file[7896] <= 8'h00
            reg_file[7897] <= 8'h00
            reg_file[7898] <= 8'h00
            reg_file[7899] <= 8'h00
            reg_file[7900] <= 8'h00
            reg_file[7901] <= 8'h00
            reg_file[7902] <= 8'h00
            reg_file[7903] <= 8'h00
            reg_file[7904] <= 8'h00
            reg_file[7905] <= 8'h00
            reg_file[7906] <= 8'h00
            reg_file[7907] <= 8'h00
            reg_file[7908] <= 8'h00
            reg_file[7909] <= 8'h00
            reg_file[7910] <= 8'h00
            reg_file[7911] <= 8'h00
            reg_file[7912] <= 8'h00
            reg_file[7913] <= 8'h00
            reg_file[7914] <= 8'h00
            reg_file[7915] <= 8'h00
            reg_file[7916] <= 8'h00
            reg_file[7917] <= 8'h00
            reg_file[7918] <= 8'h00
            reg_file[7919] <= 8'h00
            reg_file[7920] <= 8'h00
            reg_file[7921] <= 8'h00
            reg_file[7922] <= 8'h00
            reg_file[7923] <= 8'h00
            reg_file[7924] <= 8'h00
            reg_file[7925] <= 8'h00
            reg_file[7926] <= 8'h00
            reg_file[7927] <= 8'h00
            reg_file[7928] <= 8'h00
            reg_file[7929] <= 8'h00
            reg_file[7930] <= 8'h00
            reg_file[7931] <= 8'h00
            reg_file[7932] <= 8'h00
            reg_file[7933] <= 8'h00
            reg_file[7934] <= 8'h00
            reg_file[7935] <= 8'h00
            reg_file[7936] <= 8'h00
            reg_file[7937] <= 8'h00
            reg_file[7938] <= 8'h00
            reg_file[7939] <= 8'h00
            reg_file[7940] <= 8'h00
            reg_file[7941] <= 8'h00
            reg_file[7942] <= 8'h00
            reg_file[7943] <= 8'h00
            reg_file[7944] <= 8'h00
            reg_file[7945] <= 8'h00
            reg_file[7946] <= 8'h00
            reg_file[7947] <= 8'h00
            reg_file[7948] <= 8'h00
            reg_file[7949] <= 8'h00
            reg_file[7950] <= 8'h00
            reg_file[7951] <= 8'h00
            reg_file[7952] <= 8'h00
            reg_file[7953] <= 8'h00
            reg_file[7954] <= 8'h00
            reg_file[7955] <= 8'h00
            reg_file[7956] <= 8'h00
            reg_file[7957] <= 8'h00
            reg_file[7958] <= 8'h00
            reg_file[7959] <= 8'h00
            reg_file[7960] <= 8'h00
            reg_file[7961] <= 8'h00
            reg_file[7962] <= 8'h00
            reg_file[7963] <= 8'h00
            reg_file[7964] <= 8'h00
            reg_file[7965] <= 8'h00
            reg_file[7966] <= 8'h00
            reg_file[7967] <= 8'h00
            reg_file[7968] <= 8'h00
            reg_file[7969] <= 8'h00
            reg_file[7970] <= 8'h00
            reg_file[7971] <= 8'h00
            reg_file[7972] <= 8'h00
            reg_file[7973] <= 8'h00
            reg_file[7974] <= 8'h00
            reg_file[7975] <= 8'h00
            reg_file[7976] <= 8'h00
            reg_file[7977] <= 8'h00
            reg_file[7978] <= 8'h00
            reg_file[7979] <= 8'h00
            reg_file[7980] <= 8'h00
            reg_file[7981] <= 8'h00
            reg_file[7982] <= 8'h00
            reg_file[7983] <= 8'h00
            reg_file[7984] <= 8'h00
            reg_file[7985] <= 8'h00
            reg_file[7986] <= 8'h00
            reg_file[7987] <= 8'h00
            reg_file[7988] <= 8'h00
            reg_file[7989] <= 8'h00
            reg_file[7990] <= 8'h00
            reg_file[7991] <= 8'h00
            reg_file[7992] <= 8'h00
            reg_file[7993] <= 8'h00
            reg_file[7994] <= 8'h00
            reg_file[7995] <= 8'h00
            reg_file[7996] <= 8'h00
            reg_file[7997] <= 8'h00
            reg_file[7998] <= 8'h00
            reg_file[7999] <= 8'h00
            reg_file[8000] <= 8'h00
            reg_file[8001] <= 8'h00
            reg_file[8002] <= 8'h00
            reg_file[8003] <= 8'h00
            reg_file[8004] <= 8'h00
            reg_file[8005] <= 8'h00
            reg_file[8006] <= 8'h00
            reg_file[8007] <= 8'h00
            reg_file[8008] <= 8'h00
            reg_file[8009] <= 8'h00
            reg_file[8010] <= 8'h00
            reg_file[8011] <= 8'h00
            reg_file[8012] <= 8'h00
            reg_file[8013] <= 8'h00
            reg_file[8014] <= 8'h00
            reg_file[8015] <= 8'h00
            reg_file[8016] <= 8'h00
            reg_file[8017] <= 8'h00
            reg_file[8018] <= 8'h00
            reg_file[8019] <= 8'h00
            reg_file[8020] <= 8'h00
            reg_file[8021] <= 8'h00
            reg_file[8022] <= 8'h00
            reg_file[8023] <= 8'h00
            reg_file[8024] <= 8'h00
            reg_file[8025] <= 8'h00
            reg_file[8026] <= 8'h00
            reg_file[8027] <= 8'h00
            reg_file[8028] <= 8'h00
            reg_file[8029] <= 8'h00
            reg_file[8030] <= 8'h00
            reg_file[8031] <= 8'h00
            reg_file[8032] <= 8'h00
            reg_file[8033] <= 8'h00
            reg_file[8034] <= 8'h00
            reg_file[8035] <= 8'h00
            reg_file[8036] <= 8'h00
            reg_file[8037] <= 8'h00
            reg_file[8038] <= 8'h00
            reg_file[8039] <= 8'h00
            reg_file[8040] <= 8'h00
            reg_file[8041] <= 8'h00
            reg_file[8042] <= 8'h00
            reg_file[8043] <= 8'h00
            reg_file[8044] <= 8'h00
            reg_file[8045] <= 8'h00
            reg_file[8046] <= 8'h00
            reg_file[8047] <= 8'h00
            reg_file[8048] <= 8'h00
            reg_file[8049] <= 8'h00
            reg_file[8050] <= 8'h00
            reg_file[8051] <= 8'h00
            reg_file[8052] <= 8'h00
            reg_file[8053] <= 8'h00
            reg_file[8054] <= 8'h00
            reg_file[8055] <= 8'h00
            reg_file[8056] <= 8'h00
            reg_file[8057] <= 8'h00
            reg_file[8058] <= 8'h00
            reg_file[8059] <= 8'h00
            reg_file[8060] <= 8'h00
            reg_file[8061] <= 8'h00
            reg_file[8062] <= 8'h00
            reg_file[8063] <= 8'h00
            reg_file[8064] <= 8'h00
            reg_file[8065] <= 8'h00
            reg_file[8066] <= 8'h00
            reg_file[8067] <= 8'h00
            reg_file[8068] <= 8'h00
            reg_file[8069] <= 8'h00
            reg_file[8070] <= 8'h00
            reg_file[8071] <= 8'h00
            reg_file[8072] <= 8'h00
            reg_file[8073] <= 8'h00
            reg_file[8074] <= 8'h00
            reg_file[8075] <= 8'h00
            reg_file[8076] <= 8'h00
            reg_file[8077] <= 8'h00
            reg_file[8078] <= 8'h00
            reg_file[8079] <= 8'h00
            reg_file[8080] <= 8'h00
            reg_file[8081] <= 8'h00
            reg_file[8082] <= 8'h00
            reg_file[8083] <= 8'h00
            reg_file[8084] <= 8'h00
            reg_file[8085] <= 8'h00
            reg_file[8086] <= 8'h00
            reg_file[8087] <= 8'h00
            reg_file[8088] <= 8'h00
            reg_file[8089] <= 8'h00
            reg_file[8090] <= 8'h00
            reg_file[8091] <= 8'h00
            reg_file[8092] <= 8'h00
            reg_file[8093] <= 8'h00
            reg_file[8094] <= 8'h00
            reg_file[8095] <= 8'h00
            reg_file[8096] <= 8'h00
            reg_file[8097] <= 8'h00
            reg_file[8098] <= 8'h00
            reg_file[8099] <= 8'h00
            reg_file[8100] <= 8'h00
            reg_file[8101] <= 8'h00
            reg_file[8102] <= 8'h00
            reg_file[8103] <= 8'h00
            reg_file[8104] <= 8'h00
            reg_file[8105] <= 8'h00
            reg_file[8106] <= 8'h00
            reg_file[8107] <= 8'h00
            reg_file[8108] <= 8'h00
            reg_file[8109] <= 8'h00
            reg_file[8110] <= 8'h00
            reg_file[8111] <= 8'h00
            reg_file[8112] <= 8'h00
            reg_file[8113] <= 8'h00
            reg_file[8114] <= 8'h00
            reg_file[8115] <= 8'h00
            reg_file[8116] <= 8'h00
            reg_file[8117] <= 8'h00
            reg_file[8118] <= 8'h00
            reg_file[8119] <= 8'h00
            reg_file[8120] <= 8'h00
            reg_file[8121] <= 8'h00
            reg_file[8122] <= 8'h00
            reg_file[8123] <= 8'h00
            reg_file[8124] <= 8'h00
            reg_file[8125] <= 8'h00
            reg_file[8126] <= 8'h00
            reg_file[8127] <= 8'h00
            reg_file[8128] <= 8'h00
            reg_file[8129] <= 8'h00
            reg_file[8130] <= 8'h00
            reg_file[8131] <= 8'h00
            reg_file[8132] <= 8'h00
            reg_file[8133] <= 8'h00
            reg_file[8134] <= 8'h00
            reg_file[8135] <= 8'h00
            reg_file[8136] <= 8'h00
            reg_file[8137] <= 8'h00
            reg_file[8138] <= 8'h00
            reg_file[8139] <= 8'h00
            reg_file[8140] <= 8'h00
            reg_file[8141] <= 8'h00
            reg_file[8142] <= 8'h00
            reg_file[8143] <= 8'h00
            reg_file[8144] <= 8'h00
            reg_file[8145] <= 8'h00
            reg_file[8146] <= 8'h00
            reg_file[8147] <= 8'h00
            reg_file[8148] <= 8'h00
            reg_file[8149] <= 8'h00
            reg_file[8150] <= 8'h00
            reg_file[8151] <= 8'h00
            reg_file[8152] <= 8'h00
            reg_file[8153] <= 8'h00
            reg_file[8154] <= 8'h00
            reg_file[8155] <= 8'h00
            reg_file[8156] <= 8'h00
            reg_file[8157] <= 8'h00
            reg_file[8158] <= 8'h00
            reg_file[8159] <= 8'h00
            reg_file[8160] <= 8'h00
            reg_file[8161] <= 8'h00
            reg_file[8162] <= 8'h00
            reg_file[8163] <= 8'h00
            reg_file[8164] <= 8'h00
            reg_file[8165] <= 8'h00
            reg_file[8166] <= 8'h00
            reg_file[8167] <= 8'h00
            reg_file[8168] <= 8'h00
            reg_file[8169] <= 8'h00
            reg_file[8170] <= 8'h00
            reg_file[8171] <= 8'h00
            reg_file[8172] <= 8'h00
            reg_file[8173] <= 8'h00
            reg_file[8174] <= 8'h00
            reg_file[8175] <= 8'h00
            reg_file[8176] <= 8'h00
            reg_file[8177] <= 8'h00
            reg_file[8178] <= 8'h00
            reg_file[8179] <= 8'h00
            reg_file[8180] <= 8'h00
            reg_file[8181] <= 8'h00
            reg_file[8182] <= 8'h00
            reg_file[8183] <= 8'h00
            reg_file[8184] <= 8'h00
            reg_file[8185] <= 8'h00
            reg_file[8186] <= 8'h00
            reg_file[8187] <= 8'h00
            reg_file[8188] <= 8'h00
            reg_file[8189] <= 8'h00
            reg_file[8190] <= 8'h00
            reg_file[8191] <= 8'h00
            reg_file[8192] <= 8'h00
            reg_file[8193] <= 8'h00
            reg_file[8194] <= 8'h00
            reg_file[8195] <= 8'h00
            reg_file[8196] <= 8'h00
            reg_file[8197] <= 8'h00
            reg_file[8198] <= 8'h00
            reg_file[8199] <= 8'h00
            reg_file[8200] <= 8'h00
            reg_file[8201] <= 8'h00
            reg_file[8202] <= 8'h00
            reg_file[8203] <= 8'h00
            reg_file[8204] <= 8'h00
            reg_file[8205] <= 8'h00
            reg_file[8206] <= 8'h00
            reg_file[8207] <= 8'h00
            reg_file[8208] <= 8'h00
            reg_file[8209] <= 8'h00
            reg_file[8210] <= 8'h00
            reg_file[8211] <= 8'h00
            reg_file[8212] <= 8'h00
            reg_file[8213] <= 8'h00
            reg_file[8214] <= 8'h00
            reg_file[8215] <= 8'h00
            reg_file[8216] <= 8'h00
            reg_file[8217] <= 8'h00
            reg_file[8218] <= 8'h00
            reg_file[8219] <= 8'h00
            reg_file[8220] <= 8'h00
            reg_file[8221] <= 8'h00
            reg_file[8222] <= 8'h00
            reg_file[8223] <= 8'h00
            reg_file[8224] <= 8'h00
            reg_file[8225] <= 8'h00
            reg_file[8226] <= 8'h00
            reg_file[8227] <= 8'h00
            reg_file[8228] <= 8'h00
            reg_file[8229] <= 8'h00
            reg_file[8230] <= 8'h00
            reg_file[8231] <= 8'h00
            reg_file[8232] <= 8'h00
            reg_file[8233] <= 8'h00
            reg_file[8234] <= 8'h00
            reg_file[8235] <= 8'h00
            reg_file[8236] <= 8'h00
            reg_file[8237] <= 8'h00
            reg_file[8238] <= 8'h00
            reg_file[8239] <= 8'h00
            reg_file[8240] <= 8'h00
            reg_file[8241] <= 8'h00
            reg_file[8242] <= 8'h00
            reg_file[8243] <= 8'h00
            reg_file[8244] <= 8'h00
            reg_file[8245] <= 8'h00
            reg_file[8246] <= 8'h00
            reg_file[8247] <= 8'h00
            reg_file[8248] <= 8'h00
            reg_file[8249] <= 8'h00
            reg_file[8250] <= 8'h00
            reg_file[8251] <= 8'h00
            reg_file[8252] <= 8'h00
            reg_file[8253] <= 8'h00
            reg_file[8254] <= 8'h00
            reg_file[8255] <= 8'h00
            reg_file[8256] <= 8'h00
            reg_file[8257] <= 8'h00
            reg_file[8258] <= 8'h00
            reg_file[8259] <= 8'h00
            reg_file[8260] <= 8'h00
            reg_file[8261] <= 8'h00
            reg_file[8262] <= 8'h00
            reg_file[8263] <= 8'h00
            reg_file[8264] <= 8'h00
            reg_file[8265] <= 8'h00
            reg_file[8266] <= 8'h00
            reg_file[8267] <= 8'h00
            reg_file[8268] <= 8'h00
            reg_file[8269] <= 8'h00
            reg_file[8270] <= 8'h00
            reg_file[8271] <= 8'h00
            reg_file[8272] <= 8'h00
            reg_file[8273] <= 8'h00
            reg_file[8274] <= 8'h00
            reg_file[8275] <= 8'h00
            reg_file[8276] <= 8'h00
            reg_file[8277] <= 8'h00
            reg_file[8278] <= 8'h00
            reg_file[8279] <= 8'h00
            reg_file[8280] <= 8'h00
            reg_file[8281] <= 8'h00
            reg_file[8282] <= 8'h00
            reg_file[8283] <= 8'h00
            reg_file[8284] <= 8'h00
            reg_file[8285] <= 8'h00
            reg_file[8286] <= 8'h00
            reg_file[8287] <= 8'h00
            reg_file[8288] <= 8'h00
            reg_file[8289] <= 8'h00
            reg_file[8290] <= 8'h00
            reg_file[8291] <= 8'h00
            reg_file[8292] <= 8'h00
            reg_file[8293] <= 8'h00
            reg_file[8294] <= 8'h00
            reg_file[8295] <= 8'h00
            reg_file[8296] <= 8'h00
            reg_file[8297] <= 8'h00
            reg_file[8298] <= 8'h00
            reg_file[8299] <= 8'h00
            reg_file[8300] <= 8'h00
            reg_file[8301] <= 8'h00
            reg_file[8302] <= 8'h00
            reg_file[8303] <= 8'h00
            reg_file[8304] <= 8'h00
            reg_file[8305] <= 8'h00
            reg_file[8306] <= 8'h00
            reg_file[8307] <= 8'h00
            reg_file[8308] <= 8'h00
            reg_file[8309] <= 8'h00
            reg_file[8310] <= 8'h00
            reg_file[8311] <= 8'h00
            reg_file[8312] <= 8'h00
            reg_file[8313] <= 8'h00
            reg_file[8314] <= 8'h00
            reg_file[8315] <= 8'h00
            reg_file[8316] <= 8'h00
            reg_file[8317] <= 8'h00
            reg_file[8318] <= 8'h00
            reg_file[8319] <= 8'h00
            reg_file[8320] <= 8'h00
            reg_file[8321] <= 8'h00
            reg_file[8322] <= 8'h00
            reg_file[8323] <= 8'h00
            reg_file[8324] <= 8'h00
            reg_file[8325] <= 8'h00
            reg_file[8326] <= 8'h00
            reg_file[8327] <= 8'h00
            reg_file[8328] <= 8'h00
            reg_file[8329] <= 8'h00
            reg_file[8330] <= 8'h00
            reg_file[8331] <= 8'h00
            reg_file[8332] <= 8'h00
            reg_file[8333] <= 8'h00
            reg_file[8334] <= 8'h00
            reg_file[8335] <= 8'h00
            reg_file[8336] <= 8'h00
            reg_file[8337] <= 8'h00
            reg_file[8338] <= 8'h00
            reg_file[8339] <= 8'h00
            reg_file[8340] <= 8'h00
            reg_file[8341] <= 8'h00
            reg_file[8342] <= 8'h00
            reg_file[8343] <= 8'h00
            reg_file[8344] <= 8'h00
            reg_file[8345] <= 8'h00
            reg_file[8346] <= 8'h00
            reg_file[8347] <= 8'h00
            reg_file[8348] <= 8'h00
            reg_file[8349] <= 8'h00
            reg_file[8350] <= 8'h00
            reg_file[8351] <= 8'h00
            reg_file[8352] <= 8'h00
            reg_file[8353] <= 8'h00
            reg_file[8354] <= 8'h00
            reg_file[8355] <= 8'h00
            reg_file[8356] <= 8'h00
            reg_file[8357] <= 8'h00
            reg_file[8358] <= 8'h00
            reg_file[8359] <= 8'h00
            reg_file[8360] <= 8'h00
            reg_file[8361] <= 8'h00
            reg_file[8362] <= 8'h00
            reg_file[8363] <= 8'h00
            reg_file[8364] <= 8'h00
            reg_file[8365] <= 8'h00
            reg_file[8366] <= 8'h00
            reg_file[8367] <= 8'h00
            reg_file[8368] <= 8'h00
            reg_file[8369] <= 8'h00
            reg_file[8370] <= 8'h00
            reg_file[8371] <= 8'h00
            reg_file[8372] <= 8'h00
            reg_file[8373] <= 8'h00
            reg_file[8374] <= 8'h00
            reg_file[8375] <= 8'h00
            reg_file[8376] <= 8'h00
            reg_file[8377] <= 8'h00
            reg_file[8378] <= 8'h00
            reg_file[8379] <= 8'h00
            reg_file[8380] <= 8'h00
            reg_file[8381] <= 8'h00
            reg_file[8382] <= 8'h00
            reg_file[8383] <= 8'h00
            reg_file[8384] <= 8'h00
            reg_file[8385] <= 8'h00
            reg_file[8386] <= 8'h00
            reg_file[8387] <= 8'h00
            reg_file[8388] <= 8'h00
            reg_file[8389] <= 8'h00
            reg_file[8390] <= 8'h00
            reg_file[8391] <= 8'h00
            reg_file[8392] <= 8'h00
            reg_file[8393] <= 8'h00
            reg_file[8394] <= 8'h00
            reg_file[8395] <= 8'h00
            reg_file[8396] <= 8'h00
            reg_file[8397] <= 8'h00
            reg_file[8398] <= 8'h00
            reg_file[8399] <= 8'h00
            reg_file[8400] <= 8'h00
            reg_file[8401] <= 8'h00
            reg_file[8402] <= 8'h00
            reg_file[8403] <= 8'h00
            reg_file[8404] <= 8'h00
            reg_file[8405] <= 8'h00
            reg_file[8406] <= 8'h00
            reg_file[8407] <= 8'h00
            reg_file[8408] <= 8'h00
            reg_file[8409] <= 8'h00
            reg_file[8410] <= 8'h00
            reg_file[8411] <= 8'h00
            reg_file[8412] <= 8'h00
            reg_file[8413] <= 8'h00
            reg_file[8414] <= 8'h00
            reg_file[8415] <= 8'h00
            reg_file[8416] <= 8'h00
            reg_file[8417] <= 8'h00
            reg_file[8418] <= 8'h00
            reg_file[8419] <= 8'h00
            reg_file[8420] <= 8'h00
            reg_file[8421] <= 8'h00
            reg_file[8422] <= 8'h00
            reg_file[8423] <= 8'h00
            reg_file[8424] <= 8'h00
            reg_file[8425] <= 8'h00
            reg_file[8426] <= 8'h00
            reg_file[8427] <= 8'h00
            reg_file[8428] <= 8'h00
            reg_file[8429] <= 8'h00
            reg_file[8430] <= 8'h00
            reg_file[8431] <= 8'h00
            reg_file[8432] <= 8'h00
            reg_file[8433] <= 8'h00
            reg_file[8434] <= 8'h00
            reg_file[8435] <= 8'h00
            reg_file[8436] <= 8'h00
            reg_file[8437] <= 8'h00
            reg_file[8438] <= 8'h00
            reg_file[8439] <= 8'h00
            reg_file[8440] <= 8'h00
            reg_file[8441] <= 8'h00
            reg_file[8442] <= 8'h00
            reg_file[8443] <= 8'h00
            reg_file[8444] <= 8'h00
            reg_file[8445] <= 8'h00
            reg_file[8446] <= 8'h00
            reg_file[8447] <= 8'h00
            reg_file[8448] <= 8'h00
            reg_file[8449] <= 8'h00
            reg_file[8450] <= 8'h00
            reg_file[8451] <= 8'h00
            reg_file[8452] <= 8'h00
            reg_file[8453] <= 8'h00
            reg_file[8454] <= 8'h00
            reg_file[8455] <= 8'h00
            reg_file[8456] <= 8'h00
            reg_file[8457] <= 8'h00
            reg_file[8458] <= 8'h00
            reg_file[8459] <= 8'h00
            reg_file[8460] <= 8'h00
            reg_file[8461] <= 8'h00
            reg_file[8462] <= 8'h00
            reg_file[8463] <= 8'h00
            reg_file[8464] <= 8'h00
            reg_file[8465] <= 8'h00
            reg_file[8466] <= 8'h00
            reg_file[8467] <= 8'h00
            reg_file[8468] <= 8'h00
            reg_file[8469] <= 8'h00
            reg_file[8470] <= 8'h00
            reg_file[8471] <= 8'h00
            reg_file[8472] <= 8'h00
            reg_file[8473] <= 8'h00
            reg_file[8474] <= 8'h00
            reg_file[8475] <= 8'h00
            reg_file[8476] <= 8'h00
            reg_file[8477] <= 8'h00
            reg_file[8478] <= 8'h00
            reg_file[8479] <= 8'h00
            reg_file[8480] <= 8'h00
            reg_file[8481] <= 8'h00
            reg_file[8482] <= 8'h00
            reg_file[8483] <= 8'h00
            reg_file[8484] <= 8'h00
            reg_file[8485] <= 8'h00
            reg_file[8486] <= 8'h00
            reg_file[8487] <= 8'h00
            reg_file[8488] <= 8'h00
            reg_file[8489] <= 8'h00
            reg_file[8490] <= 8'h00
            reg_file[8491] <= 8'h00
            reg_file[8492] <= 8'h00
            reg_file[8493] <= 8'h00
            reg_file[8494] <= 8'h00
            reg_file[8495] <= 8'h00
            reg_file[8496] <= 8'h00
            reg_file[8497] <= 8'h00
            reg_file[8498] <= 8'h00
            reg_file[8499] <= 8'h00
            reg_file[8500] <= 8'h00
            reg_file[8501] <= 8'h00
            reg_file[8502] <= 8'h00
            reg_file[8503] <= 8'h00
            reg_file[8504] <= 8'h00
            reg_file[8505] <= 8'h00
            reg_file[8506] <= 8'h00
            reg_file[8507] <= 8'h00
            reg_file[8508] <= 8'h00
            reg_file[8509] <= 8'h00
            reg_file[8510] <= 8'h00
            reg_file[8511] <= 8'h00
            reg_file[8512] <= 8'h00
            reg_file[8513] <= 8'h00
            reg_file[8514] <= 8'h00
            reg_file[8515] <= 8'h00
            reg_file[8516] <= 8'h00
            reg_file[8517] <= 8'h00
            reg_file[8518] <= 8'h00
            reg_file[8519] <= 8'h00
            reg_file[8520] <= 8'h00
            reg_file[8521] <= 8'h00
            reg_file[8522] <= 8'h00
            reg_file[8523] <= 8'h00
            reg_file[8524] <= 8'h00
            reg_file[8525] <= 8'h00
            reg_file[8526] <= 8'h00
            reg_file[8527] <= 8'h00
            reg_file[8528] <= 8'h00
            reg_file[8529] <= 8'h00
            reg_file[8530] <= 8'h00
            reg_file[8531] <= 8'h00
            reg_file[8532] <= 8'h00
            reg_file[8533] <= 8'h00
            reg_file[8534] <= 8'h00
            reg_file[8535] <= 8'h00
            reg_file[8536] <= 8'h00
            reg_file[8537] <= 8'h00
            reg_file[8538] <= 8'h00
            reg_file[8539] <= 8'h00
            reg_file[8540] <= 8'h00
            reg_file[8541] <= 8'h00
            reg_file[8542] <= 8'h00
            reg_file[8543] <= 8'h00
            reg_file[8544] <= 8'h00
            reg_file[8545] <= 8'h00
            reg_file[8546] <= 8'h00
            reg_file[8547] <= 8'h00
            reg_file[8548] <= 8'h00
            reg_file[8549] <= 8'h00
            reg_file[8550] <= 8'h00
            reg_file[8551] <= 8'h00
            reg_file[8552] <= 8'h00
            reg_file[8553] <= 8'h00
            reg_file[8554] <= 8'h00
            reg_file[8555] <= 8'h00
            reg_file[8556] <= 8'h00
            reg_file[8557] <= 8'h00
            reg_file[8558] <= 8'h00
            reg_file[8559] <= 8'h00
            reg_file[8560] <= 8'h00
            reg_file[8561] <= 8'h00
            reg_file[8562] <= 8'h00
            reg_file[8563] <= 8'h00
            reg_file[8564] <= 8'h00
            reg_file[8565] <= 8'h00
            reg_file[8566] <= 8'h00
            reg_file[8567] <= 8'h00
            reg_file[8568] <= 8'h00
            reg_file[8569] <= 8'h00
            reg_file[8570] <= 8'h00
            reg_file[8571] <= 8'h00
            reg_file[8572] <= 8'h00
            reg_file[8573] <= 8'h00
            reg_file[8574] <= 8'h00
            reg_file[8575] <= 8'h00
            reg_file[8576] <= 8'h00
            reg_file[8577] <= 8'h00
            reg_file[8578] <= 8'h00
            reg_file[8579] <= 8'h00
            reg_file[8580] <= 8'h00
            reg_file[8581] <= 8'h00
            reg_file[8582] <= 8'h00
            reg_file[8583] <= 8'h00
            reg_file[8584] <= 8'h00
            reg_file[8585] <= 8'h00
            reg_file[8586] <= 8'h00
            reg_file[8587] <= 8'h00
            reg_file[8588] <= 8'h00
            reg_file[8589] <= 8'h00
            reg_file[8590] <= 8'h00
            reg_file[8591] <= 8'h00
            reg_file[8592] <= 8'h00
            reg_file[8593] <= 8'h00
            reg_file[8594] <= 8'h00
            reg_file[8595] <= 8'h00
            reg_file[8596] <= 8'h00
            reg_file[8597] <= 8'h00
            reg_file[8598] <= 8'h00
            reg_file[8599] <= 8'h00
            reg_file[8600] <= 8'h00
            reg_file[8601] <= 8'h00
            reg_file[8602] <= 8'h00
            reg_file[8603] <= 8'h00
            reg_file[8604] <= 8'h00
            reg_file[8605] <= 8'h00
            reg_file[8606] <= 8'h00
            reg_file[8607] <= 8'h00
            reg_file[8608] <= 8'h00
            reg_file[8609] <= 8'h00
            reg_file[8610] <= 8'h00
            reg_file[8611] <= 8'h00
            reg_file[8612] <= 8'h00
            reg_file[8613] <= 8'h00
            reg_file[8614] <= 8'h00
            reg_file[8615] <= 8'h00
            reg_file[8616] <= 8'h00
            reg_file[8617] <= 8'h00
            reg_file[8618] <= 8'h00
            reg_file[8619] <= 8'h00
            reg_file[8620] <= 8'h00
            reg_file[8621] <= 8'h00
            reg_file[8622] <= 8'h00
            reg_file[8623] <= 8'h00
            reg_file[8624] <= 8'h00
            reg_file[8625] <= 8'h00
            reg_file[8626] <= 8'h00
            reg_file[8627] <= 8'h00
            reg_file[8628] <= 8'h00
            reg_file[8629] <= 8'h00
            reg_file[8630] <= 8'h00
            reg_file[8631] <= 8'h00
            reg_file[8632] <= 8'h00
            reg_file[8633] <= 8'h00
            reg_file[8634] <= 8'h00
            reg_file[8635] <= 8'h00
            reg_file[8636] <= 8'h00
            reg_file[8637] <= 8'h00
            reg_file[8638] <= 8'h00
            reg_file[8639] <= 8'h00
            reg_file[8640] <= 8'h00
            reg_file[8641] <= 8'h00
            reg_file[8642] <= 8'h00
            reg_file[8643] <= 8'h00
            reg_file[8644] <= 8'h00
            reg_file[8645] <= 8'h00
            reg_file[8646] <= 8'h00
            reg_file[8647] <= 8'h00
            reg_file[8648] <= 8'h00
            reg_file[8649] <= 8'h00
            reg_file[8650] <= 8'h00
            reg_file[8651] <= 8'h00
            reg_file[8652] <= 8'h00
            reg_file[8653] <= 8'h00
            reg_file[8654] <= 8'h00
            reg_file[8655] <= 8'h00
            reg_file[8656] <= 8'h00
            reg_file[8657] <= 8'h00
            reg_file[8658] <= 8'h00
            reg_file[8659] <= 8'h00
            reg_file[8660] <= 8'h00
            reg_file[8661] <= 8'h00
            reg_file[8662] <= 8'h00
            reg_file[8663] <= 8'h00
            reg_file[8664] <= 8'h00
            reg_file[8665] <= 8'h00
            reg_file[8666] <= 8'h00
            reg_file[8667] <= 8'h00
            reg_file[8668] <= 8'h00
            reg_file[8669] <= 8'h00
            reg_file[8670] <= 8'h00
            reg_file[8671] <= 8'h00
            reg_file[8672] <= 8'h00
            reg_file[8673] <= 8'h00
            reg_file[8674] <= 8'h00
            reg_file[8675] <= 8'h00
            reg_file[8676] <= 8'h00
            reg_file[8677] <= 8'h00
            reg_file[8678] <= 8'h00
            reg_file[8679] <= 8'h00
            reg_file[8680] <= 8'h00
            reg_file[8681] <= 8'h00
            reg_file[8682] <= 8'h00
            reg_file[8683] <= 8'h00
            reg_file[8684] <= 8'h00
            reg_file[8685] <= 8'h00
            reg_file[8686] <= 8'h00
            reg_file[8687] <= 8'h00
            reg_file[8688] <= 8'h00
            reg_file[8689] <= 8'h00
            reg_file[8690] <= 8'h00
            reg_file[8691] <= 8'h00
            reg_file[8692] <= 8'h00
            reg_file[8693] <= 8'h00
            reg_file[8694] <= 8'h00
            reg_file[8695] <= 8'h00
            reg_file[8696] <= 8'h00
            reg_file[8697] <= 8'h00
            reg_file[8698] <= 8'h00
            reg_file[8699] <= 8'h00
            reg_file[8700] <= 8'h00
            reg_file[8701] <= 8'h00
            reg_file[8702] <= 8'h00
            reg_file[8703] <= 8'h00
            reg_file[8704] <= 8'h00
            reg_file[8705] <= 8'h00
            reg_file[8706] <= 8'h00
            reg_file[8707] <= 8'h00
            reg_file[8708] <= 8'h00
            reg_file[8709] <= 8'h00
            reg_file[8710] <= 8'h00
            reg_file[8711] <= 8'h00
            reg_file[8712] <= 8'h00
            reg_file[8713] <= 8'h00
            reg_file[8714] <= 8'h00
            reg_file[8715] <= 8'h00
            reg_file[8716] <= 8'h00
            reg_file[8717] <= 8'h00
            reg_file[8718] <= 8'h00
            reg_file[8719] <= 8'h00
            reg_file[8720] <= 8'h00
            reg_file[8721] <= 8'h00
            reg_file[8722] <= 8'h00
            reg_file[8723] <= 8'h00
            reg_file[8724] <= 8'h00
            reg_file[8725] <= 8'h00
            reg_file[8726] <= 8'h00
            reg_file[8727] <= 8'h00
            reg_file[8728] <= 8'h00
            reg_file[8729] <= 8'h00
            reg_file[8730] <= 8'h00
            reg_file[8731] <= 8'h00
            reg_file[8732] <= 8'h00
            reg_file[8733] <= 8'h00
            reg_file[8734] <= 8'h00
            reg_file[8735] <= 8'h00
            reg_file[8736] <= 8'h00
            reg_file[8737] <= 8'h00
            reg_file[8738] <= 8'h00
            reg_file[8739] <= 8'h00
            reg_file[8740] <= 8'h00
            reg_file[8741] <= 8'h00
            reg_file[8742] <= 8'h00
            reg_file[8743] <= 8'h00
            reg_file[8744] <= 8'h00
            reg_file[8745] <= 8'h00
            reg_file[8746] <= 8'h00
            reg_file[8747] <= 8'h00
            reg_file[8748] <= 8'h00
            reg_file[8749] <= 8'h00
            reg_file[8750] <= 8'h00
            reg_file[8751] <= 8'h00
            reg_file[8752] <= 8'h00
            reg_file[8753] <= 8'h00
            reg_file[8754] <= 8'h00
            reg_file[8755] <= 8'h00
            reg_file[8756] <= 8'h00
            reg_file[8757] <= 8'h00
            reg_file[8758] <= 8'h00
            reg_file[8759] <= 8'h00
            reg_file[8760] <= 8'h00
            reg_file[8761] <= 8'h00
            reg_file[8762] <= 8'h00
            reg_file[8763] <= 8'h00
            reg_file[8764] <= 8'h00
            reg_file[8765] <= 8'h00
            reg_file[8766] <= 8'h00
            reg_file[8767] <= 8'h00
            reg_file[8768] <= 8'h00
            reg_file[8769] <= 8'h00
            reg_file[8770] <= 8'h00
            reg_file[8771] <= 8'h00
            reg_file[8772] <= 8'h00
            reg_file[8773] <= 8'h00
            reg_file[8774] <= 8'h00
            reg_file[8775] <= 8'h00
            reg_file[8776] <= 8'h00
            reg_file[8777] <= 8'h00
            reg_file[8778] <= 8'h00
            reg_file[8779] <= 8'h00
            reg_file[8780] <= 8'h00
            reg_file[8781] <= 8'h00
            reg_file[8782] <= 8'h00
            reg_file[8783] <= 8'h00
            reg_file[8784] <= 8'h00
            reg_file[8785] <= 8'h00
            reg_file[8786] <= 8'h00
            reg_file[8787] <= 8'h00
            reg_file[8788] <= 8'h00
            reg_file[8789] <= 8'h00
            reg_file[8790] <= 8'h00
            reg_file[8791] <= 8'h00
            reg_file[8792] <= 8'h00
            reg_file[8793] <= 8'h00
            reg_file[8794] <= 8'h00
            reg_file[8795] <= 8'h00
            reg_file[8796] <= 8'h00
            reg_file[8797] <= 8'h00
            reg_file[8798] <= 8'h00
            reg_file[8799] <= 8'h00
            reg_file[8800] <= 8'h00
            reg_file[8801] <= 8'h00
            reg_file[8802] <= 8'h00
            reg_file[8803] <= 8'h00
            reg_file[8804] <= 8'h00
            reg_file[8805] <= 8'h00
            reg_file[8806] <= 8'h00
            reg_file[8807] <= 8'h00
            reg_file[8808] <= 8'h00
            reg_file[8809] <= 8'h00
            reg_file[8810] <= 8'h00
            reg_file[8811] <= 8'h00
            reg_file[8812] <= 8'h00
            reg_file[8813] <= 8'h00
            reg_file[8814] <= 8'h00
            reg_file[8815] <= 8'h00
            reg_file[8816] <= 8'h00
            reg_file[8817] <= 8'h00
            reg_file[8818] <= 8'h00
            reg_file[8819] <= 8'h00
            reg_file[8820] <= 8'h00
            reg_file[8821] <= 8'h00
            reg_file[8822] <= 8'h00
            reg_file[8823] <= 8'h00
            reg_file[8824] <= 8'h00
            reg_file[8825] <= 8'h00
            reg_file[8826] <= 8'h00
            reg_file[8827] <= 8'h00
            reg_file[8828] <= 8'h00
            reg_file[8829] <= 8'h00
            reg_file[8830] <= 8'h00
            reg_file[8831] <= 8'h00
            reg_file[8832] <= 8'h00
            reg_file[8833] <= 8'h00
            reg_file[8834] <= 8'h00
            reg_file[8835] <= 8'h00
            reg_file[8836] <= 8'h00
            reg_file[8837] <= 8'h00
            reg_file[8838] <= 8'h00
            reg_file[8839] <= 8'h00
            reg_file[8840] <= 8'h00
            reg_file[8841] <= 8'h00
            reg_file[8842] <= 8'h00
            reg_file[8843] <= 8'h00
            reg_file[8844] <= 8'h00
            reg_file[8845] <= 8'h00
            reg_file[8846] <= 8'h00
            reg_file[8847] <= 8'h00
            reg_file[8848] <= 8'h00
            reg_file[8849] <= 8'h00
            reg_file[8850] <= 8'h00
            reg_file[8851] <= 8'h00
            reg_file[8852] <= 8'h00
            reg_file[8853] <= 8'h00
            reg_file[8854] <= 8'h00
            reg_file[8855] <= 8'h00
            reg_file[8856] <= 8'h00
            reg_file[8857] <= 8'h00
            reg_file[8858] <= 8'h00
            reg_file[8859] <= 8'h00
            reg_file[8860] <= 8'h00
            reg_file[8861] <= 8'h00
            reg_file[8862] <= 8'h00
            reg_file[8863] <= 8'h00
            reg_file[8864] <= 8'h00
            reg_file[8865] <= 8'h00
            reg_file[8866] <= 8'h00
            reg_file[8867] <= 8'h00
            reg_file[8868] <= 8'h00
            reg_file[8869] <= 8'h00
            reg_file[8870] <= 8'h00
            reg_file[8871] <= 8'h00
            reg_file[8872] <= 8'h00
            reg_file[8873] <= 8'h00
            reg_file[8874] <= 8'h00
            reg_file[8875] <= 8'h00
            reg_file[8876] <= 8'h00
            reg_file[8877] <= 8'h00
            reg_file[8878] <= 8'h00
            reg_file[8879] <= 8'h00
            reg_file[8880] <= 8'h00
            reg_file[8881] <= 8'h00
            reg_file[8882] <= 8'h00
            reg_file[8883] <= 8'h00
            reg_file[8884] <= 8'h00
            reg_file[8885] <= 8'h00
            reg_file[8886] <= 8'h00
            reg_file[8887] <= 8'h00
            reg_file[8888] <= 8'h00
            reg_file[8889] <= 8'h00
            reg_file[8890] <= 8'h00
            reg_file[8891] <= 8'h00
            reg_file[8892] <= 8'h00
            reg_file[8893] <= 8'h00
            reg_file[8894] <= 8'h00
            reg_file[8895] <= 8'h00
            reg_file[8896] <= 8'h00
            reg_file[8897] <= 8'h00
            reg_file[8898] <= 8'h00
            reg_file[8899] <= 8'h00
            reg_file[8900] <= 8'h00
            reg_file[8901] <= 8'h00
            reg_file[8902] <= 8'h00
            reg_file[8903] <= 8'h00
            reg_file[8904] <= 8'h00
            reg_file[8905] <= 8'h00
            reg_file[8906] <= 8'h00
            reg_file[8907] <= 8'h00
            reg_file[8908] <= 8'h00
            reg_file[8909] <= 8'h00
            reg_file[8910] <= 8'h00
            reg_file[8911] <= 8'h00
            reg_file[8912] <= 8'h00
            reg_file[8913] <= 8'h00
            reg_file[8914] <= 8'h00
            reg_file[8915] <= 8'h00
            reg_file[8916] <= 8'h00
            reg_file[8917] <= 8'h00
            reg_file[8918] <= 8'h00
            reg_file[8919] <= 8'h00
            reg_file[8920] <= 8'h00
            reg_file[8921] <= 8'h00
            reg_file[8922] <= 8'h00
            reg_file[8923] <= 8'h00
            reg_file[8924] <= 8'h00
            reg_file[8925] <= 8'h00
            reg_file[8926] <= 8'h00
            reg_file[8927] <= 8'h00
            reg_file[8928] <= 8'h00
            reg_file[8929] <= 8'h00
            reg_file[8930] <= 8'h00
            reg_file[8931] <= 8'h00
            reg_file[8932] <= 8'h00
            reg_file[8933] <= 8'h00
            reg_file[8934] <= 8'h00
            reg_file[8935] <= 8'h00
            reg_file[8936] <= 8'h00
            reg_file[8937] <= 8'h00
            reg_file[8938] <= 8'h00
            reg_file[8939] <= 8'h00
            reg_file[8940] <= 8'h00
            reg_file[8941] <= 8'h00
            reg_file[8942] <= 8'h00
            reg_file[8943] <= 8'h00
            reg_file[8944] <= 8'h00
            reg_file[8945] <= 8'h00
            reg_file[8946] <= 8'h00
            reg_file[8947] <= 8'h00
            reg_file[8948] <= 8'h00
            reg_file[8949] <= 8'h00
            reg_file[8950] <= 8'h00
            reg_file[8951] <= 8'h00
            reg_file[8952] <= 8'h00
            reg_file[8953] <= 8'h00
            reg_file[8954] <= 8'h00
            reg_file[8955] <= 8'h00
            reg_file[8956] <= 8'h00
            reg_file[8957] <= 8'h00
            reg_file[8958] <= 8'h00
            reg_file[8959] <= 8'h00
            reg_file[8960] <= 8'h00
            reg_file[8961] <= 8'h00
            reg_file[8962] <= 8'h00
            reg_file[8963] <= 8'h00
            reg_file[8964] <= 8'h00
            reg_file[8965] <= 8'h00
            reg_file[8966] <= 8'h00
            reg_file[8967] <= 8'h00
            reg_file[8968] <= 8'h00
            reg_file[8969] <= 8'h00
            reg_file[8970] <= 8'h00
            reg_file[8971] <= 8'h00
            reg_file[8972] <= 8'h00
            reg_file[8973] <= 8'h00
            reg_file[8974] <= 8'h00
            reg_file[8975] <= 8'h00
            reg_file[8976] <= 8'h00
            reg_file[8977] <= 8'h00
            reg_file[8978] <= 8'h00
            reg_file[8979] <= 8'h00
            reg_file[8980] <= 8'h00
            reg_file[8981] <= 8'h00
            reg_file[8982] <= 8'h00
            reg_file[8983] <= 8'h00
            reg_file[8984] <= 8'h00
            reg_file[8985] <= 8'h00
            reg_file[8986] <= 8'h00
            reg_file[8987] <= 8'h00
            reg_file[8988] <= 8'h00
            reg_file[8989] <= 8'h00
            reg_file[8990] <= 8'h00
            reg_file[8991] <= 8'h00
            reg_file[8992] <= 8'h00
            reg_file[8993] <= 8'h00
            reg_file[8994] <= 8'h00
            reg_file[8995] <= 8'h00
            reg_file[8996] <= 8'h00
            reg_file[8997] <= 8'h00
            reg_file[8998] <= 8'h00
            reg_file[8999] <= 8'h00
            reg_file[9000] <= 8'h00
            reg_file[9001] <= 8'h00
            reg_file[9002] <= 8'h00
            reg_file[9003] <= 8'h00
            reg_file[9004] <= 8'h00
            reg_file[9005] <= 8'h00
            reg_file[9006] <= 8'h00
            reg_file[9007] <= 8'h00
            reg_file[9008] <= 8'h00
            reg_file[9009] <= 8'h00
            reg_file[9010] <= 8'h00
            reg_file[9011] <= 8'h00
            reg_file[9012] <= 8'h00
            reg_file[9013] <= 8'h00
            reg_file[9014] <= 8'h00
            reg_file[9015] <= 8'h00
            reg_file[9016] <= 8'h00
            reg_file[9017] <= 8'h00
            reg_file[9018] <= 8'h00
            reg_file[9019] <= 8'h00
            reg_file[9020] <= 8'h00
            reg_file[9021] <= 8'h00
            reg_file[9022] <= 8'h00
            reg_file[9023] <= 8'h00
            reg_file[9024] <= 8'h00
            reg_file[9025] <= 8'h00
            reg_file[9026] <= 8'h00
            reg_file[9027] <= 8'h00
            reg_file[9028] <= 8'h00
            reg_file[9029] <= 8'h00
            reg_file[9030] <= 8'h00
            reg_file[9031] <= 8'h00
            reg_file[9032] <= 8'h00
            reg_file[9033] <= 8'h00
            reg_file[9034] <= 8'h00
            reg_file[9035] <= 8'h00
            reg_file[9036] <= 8'h00
            reg_file[9037] <= 8'h00
            reg_file[9038] <= 8'h00
            reg_file[9039] <= 8'h00
            reg_file[9040] <= 8'h00
            reg_file[9041] <= 8'h00
            reg_file[9042] <= 8'h00
            reg_file[9043] <= 8'h00
            reg_file[9044] <= 8'h00
            reg_file[9045] <= 8'h00
            reg_file[9046] <= 8'h00
            reg_file[9047] <= 8'h00
            reg_file[9048] <= 8'h00
            reg_file[9049] <= 8'h00
            reg_file[9050] <= 8'h00
            reg_file[9051] <= 8'h00
            reg_file[9052] <= 8'h00
            reg_file[9053] <= 8'h00
            reg_file[9054] <= 8'h00
            reg_file[9055] <= 8'h00
            reg_file[9056] <= 8'h00
            reg_file[9057] <= 8'h00
            reg_file[9058] <= 8'h00
            reg_file[9059] <= 8'h00
            reg_file[9060] <= 8'h00
            reg_file[9061] <= 8'h00
            reg_file[9062] <= 8'h00
            reg_file[9063] <= 8'h00
            reg_file[9064] <= 8'h00
            reg_file[9065] <= 8'h00
            reg_file[9066] <= 8'h00
            reg_file[9067] <= 8'h00
            reg_file[9068] <= 8'h00
            reg_file[9069] <= 8'h00
            reg_file[9070] <= 8'h00
            reg_file[9071] <= 8'h00
            reg_file[9072] <= 8'h00
            reg_file[9073] <= 8'h00
            reg_file[9074] <= 8'h00
            reg_file[9075] <= 8'h00
            reg_file[9076] <= 8'h00
            reg_file[9077] <= 8'h00
            reg_file[9078] <= 8'h00
            reg_file[9079] <= 8'h00
            reg_file[9080] <= 8'h00
            reg_file[9081] <= 8'h00
            reg_file[9082] <= 8'h00
            reg_file[9083] <= 8'h00
            reg_file[9084] <= 8'h00
            reg_file[9085] <= 8'h00
            reg_file[9086] <= 8'h00
            reg_file[9087] <= 8'h00
            reg_file[9088] <= 8'h00
            reg_file[9089] <= 8'h00
            reg_file[9090] <= 8'h00
            reg_file[9091] <= 8'h00
            reg_file[9092] <= 8'h00
            reg_file[9093] <= 8'h00
            reg_file[9094] <= 8'h00
            reg_file[9095] <= 8'h00
            reg_file[9096] <= 8'h00
            reg_file[9097] <= 8'h00
            reg_file[9098] <= 8'h00
            reg_file[9099] <= 8'h00
            reg_file[9100] <= 8'h00
            reg_file[9101] <= 8'h00
            reg_file[9102] <= 8'h00
            reg_file[9103] <= 8'h00
            reg_file[9104] <= 8'h00
            reg_file[9105] <= 8'h00
            reg_file[9106] <= 8'h00
            reg_file[9107] <= 8'h00
            reg_file[9108] <= 8'h00
            reg_file[9109] <= 8'h00
            reg_file[9110] <= 8'h00
            reg_file[9111] <= 8'h00
            reg_file[9112] <= 8'h00
            reg_file[9113] <= 8'h00
            reg_file[9114] <= 8'h00
            reg_file[9115] <= 8'h00
            reg_file[9116] <= 8'h00
            reg_file[9117] <= 8'h00
            reg_file[9118] <= 8'h00
            reg_file[9119] <= 8'h00
            reg_file[9120] <= 8'h00
            reg_file[9121] <= 8'h00
            reg_file[9122] <= 8'h00
            reg_file[9123] <= 8'h00
            reg_file[9124] <= 8'h00
            reg_file[9125] <= 8'h00
            reg_file[9126] <= 8'h00
            reg_file[9127] <= 8'h00
            reg_file[9128] <= 8'h00
            reg_file[9129] <= 8'h00
            reg_file[9130] <= 8'h00
            reg_file[9131] <= 8'h00
            reg_file[9132] <= 8'h00
            reg_file[9133] <= 8'h00
            reg_file[9134] <= 8'h00
            reg_file[9135] <= 8'h00
            reg_file[9136] <= 8'h00
            reg_file[9137] <= 8'h00
            reg_file[9138] <= 8'h00
            reg_file[9139] <= 8'h00
            reg_file[9140] <= 8'h00
            reg_file[9141] <= 8'h00
            reg_file[9142] <= 8'h00
            reg_file[9143] <= 8'h00
            reg_file[9144] <= 8'h00
            reg_file[9145] <= 8'h00
            reg_file[9146] <= 8'h00
            reg_file[9147] <= 8'h00
            reg_file[9148] <= 8'h00
            reg_file[9149] <= 8'h00
            reg_file[9150] <= 8'h00
            reg_file[9151] <= 8'h00
            reg_file[9152] <= 8'h00
            reg_file[9153] <= 8'h00
            reg_file[9154] <= 8'h00
            reg_file[9155] <= 8'h00
            reg_file[9156] <= 8'h00
            reg_file[9157] <= 8'h00
            reg_file[9158] <= 8'h00
            reg_file[9159] <= 8'h00
            reg_file[9160] <= 8'h00
            reg_file[9161] <= 8'h00
            reg_file[9162] <= 8'h00
            reg_file[9163] <= 8'h00
            reg_file[9164] <= 8'h00
            reg_file[9165] <= 8'h00
            reg_file[9166] <= 8'h00
            reg_file[9167] <= 8'h00
            reg_file[9168] <= 8'h00
            reg_file[9169] <= 8'h00
            reg_file[9170] <= 8'h00
            reg_file[9171] <= 8'h00
            reg_file[9172] <= 8'h00
            reg_file[9173] <= 8'h00
            reg_file[9174] <= 8'h00
            reg_file[9175] <= 8'h00
            reg_file[9176] <= 8'h00
            reg_file[9177] <= 8'h00
            reg_file[9178] <= 8'h00
            reg_file[9179] <= 8'h00
            reg_file[9180] <= 8'h00
            reg_file[9181] <= 8'h00
            reg_file[9182] <= 8'h00
            reg_file[9183] <= 8'h00
            reg_file[9184] <= 8'h00
            reg_file[9185] <= 8'h00
            reg_file[9186] <= 8'h00
            reg_file[9187] <= 8'h00
            reg_file[9188] <= 8'h00
            reg_file[9189] <= 8'h00
            reg_file[9190] <= 8'h00
            reg_file[9191] <= 8'h00
            reg_file[9192] <= 8'h00
            reg_file[9193] <= 8'h00
            reg_file[9194] <= 8'h00
            reg_file[9195] <= 8'h00
            reg_file[9196] <= 8'h00
            reg_file[9197] <= 8'h00
            reg_file[9198] <= 8'h00
            reg_file[9199] <= 8'h00
            reg_file[9200] <= 8'h00
            reg_file[9201] <= 8'h00
            reg_file[9202] <= 8'h00
            reg_file[9203] <= 8'h00
            reg_file[9204] <= 8'h00
            reg_file[9205] <= 8'h00
            reg_file[9206] <= 8'h00
            reg_file[9207] <= 8'h00
            reg_file[9208] <= 8'h00
            reg_file[9209] <= 8'h00
            reg_file[9210] <= 8'h00
            reg_file[9211] <= 8'h00
            reg_file[9212] <= 8'h00
            reg_file[9213] <= 8'h00
            reg_file[9214] <= 8'h00
            reg_file[9215] <= 8'h00
            reg_file[9216] <= 8'h00
            reg_file[9217] <= 8'h00
            reg_file[9218] <= 8'h00
            reg_file[9219] <= 8'h00
            reg_file[9220] <= 8'h00
            reg_file[9221] <= 8'h00
            reg_file[9222] <= 8'h00
            reg_file[9223] <= 8'h00
            reg_file[9224] <= 8'h00
            reg_file[9225] <= 8'h00
            reg_file[9226] <= 8'h00
            reg_file[9227] <= 8'h00
            reg_file[9228] <= 8'h00
            reg_file[9229] <= 8'h00
            reg_file[9230] <= 8'h00
            reg_file[9231] <= 8'h00
            reg_file[9232] <= 8'h00
            reg_file[9233] <= 8'h00
            reg_file[9234] <= 8'h00
            reg_file[9235] <= 8'h00
            reg_file[9236] <= 8'h00
            reg_file[9237] <= 8'h00
            reg_file[9238] <= 8'h00
            reg_file[9239] <= 8'h00
            reg_file[9240] <= 8'h00
            reg_file[9241] <= 8'h00
            reg_file[9242] <= 8'h00
            reg_file[9243] <= 8'h00
            reg_file[9244] <= 8'h00
            reg_file[9245] <= 8'h00
            reg_file[9246] <= 8'h00
            reg_file[9247] <= 8'h00
            reg_file[9248] <= 8'h00
            reg_file[9249] <= 8'h00
            reg_file[9250] <= 8'h00
            reg_file[9251] <= 8'h00
            reg_file[9252] <= 8'h00
            reg_file[9253] <= 8'h00
            reg_file[9254] <= 8'h00
            reg_file[9255] <= 8'h00
            reg_file[9256] <= 8'h00
            reg_file[9257] <= 8'h00
            reg_file[9258] <= 8'h00
            reg_file[9259] <= 8'h00
            reg_file[9260] <= 8'h00
            reg_file[9261] <= 8'h00
            reg_file[9262] <= 8'h00
            reg_file[9263] <= 8'h00
            reg_file[9264] <= 8'h00
            reg_file[9265] <= 8'h00
            reg_file[9266] <= 8'h00
            reg_file[9267] <= 8'h00
            reg_file[9268] <= 8'h00
            reg_file[9269] <= 8'h00
            reg_file[9270] <= 8'h00
            reg_file[9271] <= 8'h00
            reg_file[9272] <= 8'h00
            reg_file[9273] <= 8'h00
            reg_file[9274] <= 8'h00
            reg_file[9275] <= 8'h00
            reg_file[9276] <= 8'h00
            reg_file[9277] <= 8'h00
            reg_file[9278] <= 8'h00
            reg_file[9279] <= 8'h00
            reg_file[9280] <= 8'h00
            reg_file[9281] <= 8'h00
            reg_file[9282] <= 8'h00
            reg_file[9283] <= 8'h00
            reg_file[9284] <= 8'h00
            reg_file[9285] <= 8'h00
            reg_file[9286] <= 8'h00
            reg_file[9287] <= 8'h00
            reg_file[9288] <= 8'h00
            reg_file[9289] <= 8'h00
            reg_file[9290] <= 8'h00
            reg_file[9291] <= 8'h00
            reg_file[9292] <= 8'h00
            reg_file[9293] <= 8'h00
            reg_file[9294] <= 8'h00
            reg_file[9295] <= 8'h00
            reg_file[9296] <= 8'h00
            reg_file[9297] <= 8'h00
            reg_file[9298] <= 8'h00
            reg_file[9299] <= 8'h00
            reg_file[9300] <= 8'h00
            reg_file[9301] <= 8'h00
            reg_file[9302] <= 8'h00
            reg_file[9303] <= 8'h00
            reg_file[9304] <= 8'h00
            reg_file[9305] <= 8'h00
            reg_file[9306] <= 8'h00
            reg_file[9307] <= 8'h00
            reg_file[9308] <= 8'h00
            reg_file[9309] <= 8'h00
            reg_file[9310] <= 8'h00
            reg_file[9311] <= 8'h00
            reg_file[9312] <= 8'h00
            reg_file[9313] <= 8'h00
            reg_file[9314] <= 8'h00
            reg_file[9315] <= 8'h00
            reg_file[9316] <= 8'h00
            reg_file[9317] <= 8'h00
            reg_file[9318] <= 8'h00
            reg_file[9319] <= 8'h00
            reg_file[9320] <= 8'h00
            reg_file[9321] <= 8'h00
            reg_file[9322] <= 8'h00
            reg_file[9323] <= 8'h00
            reg_file[9324] <= 8'h00
            reg_file[9325] <= 8'h00
            reg_file[9326] <= 8'h00
            reg_file[9327] <= 8'h00
            reg_file[9328] <= 8'h00
            reg_file[9329] <= 8'h00
            reg_file[9330] <= 8'h00
            reg_file[9331] <= 8'h00
            reg_file[9332] <= 8'h00
            reg_file[9333] <= 8'h00
            reg_file[9334] <= 8'h00
            reg_file[9335] <= 8'h00
            reg_file[9336] <= 8'h00
            reg_file[9337] <= 8'h00
            reg_file[9338] <= 8'h00
            reg_file[9339] <= 8'h00
            reg_file[9340] <= 8'h00
            reg_file[9341] <= 8'h00
            reg_file[9342] <= 8'h00
            reg_file[9343] <= 8'h00
            reg_file[9344] <= 8'h00
            reg_file[9345] <= 8'h00
            reg_file[9346] <= 8'h00
            reg_file[9347] <= 8'h00
            reg_file[9348] <= 8'h00
            reg_file[9349] <= 8'h00
            reg_file[9350] <= 8'h00
            reg_file[9351] <= 8'h00
            reg_file[9352] <= 8'h00
            reg_file[9353] <= 8'h00
            reg_file[9354] <= 8'h00
            reg_file[9355] <= 8'h00
            reg_file[9356] <= 8'h00
            reg_file[9357] <= 8'h00
            reg_file[9358] <= 8'h00
            reg_file[9359] <= 8'h00
            reg_file[9360] <= 8'h00
            reg_file[9361] <= 8'h00
            reg_file[9362] <= 8'h00
            reg_file[9363] <= 8'h00
            reg_file[9364] <= 8'h00
            reg_file[9365] <= 8'h00
            reg_file[9366] <= 8'h00
            reg_file[9367] <= 8'h00
            reg_file[9368] <= 8'h00
            reg_file[9369] <= 8'h00
            reg_file[9370] <= 8'h00
            reg_file[9371] <= 8'h00
            reg_file[9372] <= 8'h00
            reg_file[9373] <= 8'h00
            reg_file[9374] <= 8'h00
            reg_file[9375] <= 8'h00
            reg_file[9376] <= 8'h00
            reg_file[9377] <= 8'h00
            reg_file[9378] <= 8'h00
            reg_file[9379] <= 8'h00
            reg_file[9380] <= 8'h00
            reg_file[9381] <= 8'h00
            reg_file[9382] <= 8'h00
            reg_file[9383] <= 8'h00
            reg_file[9384] <= 8'h00
            reg_file[9385] <= 8'h00
            reg_file[9386] <= 8'h00
            reg_file[9387] <= 8'h00
            reg_file[9388] <= 8'h00
            reg_file[9389] <= 8'h00
            reg_file[9390] <= 8'h00
            reg_file[9391] <= 8'h00
            reg_file[9392] <= 8'h00
            reg_file[9393] <= 8'h00
            reg_file[9394] <= 8'h00
            reg_file[9395] <= 8'h00
            reg_file[9396] <= 8'h00
            reg_file[9397] <= 8'h00
            reg_file[9398] <= 8'h00
            reg_file[9399] <= 8'h00
            reg_file[9400] <= 8'h00
            reg_file[9401] <= 8'h00
            reg_file[9402] <= 8'h00
            reg_file[9403] <= 8'h00
            reg_file[9404] <= 8'h00
            reg_file[9405] <= 8'h00
            reg_file[9406] <= 8'h00
            reg_file[9407] <= 8'h00
            reg_file[9408] <= 8'h00
            reg_file[9409] <= 8'h00
            reg_file[9410] <= 8'h00
            reg_file[9411] <= 8'h00
            reg_file[9412] <= 8'h00
            reg_file[9413] <= 8'h00
            reg_file[9414] <= 8'h00
            reg_file[9415] <= 8'h00
            reg_file[9416] <= 8'h00
            reg_file[9417] <= 8'h00
            reg_file[9418] <= 8'h00
            reg_file[9419] <= 8'h00
            reg_file[9420] <= 8'h00
            reg_file[9421] <= 8'h00
            reg_file[9422] <= 8'h00
            reg_file[9423] <= 8'h00
            reg_file[9424] <= 8'h00
            reg_file[9425] <= 8'h00
            reg_file[9426] <= 8'h00
            reg_file[9427] <= 8'h00
            reg_file[9428] <= 8'h00
            reg_file[9429] <= 8'h00
            reg_file[9430] <= 8'h00
            reg_file[9431] <= 8'h00
            reg_file[9432] <= 8'h00
            reg_file[9433] <= 8'h00
            reg_file[9434] <= 8'h00
            reg_file[9435] <= 8'h00
            reg_file[9436] <= 8'h00
            reg_file[9437] <= 8'h00
            reg_file[9438] <= 8'h00
            reg_file[9439] <= 8'h00
            reg_file[9440] <= 8'h00
            reg_file[9441] <= 8'h00
            reg_file[9442] <= 8'h00
            reg_file[9443] <= 8'h00
            reg_file[9444] <= 8'h00
            reg_file[9445] <= 8'h00
            reg_file[9446] <= 8'h00
            reg_file[9447] <= 8'h00
            reg_file[9448] <= 8'h00
            reg_file[9449] <= 8'h00
            reg_file[9450] <= 8'h00
            reg_file[9451] <= 8'h00
            reg_file[9452] <= 8'h00
            reg_file[9453] <= 8'h00
            reg_file[9454] <= 8'h00
            reg_file[9455] <= 8'h00
            reg_file[9456] <= 8'h00
            reg_file[9457] <= 8'h00
            reg_file[9458] <= 8'h00
            reg_file[9459] <= 8'h00
            reg_file[9460] <= 8'h00
            reg_file[9461] <= 8'h00
            reg_file[9462] <= 8'h00
            reg_file[9463] <= 8'h00
            reg_file[9464] <= 8'h00
            reg_file[9465] <= 8'h00
            reg_file[9466] <= 8'h00
            reg_file[9467] <= 8'h00
            reg_file[9468] <= 8'h00
            reg_file[9469] <= 8'h00
            reg_file[9470] <= 8'h00
            reg_file[9471] <= 8'h00
            reg_file[9472] <= 8'h00
            reg_file[9473] <= 8'h00
            reg_file[9474] <= 8'h00
            reg_file[9475] <= 8'h00
            reg_file[9476] <= 8'h00
            reg_file[9477] <= 8'h00
            reg_file[9478] <= 8'h00
            reg_file[9479] <= 8'h00
            reg_file[9480] <= 8'h00
            reg_file[9481] <= 8'h00
            reg_file[9482] <= 8'h00
            reg_file[9483] <= 8'h00
            reg_file[9484] <= 8'h00
            reg_file[9485] <= 8'h00
            reg_file[9486] <= 8'h00
            reg_file[9487] <= 8'h00
            reg_file[9488] <= 8'h00
            reg_file[9489] <= 8'h00
            reg_file[9490] <= 8'h00
            reg_file[9491] <= 8'h00
            reg_file[9492] <= 8'h00
            reg_file[9493] <= 8'h00
            reg_file[9494] <= 8'h00
            reg_file[9495] <= 8'h00
            reg_file[9496] <= 8'h00
            reg_file[9497] <= 8'h00
            reg_file[9498] <= 8'h00
            reg_file[9499] <= 8'h00
            reg_file[9500] <= 8'h00
            reg_file[9501] <= 8'h00
            reg_file[9502] <= 8'h00
            reg_file[9503] <= 8'h00
            reg_file[9504] <= 8'h00
            reg_file[9505] <= 8'h00
            reg_file[9506] <= 8'h00
            reg_file[9507] <= 8'h00
            reg_file[9508] <= 8'h00
            reg_file[9509] <= 8'h00
            reg_file[9510] <= 8'h00
            reg_file[9511] <= 8'h00
            reg_file[9512] <= 8'h00
            reg_file[9513] <= 8'h00
            reg_file[9514] <= 8'h00
            reg_file[9515] <= 8'h00
            reg_file[9516] <= 8'h00
            reg_file[9517] <= 8'h00
            reg_file[9518] <= 8'h00
            reg_file[9519] <= 8'h00
            reg_file[9520] <= 8'h00
            reg_file[9521] <= 8'h00
            reg_file[9522] <= 8'h00
            reg_file[9523] <= 8'h00
            reg_file[9524] <= 8'h00
            reg_file[9525] <= 8'h00
            reg_file[9526] <= 8'h00
            reg_file[9527] <= 8'h00
            reg_file[9528] <= 8'h00
            reg_file[9529] <= 8'h00
            reg_file[9530] <= 8'h00
            reg_file[9531] <= 8'h00
            reg_file[9532] <= 8'h00
            reg_file[9533] <= 8'h00
            reg_file[9534] <= 8'h00
            reg_file[9535] <= 8'h00
            reg_file[9536] <= 8'h00
            reg_file[9537] <= 8'h00
            reg_file[9538] <= 8'h00
            reg_file[9539] <= 8'h00
            reg_file[9540] <= 8'h00
            reg_file[9541] <= 8'h00
            reg_file[9542] <= 8'h00
            reg_file[9543] <= 8'h00
            reg_file[9544] <= 8'h00
            reg_file[9545] <= 8'h00
            reg_file[9546] <= 8'h00
            reg_file[9547] <= 8'h00
            reg_file[9548] <= 8'h00
            reg_file[9549] <= 8'h00
            reg_file[9550] <= 8'h00
            reg_file[9551] <= 8'h00
            reg_file[9552] <= 8'h00
            reg_file[9553] <= 8'h00
            reg_file[9554] <= 8'h00
            reg_file[9555] <= 8'h00
            reg_file[9556] <= 8'h00
            reg_file[9557] <= 8'h00
            reg_file[9558] <= 8'h00
            reg_file[9559] <= 8'h00
            reg_file[9560] <= 8'h00
            reg_file[9561] <= 8'h00
            reg_file[9562] <= 8'h00
            reg_file[9563] <= 8'h00
            reg_file[9564] <= 8'h00
            reg_file[9565] <= 8'h00
            reg_file[9566] <= 8'h00
            reg_file[9567] <= 8'h00
            reg_file[9568] <= 8'h00
            reg_file[9569] <= 8'h00
            reg_file[9570] <= 8'h00
            reg_file[9571] <= 8'h00
            reg_file[9572] <= 8'h00
            reg_file[9573] <= 8'h00
            reg_file[9574] <= 8'h00
            reg_file[9575] <= 8'h00
            reg_file[9576] <= 8'h00
            reg_file[9577] <= 8'h00
            reg_file[9578] <= 8'h00
            reg_file[9579] <= 8'h00
            reg_file[9580] <= 8'h00
            reg_file[9581] <= 8'h00
            reg_file[9582] <= 8'h00
            reg_file[9583] <= 8'h00
            reg_file[9584] <= 8'h00
            reg_file[9585] <= 8'h00
            reg_file[9586] <= 8'h00
            reg_file[9587] <= 8'h00
            reg_file[9588] <= 8'h00
            reg_file[9589] <= 8'h00
            reg_file[9590] <= 8'h00
            reg_file[9591] <= 8'h00
            reg_file[9592] <= 8'h00
            reg_file[9593] <= 8'h00
            reg_file[9594] <= 8'h00
            reg_file[9595] <= 8'h00
            reg_file[9596] <= 8'h00
            reg_file[9597] <= 8'h00
            reg_file[9598] <= 8'h00
            reg_file[9599] <= 8'h00
            reg_file[9600] <= 8'h00
            reg_file[9601] <= 8'h00
            reg_file[9602] <= 8'h00
            reg_file[9603] <= 8'h00
            reg_file[9604] <= 8'h00
            reg_file[9605] <= 8'h00
            reg_file[9606] <= 8'h00
            reg_file[9607] <= 8'h00
            reg_file[9608] <= 8'h00
            reg_file[9609] <= 8'h00
            reg_file[9610] <= 8'h00
            reg_file[9611] <= 8'h00
            reg_file[9612] <= 8'h00
            reg_file[9613] <= 8'h00
            reg_file[9614] <= 8'h00
            reg_file[9615] <= 8'h00
            reg_file[9616] <= 8'h00
            reg_file[9617] <= 8'h00
            reg_file[9618] <= 8'h00
            reg_file[9619] <= 8'h00
            reg_file[9620] <= 8'h00
            reg_file[9621] <= 8'h00
            reg_file[9622] <= 8'h00
            reg_file[9623] <= 8'h00
            reg_file[9624] <= 8'h00
            reg_file[9625] <= 8'h00
            reg_file[9626] <= 8'h00
            reg_file[9627] <= 8'h00
            reg_file[9628] <= 8'h00
            reg_file[9629] <= 8'h00
            reg_file[9630] <= 8'h00
            reg_file[9631] <= 8'h00
            reg_file[9632] <= 8'h00
            reg_file[9633] <= 8'h00
            reg_file[9634] <= 8'h00
            reg_file[9635] <= 8'h00
            reg_file[9636] <= 8'h00
            reg_file[9637] <= 8'h00
            reg_file[9638] <= 8'h00
            reg_file[9639] <= 8'h00
            reg_file[9640] <= 8'h00
            reg_file[9641] <= 8'h00
            reg_file[9642] <= 8'h00
            reg_file[9643] <= 8'h00
            reg_file[9644] <= 8'h00
            reg_file[9645] <= 8'h00
            reg_file[9646] <= 8'h00
            reg_file[9647] <= 8'h00
            reg_file[9648] <= 8'h00
            reg_file[9649] <= 8'h00
            reg_file[9650] <= 8'h00
            reg_file[9651] <= 8'h00
            reg_file[9652] <= 8'h00
            reg_file[9653] <= 8'h00
            reg_file[9654] <= 8'h00
            reg_file[9655] <= 8'h00
            reg_file[9656] <= 8'h00
            reg_file[9657] <= 8'h00
            reg_file[9658] <= 8'h00
            reg_file[9659] <= 8'h00
            reg_file[9660] <= 8'h00
            reg_file[9661] <= 8'h00
            reg_file[9662] <= 8'h00
            reg_file[9663] <= 8'h00
            reg_file[9664] <= 8'h00
            reg_file[9665] <= 8'h00
            reg_file[9666] <= 8'h00
            reg_file[9667] <= 8'h00
            reg_file[9668] <= 8'h00
            reg_file[9669] <= 8'h00
            reg_file[9670] <= 8'h00
            reg_file[9671] <= 8'h00
            reg_file[9672] <= 8'h00
            reg_file[9673] <= 8'h00
            reg_file[9674] <= 8'h00
            reg_file[9675] <= 8'h00
            reg_file[9676] <= 8'h00
            reg_file[9677] <= 8'h00
            reg_file[9678] <= 8'h00
            reg_file[9679] <= 8'h00
            reg_file[9680] <= 8'h00
            reg_file[9681] <= 8'h00
            reg_file[9682] <= 8'h00
            reg_file[9683] <= 8'h00
            reg_file[9684] <= 8'h00
            reg_file[9685] <= 8'h00
            reg_file[9686] <= 8'h00
            reg_file[9687] <= 8'h00
            reg_file[9688] <= 8'h00
            reg_file[9689] <= 8'h00
            reg_file[9690] <= 8'h00
            reg_file[9691] <= 8'h00
            reg_file[9692] <= 8'h00
            reg_file[9693] <= 8'h00
            reg_file[9694] <= 8'h00
            reg_file[9695] <= 8'h00
            reg_file[9696] <= 8'h00
            reg_file[9697] <= 8'h00
            reg_file[9698] <= 8'h00
            reg_file[9699] <= 8'h00
            reg_file[9700] <= 8'h00
            reg_file[9701] <= 8'h00
            reg_file[9702] <= 8'h00
            reg_file[9703] <= 8'h00
            reg_file[9704] <= 8'h00
            reg_file[9705] <= 8'h00
            reg_file[9706] <= 8'h00
            reg_file[9707] <= 8'h00
            reg_file[9708] <= 8'h00
            reg_file[9709] <= 8'h00
            reg_file[9710] <= 8'h00
            reg_file[9711] <= 8'h00
            reg_file[9712] <= 8'h00
            reg_file[9713] <= 8'h00
            reg_file[9714] <= 8'h00
            reg_file[9715] <= 8'h00
            reg_file[9716] <= 8'h00
            reg_file[9717] <= 8'h00
            reg_file[9718] <= 8'h00
            reg_file[9719] <= 8'h00
            reg_file[9720] <= 8'h00
            reg_file[9721] <= 8'h00
            reg_file[9722] <= 8'h00
            reg_file[9723] <= 8'h00
            reg_file[9724] <= 8'h00
            reg_file[9725] <= 8'h00
            reg_file[9726] <= 8'h00
            reg_file[9727] <= 8'h00
            reg_file[9728] <= 8'h00
            reg_file[9729] <= 8'h00
            reg_file[9730] <= 8'h00
            reg_file[9731] <= 8'h00
            reg_file[9732] <= 8'h00
            reg_file[9733] <= 8'h00
            reg_file[9734] <= 8'h00
            reg_file[9735] <= 8'h00
            reg_file[9736] <= 8'h00
            reg_file[9737] <= 8'h00
            reg_file[9738] <= 8'h00
            reg_file[9739] <= 8'h00
            reg_file[9740] <= 8'h00
            reg_file[9741] <= 8'h00
            reg_file[9742] <= 8'h00
            reg_file[9743] <= 8'h00
            reg_file[9744] <= 8'h00
            reg_file[9745] <= 8'h00
            reg_file[9746] <= 8'h00
            reg_file[9747] <= 8'h00
            reg_file[9748] <= 8'h00
            reg_file[9749] <= 8'h00
            reg_file[9750] <= 8'h00
            reg_file[9751] <= 8'h00
            reg_file[9752] <= 8'h00
            reg_file[9753] <= 8'h00
            reg_file[9754] <= 8'h00
            reg_file[9755] <= 8'h00
            reg_file[9756] <= 8'h00
            reg_file[9757] <= 8'h00
            reg_file[9758] <= 8'h00
            reg_file[9759] <= 8'h00
            reg_file[9760] <= 8'h00
            reg_file[9761] <= 8'h00
            reg_file[9762] <= 8'h00
            reg_file[9763] <= 8'h00
            reg_file[9764] <= 8'h00
            reg_file[9765] <= 8'h00
            reg_file[9766] <= 8'h00
            reg_file[9767] <= 8'h00
            reg_file[9768] <= 8'h00
            reg_file[9769] <= 8'h00
            reg_file[9770] <= 8'h00
            reg_file[9771] <= 8'h00
            reg_file[9772] <= 8'h00
            reg_file[9773] <= 8'h00
            reg_file[9774] <= 8'h00
            reg_file[9775] <= 8'h00
            reg_file[9776] <= 8'h00
            reg_file[9777] <= 8'h00
            reg_file[9778] <= 8'h00
            reg_file[9779] <= 8'h00
            reg_file[9780] <= 8'h00
            reg_file[9781] <= 8'h00
            reg_file[9782] <= 8'h00
            reg_file[9783] <= 8'h00
            reg_file[9784] <= 8'h00
            reg_file[9785] <= 8'h00
            reg_file[9786] <= 8'h00
            reg_file[9787] <= 8'h00
            reg_file[9788] <= 8'h00
            reg_file[9789] <= 8'h00
            reg_file[9790] <= 8'h00
            reg_file[9791] <= 8'h00
            reg_file[9792] <= 8'h00
            reg_file[9793] <= 8'h00
            reg_file[9794] <= 8'h00
            reg_file[9795] <= 8'h00
            reg_file[9796] <= 8'h00
            reg_file[9797] <= 8'h00
            reg_file[9798] <= 8'h00
            reg_file[9799] <= 8'h00
            reg_file[9800] <= 8'h00
            reg_file[9801] <= 8'h00
            reg_file[9802] <= 8'h00
            reg_file[9803] <= 8'h00
            reg_file[9804] <= 8'h00
            reg_file[9805] <= 8'h00
            reg_file[9806] <= 8'h00
            reg_file[9807] <= 8'h00
            reg_file[9808] <= 8'h00
            reg_file[9809] <= 8'h00
            reg_file[9810] <= 8'h00
            reg_file[9811] <= 8'h00
            reg_file[9812] <= 8'h00
            reg_file[9813] <= 8'h00
            reg_file[9814] <= 8'h00
            reg_file[9815] <= 8'h00
            reg_file[9816] <= 8'h00
            reg_file[9817] <= 8'h00
            reg_file[9818] <= 8'h00
            reg_file[9819] <= 8'h00
            reg_file[9820] <= 8'h00
            reg_file[9821] <= 8'h00
            reg_file[9822] <= 8'h00
            reg_file[9823] <= 8'h00
            reg_file[9824] <= 8'h00
            reg_file[9825] <= 8'h00
            reg_file[9826] <= 8'h00
            reg_file[9827] <= 8'h00
            reg_file[9828] <= 8'h00
            reg_file[9829] <= 8'h00
            reg_file[9830] <= 8'h00
            reg_file[9831] <= 8'h00
            reg_file[9832] <= 8'h00
            reg_file[9833] <= 8'h00
            reg_file[9834] <= 8'h00
            reg_file[9835] <= 8'h00
            reg_file[9836] <= 8'h00
            reg_file[9837] <= 8'h00
            reg_file[9838] <= 8'h00
            reg_file[9839] <= 8'h00
            reg_file[9840] <= 8'h00
            reg_file[9841] <= 8'h00
            reg_file[9842] <= 8'h00
            reg_file[9843] <= 8'h00
            reg_file[9844] <= 8'h00
            reg_file[9845] <= 8'h00
            reg_file[9846] <= 8'h00
            reg_file[9847] <= 8'h00
            reg_file[9848] <= 8'h00
            reg_file[9849] <= 8'h00
            reg_file[9850] <= 8'h00
            reg_file[9851] <= 8'h00
            reg_file[9852] <= 8'h00
            reg_file[9853] <= 8'h00
            reg_file[9854] <= 8'h00
            reg_file[9855] <= 8'h00
            reg_file[9856] <= 8'h00
            reg_file[9857] <= 8'h00
            reg_file[9858] <= 8'h00
            reg_file[9859] <= 8'h00
            reg_file[9860] <= 8'h00
            reg_file[9861] <= 8'h00
            reg_file[9862] <= 8'h00
            reg_file[9863] <= 8'h00
            reg_file[9864] <= 8'h00
            reg_file[9865] <= 8'h00
            reg_file[9866] <= 8'h00
            reg_file[9867] <= 8'h00
            reg_file[9868] <= 8'h00
            reg_file[9869] <= 8'h00
            reg_file[9870] <= 8'h00
            reg_file[9871] <= 8'h00
            reg_file[9872] <= 8'h00
            reg_file[9873] <= 8'h00
            reg_file[9874] <= 8'h00
            reg_file[9875] <= 8'h00
            reg_file[9876] <= 8'h00
            reg_file[9877] <= 8'h00
            reg_file[9878] <= 8'h00
            reg_file[9879] <= 8'h00
            reg_file[9880] <= 8'h00
            reg_file[9881] <= 8'h00
            reg_file[9882] <= 8'h00
            reg_file[9883] <= 8'h00
            reg_file[9884] <= 8'h00
            reg_file[9885] <= 8'h00
            reg_file[9886] <= 8'h00
            reg_file[9887] <= 8'h00
            reg_file[9888] <= 8'h00
            reg_file[9889] <= 8'h00
            reg_file[9890] <= 8'h00
            reg_file[9891] <= 8'h00
            reg_file[9892] <= 8'h00
            reg_file[9893] <= 8'h00
            reg_file[9894] <= 8'h00
            reg_file[9895] <= 8'h00
            reg_file[9896] <= 8'h00
            reg_file[9897] <= 8'h00
            reg_file[9898] <= 8'h00
            reg_file[9899] <= 8'h00
            reg_file[9900] <= 8'h00
            reg_file[9901] <= 8'h00
            reg_file[9902] <= 8'h00
            reg_file[9903] <= 8'h00
            reg_file[9904] <= 8'h00
            reg_file[9905] <= 8'h00
            reg_file[9906] <= 8'h00
            reg_file[9907] <= 8'h00
            reg_file[9908] <= 8'h00
            reg_file[9909] <= 8'h00
            reg_file[9910] <= 8'h00
            reg_file[9911] <= 8'h00
            reg_file[9912] <= 8'h00
            reg_file[9913] <= 8'h00
            reg_file[9914] <= 8'h00
            reg_file[9915] <= 8'h00
            reg_file[9916] <= 8'h00
            reg_file[9917] <= 8'h00
            reg_file[9918] <= 8'h00
            reg_file[9919] <= 8'h00
            reg_file[9920] <= 8'h00
            reg_file[9921] <= 8'h00
            reg_file[9922] <= 8'h00
            reg_file[9923] <= 8'h00
            reg_file[9924] <= 8'h00
            reg_file[9925] <= 8'h00
            reg_file[9926] <= 8'h00
            reg_file[9927] <= 8'h00
            reg_file[9928] <= 8'h00
            reg_file[9929] <= 8'h00
            reg_file[9930] <= 8'h00
            reg_file[9931] <= 8'h00
            reg_file[9932] <= 8'h00
            reg_file[9933] <= 8'h00
            reg_file[9934] <= 8'h00
            reg_file[9935] <= 8'h00
            reg_file[9936] <= 8'h00
            reg_file[9937] <= 8'h00
            reg_file[9938] <= 8'h00
            reg_file[9939] <= 8'h00
            reg_file[9940] <= 8'h00
            reg_file[9941] <= 8'h00
            reg_file[9942] <= 8'h00
            reg_file[9943] <= 8'h00
            reg_file[9944] <= 8'h00
            reg_file[9945] <= 8'h00
            reg_file[9946] <= 8'h00
            reg_file[9947] <= 8'h00
            reg_file[9948] <= 8'h00
            reg_file[9949] <= 8'h00
            reg_file[9950] <= 8'h00
            reg_file[9951] <= 8'h00
            reg_file[9952] <= 8'h00
            reg_file[9953] <= 8'h00
            reg_file[9954] <= 8'h00
            reg_file[9955] <= 8'h00
            reg_file[9956] <= 8'h00
            reg_file[9957] <= 8'h00
            reg_file[9958] <= 8'h00
            reg_file[9959] <= 8'h00
            reg_file[9960] <= 8'h00
            reg_file[9961] <= 8'h00
            reg_file[9962] <= 8'h00
            reg_file[9963] <= 8'h00
            reg_file[9964] <= 8'h00
            reg_file[9965] <= 8'h00
            reg_file[9966] <= 8'h00
            reg_file[9967] <= 8'h00
            reg_file[9968] <= 8'h00
            reg_file[9969] <= 8'h00
            reg_file[9970] <= 8'h00
            reg_file[9971] <= 8'h00
            reg_file[9972] <= 8'h00
            reg_file[9973] <= 8'h00
            reg_file[9974] <= 8'h00
            reg_file[9975] <= 8'h00
            reg_file[9976] <= 8'h00
            reg_file[9977] <= 8'h00
            reg_file[9978] <= 8'h00
            reg_file[9979] <= 8'h00
            reg_file[9980] <= 8'h00
            reg_file[9981] <= 8'h00
            reg_file[9982] <= 8'h00
            reg_file[9983] <= 8'h00
            reg_file[9984] <= 8'h00
            reg_file[9985] <= 8'h00
            reg_file[9986] <= 8'h00
            reg_file[9987] <= 8'h00
            reg_file[9988] <= 8'h00
            reg_file[9989] <= 8'h00
            reg_file[9990] <= 8'h00
            reg_file[9991] <= 8'h00
            reg_file[9992] <= 8'h00
            reg_file[9993] <= 8'h00
            reg_file[9994] <= 8'h00
            reg_file[9995] <= 8'h00
            reg_file[9996] <= 8'h00
            reg_file[9997] <= 8'h00
            reg_file[9998] <= 8'h00
            reg_file[9999] <= 8'h00
            reg_file[10000] <= 8'h00
            reg_file[10001] <= 8'h00
            reg_file[10002] <= 8'h00
            reg_file[10003] <= 8'h00
            reg_file[10004] <= 8'h00
            reg_file[10005] <= 8'h00
            reg_file[10006] <= 8'h00
            reg_file[10007] <= 8'h00
            reg_file[10008] <= 8'h00
            reg_file[10009] <= 8'h00
            reg_file[10010] <= 8'h00
            reg_file[10011] <= 8'h00
            reg_file[10012] <= 8'h00
            reg_file[10013] <= 8'h00
            reg_file[10014] <= 8'h00
            reg_file[10015] <= 8'h00
            reg_file[10016] <= 8'h00
            reg_file[10017] <= 8'h00
            reg_file[10018] <= 8'h00
            reg_file[10019] <= 8'h00
            reg_file[10020] <= 8'h00
            reg_file[10021] <= 8'h00
            reg_file[10022] <= 8'h00
            reg_file[10023] <= 8'h00
            reg_file[10024] <= 8'h00
            reg_file[10025] <= 8'h00
            reg_file[10026] <= 8'h00
            reg_file[10027] <= 8'h00
            reg_file[10028] <= 8'h00
            reg_file[10029] <= 8'h00
            reg_file[10030] <= 8'h00
            reg_file[10031] <= 8'h00
            reg_file[10032] <= 8'h00
            reg_file[10033] <= 8'h00
            reg_file[10034] <= 8'h00
            reg_file[10035] <= 8'h00
            reg_file[10036] <= 8'h00
            reg_file[10037] <= 8'h00
            reg_file[10038] <= 8'h00
            reg_file[10039] <= 8'h00
            reg_file[10040] <= 8'h00
            reg_file[10041] <= 8'h00
            reg_file[10042] <= 8'h00
            reg_file[10043] <= 8'h00
            reg_file[10044] <= 8'h00
            reg_file[10045] <= 8'h00
            reg_file[10046] <= 8'h00
            reg_file[10047] <= 8'h00
            reg_file[10048] <= 8'h00
            reg_file[10049] <= 8'h00
            reg_file[10050] <= 8'h00
            reg_file[10051] <= 8'h00
            reg_file[10052] <= 8'h00
            reg_file[10053] <= 8'h00
            reg_file[10054] <= 8'h00
            reg_file[10055] <= 8'h00
            reg_file[10056] <= 8'h00
            reg_file[10057] <= 8'h00
            reg_file[10058] <= 8'h00
            reg_file[10059] <= 8'h00
            reg_file[10060] <= 8'h00
            reg_file[10061] <= 8'h00
            reg_file[10062] <= 8'h00
            reg_file[10063] <= 8'h00
            reg_file[10064] <= 8'h00
            reg_file[10065] <= 8'h00
            reg_file[10066] <= 8'h00
            reg_file[10067] <= 8'h00
            reg_file[10068] <= 8'h00
            reg_file[10069] <= 8'h00
            reg_file[10070] <= 8'h00
            reg_file[10071] <= 8'h00
            reg_file[10072] <= 8'h00
            reg_file[10073] <= 8'h00
            reg_file[10074] <= 8'h00
            reg_file[10075] <= 8'h00
            reg_file[10076] <= 8'h00
            reg_file[10077] <= 8'h00
            reg_file[10078] <= 8'h00
            reg_file[10079] <= 8'h00
            reg_file[10080] <= 8'h00
            reg_file[10081] <= 8'h00
            reg_file[10082] <= 8'h00
            reg_file[10083] <= 8'h00
            reg_file[10084] <= 8'h00
            reg_file[10085] <= 8'h00
            reg_file[10086] <= 8'h00
            reg_file[10087] <= 8'h00
            reg_file[10088] <= 8'h00
            reg_file[10089] <= 8'h00
            reg_file[10090] <= 8'h00
            reg_file[10091] <= 8'h00
            reg_file[10092] <= 8'h00
            reg_file[10093] <= 8'h00
            reg_file[10094] <= 8'h00
            reg_file[10095] <= 8'h00
            reg_file[10096] <= 8'h00
            reg_file[10097] <= 8'h00
            reg_file[10098] <= 8'h00
            reg_file[10099] <= 8'h00
            reg_file[10100] <= 8'h00
            reg_file[10101] <= 8'h00
            reg_file[10102] <= 8'h00
            reg_file[10103] <= 8'h00
            reg_file[10104] <= 8'h00
            reg_file[10105] <= 8'h00
            reg_file[10106] <= 8'h00
            reg_file[10107] <= 8'h00
            reg_file[10108] <= 8'h00
            reg_file[10109] <= 8'h00
            reg_file[10110] <= 8'h00
            reg_file[10111] <= 8'h00
            reg_file[10112] <= 8'h00
            reg_file[10113] <= 8'h00
            reg_file[10114] <= 8'h00
            reg_file[10115] <= 8'h00
            reg_file[10116] <= 8'h00
            reg_file[10117] <= 8'h00
            reg_file[10118] <= 8'h00
            reg_file[10119] <= 8'h00
            reg_file[10120] <= 8'h00
            reg_file[10121] <= 8'h00
            reg_file[10122] <= 8'h00
            reg_file[10123] <= 8'h00
            reg_file[10124] <= 8'h00
            reg_file[10125] <= 8'h00
            reg_file[10126] <= 8'h00
            reg_file[10127] <= 8'h00
            reg_file[10128] <= 8'h00
            reg_file[10129] <= 8'h00
            reg_file[10130] <= 8'h00
            reg_file[10131] <= 8'h00
            reg_file[10132] <= 8'h00
            reg_file[10133] <= 8'h00
            reg_file[10134] <= 8'h00
            reg_file[10135] <= 8'h00
            reg_file[10136] <= 8'h00
            reg_file[10137] <= 8'h00
            reg_file[10138] <= 8'h00
            reg_file[10139] <= 8'h00
            reg_file[10140] <= 8'h00
            reg_file[10141] <= 8'h00
            reg_file[10142] <= 8'h00
            reg_file[10143] <= 8'h00
            reg_file[10144] <= 8'h00
            reg_file[10145] <= 8'h00
            reg_file[10146] <= 8'h00
            reg_file[10147] <= 8'h00
            reg_file[10148] <= 8'h00
            reg_file[10149] <= 8'h00
            reg_file[10150] <= 8'h00
            reg_file[10151] <= 8'h00
            reg_file[10152] <= 8'h00
            reg_file[10153] <= 8'h00
            reg_file[10154] <= 8'h00
            reg_file[10155] <= 8'h00
            reg_file[10156] <= 8'h00
            reg_file[10157] <= 8'h00
            reg_file[10158] <= 8'h00
            reg_file[10159] <= 8'h00
            reg_file[10160] <= 8'h00
            reg_file[10161] <= 8'h00
            reg_file[10162] <= 8'h00
            reg_file[10163] <= 8'h00
            reg_file[10164] <= 8'h00
            reg_file[10165] <= 8'h00
            reg_file[10166] <= 8'h00
            reg_file[10167] <= 8'h00
            reg_file[10168] <= 8'h00
            reg_file[10169] <= 8'h00
            reg_file[10170] <= 8'h00
            reg_file[10171] <= 8'h00
            reg_file[10172] <= 8'h00
            reg_file[10173] <= 8'h00
            reg_file[10174] <= 8'h00
            reg_file[10175] <= 8'h00
            reg_file[10176] <= 8'h00
            reg_file[10177] <= 8'h00
            reg_file[10178] <= 8'h00
            reg_file[10179] <= 8'h00
            reg_file[10180] <= 8'h00
            reg_file[10181] <= 8'h00
            reg_file[10182] <= 8'h00
            reg_file[10183] <= 8'h00
            reg_file[10184] <= 8'h00
            reg_file[10185] <= 8'h00
            reg_file[10186] <= 8'h00
            reg_file[10187] <= 8'h00
            reg_file[10188] <= 8'h00
            reg_file[10189] <= 8'h00
            reg_file[10190] <= 8'h00
            reg_file[10191] <= 8'h00
            reg_file[10192] <= 8'h00
            reg_file[10193] <= 8'h00
            reg_file[10194] <= 8'h00
            reg_file[10195] <= 8'h00
            reg_file[10196] <= 8'h00
            reg_file[10197] <= 8'h00
            reg_file[10198] <= 8'h00
            reg_file[10199] <= 8'h00
            reg_file[10200] <= 8'h00
            reg_file[10201] <= 8'h00
            reg_file[10202] <= 8'h00
            reg_file[10203] <= 8'h00
            reg_file[10204] <= 8'h00
            reg_file[10205] <= 8'h00
            reg_file[10206] <= 8'h00
            reg_file[10207] <= 8'h00
            reg_file[10208] <= 8'h00
            reg_file[10209] <= 8'h00
            reg_file[10210] <= 8'h00
            reg_file[10211] <= 8'h00
            reg_file[10212] <= 8'h00
            reg_file[10213] <= 8'h00
            reg_file[10214] <= 8'h00
            reg_file[10215] <= 8'h00
            reg_file[10216] <= 8'h00
            reg_file[10217] <= 8'h00
            reg_file[10218] <= 8'h00
            reg_file[10219] <= 8'h00
            reg_file[10220] <= 8'h00
            reg_file[10221] <= 8'h00
            reg_file[10222] <= 8'h00
            reg_file[10223] <= 8'h00
            reg_file[10224] <= 8'h00
            reg_file[10225] <= 8'h00
            reg_file[10226] <= 8'h00
            reg_file[10227] <= 8'h00
            reg_file[10228] <= 8'h00
            reg_file[10229] <= 8'h00
            reg_file[10230] <= 8'h00
            reg_file[10231] <= 8'h00
            reg_file[10232] <= 8'h00
            reg_file[10233] <= 8'h00
            reg_file[10234] <= 8'h00
            reg_file[10235] <= 8'h00
            reg_file[10236] <= 8'h00
            reg_file[10237] <= 8'h00
            reg_file[10238] <= 8'h00
            reg_file[10239] <= 8'h00
            reg_file[10240] <= 8'h00
            reg_file[10241] <= 8'h00
            reg_file[10242] <= 8'h00
            reg_file[10243] <= 8'h00
            reg_file[10244] <= 8'h00
            reg_file[10245] <= 8'h00
            reg_file[10246] <= 8'h00
            reg_file[10247] <= 8'h00
            reg_file[10248] <= 8'h00
            reg_file[10249] <= 8'h00
            reg_file[10250] <= 8'h00
            reg_file[10251] <= 8'h00
            reg_file[10252] <= 8'h00
            reg_file[10253] <= 8'h00
            reg_file[10254] <= 8'h00
            reg_file[10255] <= 8'h00
            reg_file[10256] <= 8'h00
            reg_file[10257] <= 8'h00
            reg_file[10258] <= 8'h00
            reg_file[10259] <= 8'h00
            reg_file[10260] <= 8'h00
            reg_file[10261] <= 8'h00
            reg_file[10262] <= 8'h00
            reg_file[10263] <= 8'h00
            reg_file[10264] <= 8'h00
            reg_file[10265] <= 8'h00
            reg_file[10266] <= 8'h00
            reg_file[10267] <= 8'h00
            reg_file[10268] <= 8'h00
            reg_file[10269] <= 8'h00
            reg_file[10270] <= 8'h00
            reg_file[10271] <= 8'h00
            reg_file[10272] <= 8'h00
            reg_file[10273] <= 8'h00
            reg_file[10274] <= 8'h00
            reg_file[10275] <= 8'h00
            reg_file[10276] <= 8'h00
            reg_file[10277] <= 8'h00
            reg_file[10278] <= 8'h00
            reg_file[10279] <= 8'h00
            reg_file[10280] <= 8'h00
            reg_file[10281] <= 8'h00
            reg_file[10282] <= 8'h00
            reg_file[10283] <= 8'h00
            reg_file[10284] <= 8'h00
            reg_file[10285] <= 8'h00
            reg_file[10286] <= 8'h00
            reg_file[10287] <= 8'h00
            reg_file[10288] <= 8'h00
            reg_file[10289] <= 8'h00
            reg_file[10290] <= 8'h00
            reg_file[10291] <= 8'h00
            reg_file[10292] <= 8'h00
            reg_file[10293] <= 8'h00
            reg_file[10294] <= 8'h00
            reg_file[10295] <= 8'h00
            reg_file[10296] <= 8'h00
            reg_file[10297] <= 8'h00
            reg_file[10298] <= 8'h00
            reg_file[10299] <= 8'h00
            reg_file[10300] <= 8'h00
            reg_file[10301] <= 8'h00
            reg_file[10302] <= 8'h00
            reg_file[10303] <= 8'h00
            reg_file[10304] <= 8'h00
            reg_file[10305] <= 8'h00
            reg_file[10306] <= 8'h00
            reg_file[10307] <= 8'h00
            reg_file[10308] <= 8'h00
            reg_file[10309] <= 8'h00
            reg_file[10310] <= 8'h00
            reg_file[10311] <= 8'h00
            reg_file[10312] <= 8'h00
            reg_file[10313] <= 8'h00
            reg_file[10314] <= 8'h00
            reg_file[10315] <= 8'h00
            reg_file[10316] <= 8'h00
            reg_file[10317] <= 8'h00
            reg_file[10318] <= 8'h00
            reg_file[10319] <= 8'h00
            reg_file[10320] <= 8'h00
            reg_file[10321] <= 8'h00
            reg_file[10322] <= 8'h00
            reg_file[10323] <= 8'h00
            reg_file[10324] <= 8'h00
            reg_file[10325] <= 8'h00
            reg_file[10326] <= 8'h00
            reg_file[10327] <= 8'h00
            reg_file[10328] <= 8'h00
            reg_file[10329] <= 8'h00
            reg_file[10330] <= 8'h00
            reg_file[10331] <= 8'h00
            reg_file[10332] <= 8'h00
            reg_file[10333] <= 8'h00
            reg_file[10334] <= 8'h00
            reg_file[10335] <= 8'h00
            reg_file[10336] <= 8'h00
            reg_file[10337] <= 8'h00
            reg_file[10338] <= 8'h00
            reg_file[10339] <= 8'h00
            reg_file[10340] <= 8'h00
            reg_file[10341] <= 8'h00
            reg_file[10342] <= 8'h00
            reg_file[10343] <= 8'h00
            reg_file[10344] <= 8'h00
            reg_file[10345] <= 8'h00
            reg_file[10346] <= 8'h00
            reg_file[10347] <= 8'h00
            reg_file[10348] <= 8'h00
            reg_file[10349] <= 8'h00
            reg_file[10350] <= 8'h00
            reg_file[10351] <= 8'h00
            reg_file[10352] <= 8'h00
            reg_file[10353] <= 8'h00
            reg_file[10354] <= 8'h00
            reg_file[10355] <= 8'h00
            reg_file[10356] <= 8'h00
            reg_file[10357] <= 8'h00
            reg_file[10358] <= 8'h00
            reg_file[10359] <= 8'h00
            reg_file[10360] <= 8'h00
            reg_file[10361] <= 8'h00
            reg_file[10362] <= 8'h00
            reg_file[10363] <= 8'h00
            reg_file[10364] <= 8'h00
            reg_file[10365] <= 8'h00
            reg_file[10366] <= 8'h00
            reg_file[10367] <= 8'h00
            reg_file[10368] <= 8'h00
            reg_file[10369] <= 8'h00
            reg_file[10370] <= 8'h00
            reg_file[10371] <= 8'h00
            reg_file[10372] <= 8'h00
            reg_file[10373] <= 8'h00
            reg_file[10374] <= 8'h00
            reg_file[10375] <= 8'h00
            reg_file[10376] <= 8'h00
            reg_file[10377] <= 8'h00
            reg_file[10378] <= 8'h00
            reg_file[10379] <= 8'h00
            reg_file[10380] <= 8'h00
            reg_file[10381] <= 8'h00
            reg_file[10382] <= 8'h00
            reg_file[10383] <= 8'h00
            reg_file[10384] <= 8'h00
            reg_file[10385] <= 8'h00
            reg_file[10386] <= 8'h00
            reg_file[10387] <= 8'h00
            reg_file[10388] <= 8'h00
            reg_file[10389] <= 8'h00
            reg_file[10390] <= 8'h00
            reg_file[10391] <= 8'h00
            reg_file[10392] <= 8'h00
            reg_file[10393] <= 8'h00
            reg_file[10394] <= 8'h00
            reg_file[10395] <= 8'h00
            reg_file[10396] <= 8'h00
            reg_file[10397] <= 8'h00
            reg_file[10398] <= 8'h00
            reg_file[10399] <= 8'h00
            reg_file[10400] <= 8'h00
            reg_file[10401] <= 8'h00
            reg_file[10402] <= 8'h00
            reg_file[10403] <= 8'h00
            reg_file[10404] <= 8'h00
            reg_file[10405] <= 8'h00
            reg_file[10406] <= 8'h00
            reg_file[10407] <= 8'h00
            reg_file[10408] <= 8'h00
            reg_file[10409] <= 8'h00
            reg_file[10410] <= 8'h00
            reg_file[10411] <= 8'h00
            reg_file[10412] <= 8'h00
            reg_file[10413] <= 8'h00
            reg_file[10414] <= 8'h00
            reg_file[10415] <= 8'h00
            reg_file[10416] <= 8'h00
            reg_file[10417] <= 8'h00
            reg_file[10418] <= 8'h00
            reg_file[10419] <= 8'h00
            reg_file[10420] <= 8'h00
            reg_file[10421] <= 8'h00
            reg_file[10422] <= 8'h00
            reg_file[10423] <= 8'h00
            reg_file[10424] <= 8'h00
            reg_file[10425] <= 8'h00
            reg_file[10426] <= 8'h00
            reg_file[10427] <= 8'h00
            reg_file[10428] <= 8'h00
            reg_file[10429] <= 8'h00
            reg_file[10430] <= 8'h00
            reg_file[10431] <= 8'h00
            reg_file[10432] <= 8'h00
            reg_file[10433] <= 8'h00
            reg_file[10434] <= 8'h00
            reg_file[10435] <= 8'h00
            reg_file[10436] <= 8'h00
            reg_file[10437] <= 8'h00
            reg_file[10438] <= 8'h00
            reg_file[10439] <= 8'h00
            reg_file[10440] <= 8'h00
            reg_file[10441] <= 8'h00
            reg_file[10442] <= 8'h00
            reg_file[10443] <= 8'h00
            reg_file[10444] <= 8'h00
            reg_file[10445] <= 8'h00
            reg_file[10446] <= 8'h00
            reg_file[10447] <= 8'h00
            reg_file[10448] <= 8'h00
            reg_file[10449] <= 8'h00
            reg_file[10450] <= 8'h00
            reg_file[10451] <= 8'h00
            reg_file[10452] <= 8'h00
            reg_file[10453] <= 8'h00
            reg_file[10454] <= 8'h00
            reg_file[10455] <= 8'h00
            reg_file[10456] <= 8'h00
            reg_file[10457] <= 8'h00
            reg_file[10458] <= 8'h00
            reg_file[10459] <= 8'h00
            reg_file[10460] <= 8'h00
            reg_file[10461] <= 8'h00
            reg_file[10462] <= 8'h00
            reg_file[10463] <= 8'h00
            reg_file[10464] <= 8'h00
            reg_file[10465] <= 8'h00
            reg_file[10466] <= 8'h00
            reg_file[10467] <= 8'h00
            reg_file[10468] <= 8'h00
            reg_file[10469] <= 8'h00
            reg_file[10470] <= 8'h00
            reg_file[10471] <= 8'h00
            reg_file[10472] <= 8'h00
            reg_file[10473] <= 8'h00
            reg_file[10474] <= 8'h00
            reg_file[10475] <= 8'h00
            reg_file[10476] <= 8'h00
            reg_file[10477] <= 8'h00
            reg_file[10478] <= 8'h00
            reg_file[10479] <= 8'h00
            reg_file[10480] <= 8'h00
            reg_file[10481] <= 8'h00
            reg_file[10482] <= 8'h00
            reg_file[10483] <= 8'h00
            reg_file[10484] <= 8'h00
            reg_file[10485] <= 8'h00
            reg_file[10486] <= 8'h00
            reg_file[10487] <= 8'h00
            reg_file[10488] <= 8'h00
            reg_file[10489] <= 8'h00
            reg_file[10490] <= 8'h00
            reg_file[10491] <= 8'h00
            reg_file[10492] <= 8'h00
            reg_file[10493] <= 8'h00
            reg_file[10494] <= 8'h00
            reg_file[10495] <= 8'h00
            reg_file[10496] <= 8'h00
            reg_file[10497] <= 8'h00
            reg_file[10498] <= 8'h00
            reg_file[10499] <= 8'h00
            reg_file[10500] <= 8'h00
            reg_file[10501] <= 8'h00
            reg_file[10502] <= 8'h00
            reg_file[10503] <= 8'h00
            reg_file[10504] <= 8'h00
            reg_file[10505] <= 8'h00
            reg_file[10506] <= 8'h00
            reg_file[10507] <= 8'h00
            reg_file[10508] <= 8'h00
            reg_file[10509] <= 8'h00
            reg_file[10510] <= 8'h00
            reg_file[10511] <= 8'h00
            reg_file[10512] <= 8'h00
            reg_file[10513] <= 8'h00
            reg_file[10514] <= 8'h00
            reg_file[10515] <= 8'h00
            reg_file[10516] <= 8'h00
            reg_file[10517] <= 8'h00
            reg_file[10518] <= 8'h00
            reg_file[10519] <= 8'h00
            reg_file[10520] <= 8'h00
            reg_file[10521] <= 8'h00
            reg_file[10522] <= 8'h00
            reg_file[10523] <= 8'h00
            reg_file[10524] <= 8'h00
            reg_file[10525] <= 8'h00
            reg_file[10526] <= 8'h00
            reg_file[10527] <= 8'h00
            reg_file[10528] <= 8'h00
            reg_file[10529] <= 8'h00
            reg_file[10530] <= 8'h00
            reg_file[10531] <= 8'h00
            reg_file[10532] <= 8'h00
            reg_file[10533] <= 8'h00
            reg_file[10534] <= 8'h00
            reg_file[10535] <= 8'h00
            reg_file[10536] <= 8'h00
            reg_file[10537] <= 8'h00
            reg_file[10538] <= 8'h00
            reg_file[10539] <= 8'h00
            reg_file[10540] <= 8'h00
            reg_file[10541] <= 8'h00
            reg_file[10542] <= 8'h00
            reg_file[10543] <= 8'h00
            reg_file[10544] <= 8'h00
            reg_file[10545] <= 8'h00
            reg_file[10546] <= 8'h00
            reg_file[10547] <= 8'h00
            reg_file[10548] <= 8'h00
            reg_file[10549] <= 8'h00
            reg_file[10550] <= 8'h00
            reg_file[10551] <= 8'h00
            reg_file[10552] <= 8'h00
            reg_file[10553] <= 8'h00
            reg_file[10554] <= 8'h00
            reg_file[10555] <= 8'h00
            reg_file[10556] <= 8'h00
            reg_file[10557] <= 8'h00
            reg_file[10558] <= 8'h00
            reg_file[10559] <= 8'h00
            reg_file[10560] <= 8'h00
            reg_file[10561] <= 8'h00
            reg_file[10562] <= 8'h00
            reg_file[10563] <= 8'h00
            reg_file[10564] <= 8'h00
            reg_file[10565] <= 8'h00
            reg_file[10566] <= 8'h00
            reg_file[10567] <= 8'h00
            reg_file[10568] <= 8'h00
            reg_file[10569] <= 8'h00
            reg_file[10570] <= 8'h00
            reg_file[10571] <= 8'h00
            reg_file[10572] <= 8'h00
            reg_file[10573] <= 8'h00
            reg_file[10574] <= 8'h00
            reg_file[10575] <= 8'h00
            reg_file[10576] <= 8'h00
            reg_file[10577] <= 8'h00
            reg_file[10578] <= 8'h00
            reg_file[10579] <= 8'h00
            reg_file[10580] <= 8'h00
            reg_file[10581] <= 8'h00
            reg_file[10582] <= 8'h00
            reg_file[10583] <= 8'h00
            reg_file[10584] <= 8'h00
            reg_file[10585] <= 8'h00
            reg_file[10586] <= 8'h00
            reg_file[10587] <= 8'h00
            reg_file[10588] <= 8'h00
            reg_file[10589] <= 8'h00
            reg_file[10590] <= 8'h00
            reg_file[10591] <= 8'h00
            reg_file[10592] <= 8'h00
            reg_file[10593] <= 8'h00
            reg_file[10594] <= 8'h00
            reg_file[10595] <= 8'h00
            reg_file[10596] <= 8'h00
            reg_file[10597] <= 8'h00
            reg_file[10598] <= 8'h00
            reg_file[10599] <= 8'h00
            reg_file[10600] <= 8'h00
            reg_file[10601] <= 8'h00
            reg_file[10602] <= 8'h00
            reg_file[10603] <= 8'h00
            reg_file[10604] <= 8'h00
            reg_file[10605] <= 8'h00
            reg_file[10606] <= 8'h00
            reg_file[10607] <= 8'h00
            reg_file[10608] <= 8'h00
            reg_file[10609] <= 8'h00
            reg_file[10610] <= 8'h00
            reg_file[10611] <= 8'h00
            reg_file[10612] <= 8'h00
            reg_file[10613] <= 8'h00
            reg_file[10614] <= 8'h00
            reg_file[10615] <= 8'h00
            reg_file[10616] <= 8'h00
            reg_file[10617] <= 8'h00
            reg_file[10618] <= 8'h00
            reg_file[10619] <= 8'h00
            reg_file[10620] <= 8'h00
            reg_file[10621] <= 8'h00
            reg_file[10622] <= 8'h00
            reg_file[10623] <= 8'h00
            reg_file[10624] <= 8'h00
            reg_file[10625] <= 8'h00
            reg_file[10626] <= 8'h00
            reg_file[10627] <= 8'h00
            reg_file[10628] <= 8'h00
            reg_file[10629] <= 8'h00
            reg_file[10630] <= 8'h00
            reg_file[10631] <= 8'h00
            reg_file[10632] <= 8'h00
            reg_file[10633] <= 8'h00
            reg_file[10634] <= 8'h00
            reg_file[10635] <= 8'h00
            reg_file[10636] <= 8'h00
            reg_file[10637] <= 8'h00
            reg_file[10638] <= 8'h00
            reg_file[10639] <= 8'h00
            reg_file[10640] <= 8'h00
            reg_file[10641] <= 8'h00
            reg_file[10642] <= 8'h00
            reg_file[10643] <= 8'h00
            reg_file[10644] <= 8'h00
            reg_file[10645] <= 8'h00
            reg_file[10646] <= 8'h00
            reg_file[10647] <= 8'h00
            reg_file[10648] <= 8'h00
            reg_file[10649] <= 8'h00
            reg_file[10650] <= 8'h00
            reg_file[10651] <= 8'h00
            reg_file[10652] <= 8'h00
            reg_file[10653] <= 8'h00
            reg_file[10654] <= 8'h00
            reg_file[10655] <= 8'h00
            reg_file[10656] <= 8'h00
            reg_file[10657] <= 8'h00
            reg_file[10658] <= 8'h00
            reg_file[10659] <= 8'h00
            reg_file[10660] <= 8'h00
            reg_file[10661] <= 8'h00
            reg_file[10662] <= 8'h00
            reg_file[10663] <= 8'h00
            reg_file[10664] <= 8'h00
            reg_file[10665] <= 8'h00
            reg_file[10666] <= 8'h00
            reg_file[10667] <= 8'h00
            reg_file[10668] <= 8'h00
            reg_file[10669] <= 8'h00
            reg_file[10670] <= 8'h00
            reg_file[10671] <= 8'h00
            reg_file[10672] <= 8'h00
            reg_file[10673] <= 8'h00
            reg_file[10674] <= 8'h00
            reg_file[10675] <= 8'h00
            reg_file[10676] <= 8'h00
            reg_file[10677] <= 8'h00
            reg_file[10678] <= 8'h00
            reg_file[10679] <= 8'h00
            reg_file[10680] <= 8'h00
            reg_file[10681] <= 8'h00
            reg_file[10682] <= 8'h00
            reg_file[10683] <= 8'h00
            reg_file[10684] <= 8'h00
            reg_file[10685] <= 8'h00
            reg_file[10686] <= 8'h00
            reg_file[10687] <= 8'h00
            reg_file[10688] <= 8'h00
            reg_file[10689] <= 8'h00
            reg_file[10690] <= 8'h00
            reg_file[10691] <= 8'h00
            reg_file[10692] <= 8'h00
            reg_file[10693] <= 8'h00
            reg_file[10694] <= 8'h00
            reg_file[10695] <= 8'h00
            reg_file[10696] <= 8'h00
            reg_file[10697] <= 8'h00
            reg_file[10698] <= 8'h00
            reg_file[10699] <= 8'h00
            reg_file[10700] <= 8'h00
            reg_file[10701] <= 8'h00
            reg_file[10702] <= 8'h00
            reg_file[10703] <= 8'h00
            reg_file[10704] <= 8'h00
            reg_file[10705] <= 8'h00
            reg_file[10706] <= 8'h00
            reg_file[10707] <= 8'h00
            reg_file[10708] <= 8'h00
            reg_file[10709] <= 8'h00
            reg_file[10710] <= 8'h00
            reg_file[10711] <= 8'h00
            reg_file[10712] <= 8'h00
            reg_file[10713] <= 8'h00
            reg_file[10714] <= 8'h00
            reg_file[10715] <= 8'h00
            reg_file[10716] <= 8'h00
            reg_file[10717] <= 8'h00
            reg_file[10718] <= 8'h00
            reg_file[10719] <= 8'h00
            reg_file[10720] <= 8'h00
            reg_file[10721] <= 8'h00
            reg_file[10722] <= 8'h00
            reg_file[10723] <= 8'h00
            reg_file[10724] <= 8'h00
            reg_file[10725] <= 8'h00
            reg_file[10726] <= 8'h00
            reg_file[10727] <= 8'h00
            reg_file[10728] <= 8'h00
            reg_file[10729] <= 8'h00
            reg_file[10730] <= 8'h00
            reg_file[10731] <= 8'h00
            reg_file[10732] <= 8'h00
            reg_file[10733] <= 8'h00
            reg_file[10734] <= 8'h00
            reg_file[10735] <= 8'h00
            reg_file[10736] <= 8'h00
            reg_file[10737] <= 8'h00
            reg_file[10738] <= 8'h00
            reg_file[10739] <= 8'h00
            reg_file[10740] <= 8'h00
            reg_file[10741] <= 8'h00
            reg_file[10742] <= 8'h00
            reg_file[10743] <= 8'h00
            reg_file[10744] <= 8'h00
            reg_file[10745] <= 8'h00
            reg_file[10746] <= 8'h00
            reg_file[10747] <= 8'h00
            reg_file[10748] <= 8'h00
            reg_file[10749] <= 8'h00
            reg_file[10750] <= 8'h00
            reg_file[10751] <= 8'h00
            reg_file[10752] <= 8'h00
            reg_file[10753] <= 8'h00
            reg_file[10754] <= 8'h00
            reg_file[10755] <= 8'h00
            reg_file[10756] <= 8'h00
            reg_file[10757] <= 8'h00
            reg_file[10758] <= 8'h00
            reg_file[10759] <= 8'h00
            reg_file[10760] <= 8'h00
            reg_file[10761] <= 8'h00
            reg_file[10762] <= 8'h00
            reg_file[10763] <= 8'h00
            reg_file[10764] <= 8'h00
            reg_file[10765] <= 8'h00
            reg_file[10766] <= 8'h00
            reg_file[10767] <= 8'h00
            reg_file[10768] <= 8'h00
            reg_file[10769] <= 8'h00
            reg_file[10770] <= 8'h00
            reg_file[10771] <= 8'h00
            reg_file[10772] <= 8'h00
            reg_file[10773] <= 8'h00
            reg_file[10774] <= 8'h00
            reg_file[10775] <= 8'h00
            reg_file[10776] <= 8'h00
            reg_file[10777] <= 8'h00
            reg_file[10778] <= 8'h00
            reg_file[10779] <= 8'h00
            reg_file[10780] <= 8'h00
            reg_file[10781] <= 8'h00
            reg_file[10782] <= 8'h00
            reg_file[10783] <= 8'h00
            reg_file[10784] <= 8'h00
            reg_file[10785] <= 8'h00
            reg_file[10786] <= 8'h00
            reg_file[10787] <= 8'h00
            reg_file[10788] <= 8'h00
            reg_file[10789] <= 8'h00
            reg_file[10790] <= 8'h00
            reg_file[10791] <= 8'h00
            reg_file[10792] <= 8'h00
            reg_file[10793] <= 8'h00
            reg_file[10794] <= 8'h00
            reg_file[10795] <= 8'h00
            reg_file[10796] <= 8'h00
            reg_file[10797] <= 8'h00
            reg_file[10798] <= 8'h00
            reg_file[10799] <= 8'h00
            reg_file[10800] <= 8'h00
            reg_file[10801] <= 8'h00
            reg_file[10802] <= 8'h00
            reg_file[10803] <= 8'h00
            reg_file[10804] <= 8'h00
            reg_file[10805] <= 8'h00
            reg_file[10806] <= 8'h00
            reg_file[10807] <= 8'h00
            reg_file[10808] <= 8'h00
            reg_file[10809] <= 8'h00
            reg_file[10810] <= 8'h00
            reg_file[10811] <= 8'h00
            reg_file[10812] <= 8'h00
            reg_file[10813] <= 8'h00
            reg_file[10814] <= 8'h00
            reg_file[10815] <= 8'h00
            reg_file[10816] <= 8'h00
            reg_file[10817] <= 8'h00
            reg_file[10818] <= 8'h00
            reg_file[10819] <= 8'h00
            reg_file[10820] <= 8'h00
            reg_file[10821] <= 8'h00
            reg_file[10822] <= 8'h00
            reg_file[10823] <= 8'h00
            reg_file[10824] <= 8'h00
            reg_file[10825] <= 8'h00
            reg_file[10826] <= 8'h00
            reg_file[10827] <= 8'h00
            reg_file[10828] <= 8'h00
            reg_file[10829] <= 8'h00
            reg_file[10830] <= 8'h00
            reg_file[10831] <= 8'h00
            reg_file[10832] <= 8'h00
            reg_file[10833] <= 8'h00
            reg_file[10834] <= 8'h00
            reg_file[10835] <= 8'h00
            reg_file[10836] <= 8'h00
            reg_file[10837] <= 8'h00
            reg_file[10838] <= 8'h00
            reg_file[10839] <= 8'h00
            reg_file[10840] <= 8'h00
            reg_file[10841] <= 8'h00
            reg_file[10842] <= 8'h00
            reg_file[10843] <= 8'h00
            reg_file[10844] <= 8'h00
            reg_file[10845] <= 8'h00
            reg_file[10846] <= 8'h00
            reg_file[10847] <= 8'h00
            reg_file[10848] <= 8'h00
            reg_file[10849] <= 8'h00
            reg_file[10850] <= 8'h00
            reg_file[10851] <= 8'h00
            reg_file[10852] <= 8'h00
            reg_file[10853] <= 8'h00
            reg_file[10854] <= 8'h00
            reg_file[10855] <= 8'h00
            reg_file[10856] <= 8'h00
            reg_file[10857] <= 8'h00
            reg_file[10858] <= 8'h00
            reg_file[10859] <= 8'h00
            reg_file[10860] <= 8'h00
            reg_file[10861] <= 8'h00
            reg_file[10862] <= 8'h00
            reg_file[10863] <= 8'h00
            reg_file[10864] <= 8'h00
            reg_file[10865] <= 8'h00
            reg_file[10866] <= 8'h00
            reg_file[10867] <= 8'h00
            reg_file[10868] <= 8'h00
            reg_file[10869] <= 8'h00
            reg_file[10870] <= 8'h00
            reg_file[10871] <= 8'h00
            reg_file[10872] <= 8'h00
            reg_file[10873] <= 8'h00
            reg_file[10874] <= 8'h00
            reg_file[10875] <= 8'h00
            reg_file[10876] <= 8'h00
            reg_file[10877] <= 8'h00
            reg_file[10878] <= 8'h00
            reg_file[10879] <= 8'h00
            reg_file[10880] <= 8'h00
            reg_file[10881] <= 8'h00
            reg_file[10882] <= 8'h00
            reg_file[10883] <= 8'h00
            reg_file[10884] <= 8'h00
            reg_file[10885] <= 8'h00
            reg_file[10886] <= 8'h00
            reg_file[10887] <= 8'h00
            reg_file[10888] <= 8'h00
            reg_file[10889] <= 8'h00
            reg_file[10890] <= 8'h00
            reg_file[10891] <= 8'h00
            reg_file[10892] <= 8'h00
            reg_file[10893] <= 8'h00
            reg_file[10894] <= 8'h00
            reg_file[10895] <= 8'h00
            reg_file[10896] <= 8'h00
            reg_file[10897] <= 8'h00
            reg_file[10898] <= 8'h00
            reg_file[10899] <= 8'h00
            reg_file[10900] <= 8'h00
            reg_file[10901] <= 8'h00
            reg_file[10902] <= 8'h00
            reg_file[10903] <= 8'h00
            reg_file[10904] <= 8'h00
            reg_file[10905] <= 8'h00
            reg_file[10906] <= 8'h00
            reg_file[10907] <= 8'h00
            reg_file[10908] <= 8'h00
            reg_file[10909] <= 8'h00
            reg_file[10910] <= 8'h00
            reg_file[10911] <= 8'h00
            reg_file[10912] <= 8'h00
            reg_file[10913] <= 8'h00
            reg_file[10914] <= 8'h00
            reg_file[10915] <= 8'h00
            reg_file[10916] <= 8'h00
            reg_file[10917] <= 8'h00
            reg_file[10918] <= 8'h00
            reg_file[10919] <= 8'h00
            reg_file[10920] <= 8'h00
            reg_file[10921] <= 8'h00
            reg_file[10922] <= 8'h00
            reg_file[10923] <= 8'h00
            reg_file[10924] <= 8'h00
            reg_file[10925] <= 8'h00
            reg_file[10926] <= 8'h00
            reg_file[10927] <= 8'h00
            reg_file[10928] <= 8'h00
            reg_file[10929] <= 8'h00
            reg_file[10930] <= 8'h00
            reg_file[10931] <= 8'h00
            reg_file[10932] <= 8'h00
            reg_file[10933] <= 8'h00
            reg_file[10934] <= 8'h00
            reg_file[10935] <= 8'h00
            reg_file[10936] <= 8'h00
            reg_file[10937] <= 8'h00
            reg_file[10938] <= 8'h00
            reg_file[10939] <= 8'h00
            reg_file[10940] <= 8'h00
            reg_file[10941] <= 8'h00
            reg_file[10942] <= 8'h00
            reg_file[10943] <= 8'h00
            reg_file[10944] <= 8'h00
            reg_file[10945] <= 8'h00
            reg_file[10946] <= 8'h00
            reg_file[10947] <= 8'h00
            reg_file[10948] <= 8'h00
            reg_file[10949] <= 8'h00
            reg_file[10950] <= 8'h00
            reg_file[10951] <= 8'h00
            reg_file[10952] <= 8'h00
            reg_file[10953] <= 8'h00
            reg_file[10954] <= 8'h00
            reg_file[10955] <= 8'h00
            reg_file[10956] <= 8'h00
            reg_file[10957] <= 8'h00
            reg_file[10958] <= 8'h00
            reg_file[10959] <= 8'h00
            reg_file[10960] <= 8'h00
            reg_file[10961] <= 8'h00
            reg_file[10962] <= 8'h00
            reg_file[10963] <= 8'h00
            reg_file[10964] <= 8'h00
            reg_file[10965] <= 8'h00
            reg_file[10966] <= 8'h00
            reg_file[10967] <= 8'h00
            reg_file[10968] <= 8'h00
            reg_file[10969] <= 8'h00
            reg_file[10970] <= 8'h00
            reg_file[10971] <= 8'h00
            reg_file[10972] <= 8'h00
            reg_file[10973] <= 8'h00
            reg_file[10974] <= 8'h00
            reg_file[10975] <= 8'h00
            reg_file[10976] <= 8'h00
            reg_file[10977] <= 8'h00
            reg_file[10978] <= 8'h00
            reg_file[10979] <= 8'h00
            reg_file[10980] <= 8'h00
            reg_file[10981] <= 8'h00
            reg_file[10982] <= 8'h00
            reg_file[10983] <= 8'h00
            reg_file[10984] <= 8'h00
            reg_file[10985] <= 8'h00
            reg_file[10986] <= 8'h00
            reg_file[10987] <= 8'h00
            reg_file[10988] <= 8'h00
            reg_file[10989] <= 8'h00
            reg_file[10990] <= 8'h00
            reg_file[10991] <= 8'h00
            reg_file[10992] <= 8'h00
            reg_file[10993] <= 8'h00
            reg_file[10994] <= 8'h00
            reg_file[10995] <= 8'h00
            reg_file[10996] <= 8'h00
            reg_file[10997] <= 8'h00
            reg_file[10998] <= 8'h00
            reg_file[10999] <= 8'h00
            reg_file[11000] <= 8'h00
            reg_file[11001] <= 8'h00
            reg_file[11002] <= 8'h00
            reg_file[11003] <= 8'h00
            reg_file[11004] <= 8'h00
            reg_file[11005] <= 8'h00
            reg_file[11006] <= 8'h00
            reg_file[11007] <= 8'h00
            reg_file[11008] <= 8'h00
            reg_file[11009] <= 8'h00
            reg_file[11010] <= 8'h00
            reg_file[11011] <= 8'h00
            reg_file[11012] <= 8'h00
            reg_file[11013] <= 8'h00
            reg_file[11014] <= 8'h00
            reg_file[11015] <= 8'h00
            reg_file[11016] <= 8'h00
            reg_file[11017] <= 8'h00
            reg_file[11018] <= 8'h00
            reg_file[11019] <= 8'h00
            reg_file[11020] <= 8'h00
            reg_file[11021] <= 8'h00
            reg_file[11022] <= 8'h00
            reg_file[11023] <= 8'h00
            reg_file[11024] <= 8'h00
            reg_file[11025] <= 8'h00
            reg_file[11026] <= 8'h00
            reg_file[11027] <= 8'h00
            reg_file[11028] <= 8'h00
            reg_file[11029] <= 8'h00
            reg_file[11030] <= 8'h00
            reg_file[11031] <= 8'h00
            reg_file[11032] <= 8'h00
            reg_file[11033] <= 8'h00
            reg_file[11034] <= 8'h00
            reg_file[11035] <= 8'h00
            reg_file[11036] <= 8'h00
            reg_file[11037] <= 8'h00
            reg_file[11038] <= 8'h00
            reg_file[11039] <= 8'h00
            reg_file[11040] <= 8'h00
            reg_file[11041] <= 8'h00
            reg_file[11042] <= 8'h00
            reg_file[11043] <= 8'h00
            reg_file[11044] <= 8'h00
            reg_file[11045] <= 8'h00
            reg_file[11046] <= 8'h00
            reg_file[11047] <= 8'h00
            reg_file[11048] <= 8'h00
            reg_file[11049] <= 8'h00
            reg_file[11050] <= 8'h00
            reg_file[11051] <= 8'h00
            reg_file[11052] <= 8'h00
            reg_file[11053] <= 8'h00
            reg_file[11054] <= 8'h00
            reg_file[11055] <= 8'h00
            reg_file[11056] <= 8'h00
            reg_file[11057] <= 8'h00
            reg_file[11058] <= 8'h00
            reg_file[11059] <= 8'h00
            reg_file[11060] <= 8'h00
            reg_file[11061] <= 8'h00
            reg_file[11062] <= 8'h00
            reg_file[11063] <= 8'h00
            reg_file[11064] <= 8'h00
            reg_file[11065] <= 8'h00
            reg_file[11066] <= 8'h00
            reg_file[11067] <= 8'h00
            reg_file[11068] <= 8'h00
            reg_file[11069] <= 8'h00
            reg_file[11070] <= 8'h00
            reg_file[11071] <= 8'h00
            reg_file[11072] <= 8'h00
            reg_file[11073] <= 8'h00
            reg_file[11074] <= 8'h00
            reg_file[11075] <= 8'h00
            reg_file[11076] <= 8'h00
            reg_file[11077] <= 8'h00
            reg_file[11078] <= 8'h00
            reg_file[11079] <= 8'h00
            reg_file[11080] <= 8'h00
            reg_file[11081] <= 8'h00
            reg_file[11082] <= 8'h00
            reg_file[11083] <= 8'h00
            reg_file[11084] <= 8'h00
            reg_file[11085] <= 8'h00
            reg_file[11086] <= 8'h00
            reg_file[11087] <= 8'h00
            reg_file[11088] <= 8'h00
            reg_file[11089] <= 8'h00
            reg_file[11090] <= 8'h00
            reg_file[11091] <= 8'h00
            reg_file[11092] <= 8'h00
            reg_file[11093] <= 8'h00
            reg_file[11094] <= 8'h00
            reg_file[11095] <= 8'h00
            reg_file[11096] <= 8'h00
            reg_file[11097] <= 8'h00
            reg_file[11098] <= 8'h00
            reg_file[11099] <= 8'h00
            reg_file[11100] <= 8'h00
            reg_file[11101] <= 8'h00
            reg_file[11102] <= 8'h00
            reg_file[11103] <= 8'h00
            reg_file[11104] <= 8'h00
            reg_file[11105] <= 8'h00
            reg_file[11106] <= 8'h00
            reg_file[11107] <= 8'h00
            reg_file[11108] <= 8'h00
            reg_file[11109] <= 8'h00
            reg_file[11110] <= 8'h00
            reg_file[11111] <= 8'h00
            reg_file[11112] <= 8'h00
            reg_file[11113] <= 8'h00
            reg_file[11114] <= 8'h00
            reg_file[11115] <= 8'h00
            reg_file[11116] <= 8'h00
            reg_file[11117] <= 8'h00
            reg_file[11118] <= 8'h00
            reg_file[11119] <= 8'h00
            reg_file[11120] <= 8'h00
            reg_file[11121] <= 8'h00
            reg_file[11122] <= 8'h00
            reg_file[11123] <= 8'h00
            reg_file[11124] <= 8'h00
            reg_file[11125] <= 8'h00
            reg_file[11126] <= 8'h00
            reg_file[11127] <= 8'h00
            reg_file[11128] <= 8'h00
            reg_file[11129] <= 8'h00
            reg_file[11130] <= 8'h00
            reg_file[11131] <= 8'h00
            reg_file[11132] <= 8'h00
            reg_file[11133] <= 8'h00
            reg_file[11134] <= 8'h00
            reg_file[11135] <= 8'h00
            reg_file[11136] <= 8'h00
            reg_file[11137] <= 8'h00
            reg_file[11138] <= 8'h00
            reg_file[11139] <= 8'h00
            reg_file[11140] <= 8'h00
            reg_file[11141] <= 8'h00
            reg_file[11142] <= 8'h00
            reg_file[11143] <= 8'h00
            reg_file[11144] <= 8'h00
            reg_file[11145] <= 8'h00
            reg_file[11146] <= 8'h00
            reg_file[11147] <= 8'h00
            reg_file[11148] <= 8'h00
            reg_file[11149] <= 8'h00
            reg_file[11150] <= 8'h00
            reg_file[11151] <= 8'h00
            reg_file[11152] <= 8'h00
            reg_file[11153] <= 8'h00
            reg_file[11154] <= 8'h00
            reg_file[11155] <= 8'h00
            reg_file[11156] <= 8'h00
            reg_file[11157] <= 8'h00
            reg_file[11158] <= 8'h00
            reg_file[11159] <= 8'h00
            reg_file[11160] <= 8'h00
            reg_file[11161] <= 8'h00
            reg_file[11162] <= 8'h00
            reg_file[11163] <= 8'h00
            reg_file[11164] <= 8'h00
            reg_file[11165] <= 8'h00
            reg_file[11166] <= 8'h00
            reg_file[11167] <= 8'h00
            reg_file[11168] <= 8'h00
            reg_file[11169] <= 8'h00
            reg_file[11170] <= 8'h00
            reg_file[11171] <= 8'h00
            reg_file[11172] <= 8'h00
            reg_file[11173] <= 8'h00
            reg_file[11174] <= 8'h00
            reg_file[11175] <= 8'h00
            reg_file[11176] <= 8'h00
            reg_file[11177] <= 8'h00
            reg_file[11178] <= 8'h00
            reg_file[11179] <= 8'h00
            reg_file[11180] <= 8'h00
            reg_file[11181] <= 8'h00
            reg_file[11182] <= 8'h00
            reg_file[11183] <= 8'h00
            reg_file[11184] <= 8'h00
            reg_file[11185] <= 8'h00
            reg_file[11186] <= 8'h00
            reg_file[11187] <= 8'h00
            reg_file[11188] <= 8'h00
            reg_file[11189] <= 8'h00
            reg_file[11190] <= 8'h00
            reg_file[11191] <= 8'h00
            reg_file[11192] <= 8'h00
            reg_file[11193] <= 8'h00
            reg_file[11194] <= 8'h00
            reg_file[11195] <= 8'h00
            reg_file[11196] <= 8'h00
            reg_file[11197] <= 8'h00
            reg_file[11198] <= 8'h00
            reg_file[11199] <= 8'h00
            reg_file[11200] <= 8'h00
            reg_file[11201] <= 8'h00
            reg_file[11202] <= 8'h00
            reg_file[11203] <= 8'h00
            reg_file[11204] <= 8'h00
            reg_file[11205] <= 8'h00
            reg_file[11206] <= 8'h00
            reg_file[11207] <= 8'h00
            reg_file[11208] <= 8'h00
            reg_file[11209] <= 8'h00
            reg_file[11210] <= 8'h00
            reg_file[11211] <= 8'h00
            reg_file[11212] <= 8'h00
            reg_file[11213] <= 8'h00
            reg_file[11214] <= 8'h00
            reg_file[11215] <= 8'h00
            reg_file[11216] <= 8'h00
            reg_file[11217] <= 8'h00
            reg_file[11218] <= 8'h00
            reg_file[11219] <= 8'h00
            reg_file[11220] <= 8'h00
            reg_file[11221] <= 8'h00
            reg_file[11222] <= 8'h00
            reg_file[11223] <= 8'h00
            reg_file[11224] <= 8'h00
            reg_file[11225] <= 8'h00
            reg_file[11226] <= 8'h00
            reg_file[11227] <= 8'h00
            reg_file[11228] <= 8'h00
            reg_file[11229] <= 8'h00
            reg_file[11230] <= 8'h00
            reg_file[11231] <= 8'h00
            reg_file[11232] <= 8'h00
            reg_file[11233] <= 8'h00
            reg_file[11234] <= 8'h00
            reg_file[11235] <= 8'h00
            reg_file[11236] <= 8'h00
            reg_file[11237] <= 8'h00
            reg_file[11238] <= 8'h00
            reg_file[11239] <= 8'h00
            reg_file[11240] <= 8'h00
            reg_file[11241] <= 8'h00
            reg_file[11242] <= 8'h00
            reg_file[11243] <= 8'h00
            reg_file[11244] <= 8'h00
            reg_file[11245] <= 8'h00
            reg_file[11246] <= 8'h00
            reg_file[11247] <= 8'h00
            reg_file[11248] <= 8'h00
            reg_file[11249] <= 8'h00
            reg_file[11250] <= 8'h00
            reg_file[11251] <= 8'h00
            reg_file[11252] <= 8'h00
            reg_file[11253] <= 8'h00
            reg_file[11254] <= 8'h00
            reg_file[11255] <= 8'h00
            reg_file[11256] <= 8'h00
            reg_file[11257] <= 8'h00
            reg_file[11258] <= 8'h00
            reg_file[11259] <= 8'h00
            reg_file[11260] <= 8'h00
            reg_file[11261] <= 8'h00
            reg_file[11262] <= 8'h00
            reg_file[11263] <= 8'h00
            reg_file[11264] <= 8'h00
            reg_file[11265] <= 8'h00
            reg_file[11266] <= 8'h00
            reg_file[11267] <= 8'h00
            reg_file[11268] <= 8'h00
            reg_file[11269] <= 8'h00
            reg_file[11270] <= 8'h00
            reg_file[11271] <= 8'h00
            reg_file[11272] <= 8'h00
            reg_file[11273] <= 8'h00
            reg_file[11274] <= 8'h00
            reg_file[11275] <= 8'h00
            reg_file[11276] <= 8'h00
            reg_file[11277] <= 8'h00
            reg_file[11278] <= 8'h00
            reg_file[11279] <= 8'h00
            reg_file[11280] <= 8'h00
            reg_file[11281] <= 8'h00
            reg_file[11282] <= 8'h00
            reg_file[11283] <= 8'h00
            reg_file[11284] <= 8'h00
            reg_file[11285] <= 8'h00
            reg_file[11286] <= 8'h00
            reg_file[11287] <= 8'h00
            reg_file[11288] <= 8'h00
            reg_file[11289] <= 8'h00
            reg_file[11290] <= 8'h00
            reg_file[11291] <= 8'h00
            reg_file[11292] <= 8'h00
            reg_file[11293] <= 8'h00
            reg_file[11294] <= 8'h00
            reg_file[11295] <= 8'h00
            reg_file[11296] <= 8'h00
            reg_file[11297] <= 8'h00
            reg_file[11298] <= 8'h00
            reg_file[11299] <= 8'h00
            reg_file[11300] <= 8'h00
            reg_file[11301] <= 8'h00
            reg_file[11302] <= 8'h00
            reg_file[11303] <= 8'h00
            reg_file[11304] <= 8'h00
            reg_file[11305] <= 8'h00
            reg_file[11306] <= 8'h00
            reg_file[11307] <= 8'h00
            reg_file[11308] <= 8'h00
            reg_file[11309] <= 8'h00
            reg_file[11310] <= 8'h00
            reg_file[11311] <= 8'h00
            reg_file[11312] <= 8'h00
            reg_file[11313] <= 8'h00
            reg_file[11314] <= 8'h00
            reg_file[11315] <= 8'h00
            reg_file[11316] <= 8'h00
            reg_file[11317] <= 8'h00
            reg_file[11318] <= 8'h00
            reg_file[11319] <= 8'h00
            reg_file[11320] <= 8'h00
            reg_file[11321] <= 8'h00
            reg_file[11322] <= 8'h00
            reg_file[11323] <= 8'h00
            reg_file[11324] <= 8'h00
            reg_file[11325] <= 8'h00
            reg_file[11326] <= 8'h00
            reg_file[11327] <= 8'h00
            reg_file[11328] <= 8'h00
            reg_file[11329] <= 8'h00
            reg_file[11330] <= 8'h00
            reg_file[11331] <= 8'h00
            reg_file[11332] <= 8'h00
            reg_file[11333] <= 8'h00
            reg_file[11334] <= 8'h00
            reg_file[11335] <= 8'h00
            reg_file[11336] <= 8'h00
            reg_file[11337] <= 8'h00
            reg_file[11338] <= 8'h00
            reg_file[11339] <= 8'h00
            reg_file[11340] <= 8'h00
            reg_file[11341] <= 8'h00
            reg_file[11342] <= 8'h00
            reg_file[11343] <= 8'h00
            reg_file[11344] <= 8'h00
            reg_file[11345] <= 8'h00
            reg_file[11346] <= 8'h00
            reg_file[11347] <= 8'h00
            reg_file[11348] <= 8'h00
            reg_file[11349] <= 8'h00
            reg_file[11350] <= 8'h00
            reg_file[11351] <= 8'h00
            reg_file[11352] <= 8'h00
            reg_file[11353] <= 8'h00
            reg_file[11354] <= 8'h00
            reg_file[11355] <= 8'h00
            reg_file[11356] <= 8'h00
            reg_file[11357] <= 8'h00
            reg_file[11358] <= 8'h00
            reg_file[11359] <= 8'h00
            reg_file[11360] <= 8'h00
            reg_file[11361] <= 8'h00
            reg_file[11362] <= 8'h00
            reg_file[11363] <= 8'h00
            reg_file[11364] <= 8'h00
            reg_file[11365] <= 8'h00
            reg_file[11366] <= 8'h00
            reg_file[11367] <= 8'h00
            reg_file[11368] <= 8'h00
            reg_file[11369] <= 8'h00
            reg_file[11370] <= 8'h00
            reg_file[11371] <= 8'h00
            reg_file[11372] <= 8'h00
            reg_file[11373] <= 8'h00
            reg_file[11374] <= 8'h00
            reg_file[11375] <= 8'h00
            reg_file[11376] <= 8'h00
            reg_file[11377] <= 8'h00
            reg_file[11378] <= 8'h00
            reg_file[11379] <= 8'h00
            reg_file[11380] <= 8'h00
            reg_file[11381] <= 8'h00
            reg_file[11382] <= 8'h00
            reg_file[11383] <= 8'h00
            reg_file[11384] <= 8'h00
            reg_file[11385] <= 8'h00
            reg_file[11386] <= 8'h00
            reg_file[11387] <= 8'h00
            reg_file[11388] <= 8'h00
            reg_file[11389] <= 8'h00
            reg_file[11390] <= 8'h00
            reg_file[11391] <= 8'h00
            reg_file[11392] <= 8'h00
            reg_file[11393] <= 8'h00
            reg_file[11394] <= 8'h00
            reg_file[11395] <= 8'h00
            reg_file[11396] <= 8'h00
            reg_file[11397] <= 8'h00
            reg_file[11398] <= 8'h00
            reg_file[11399] <= 8'h00
            reg_file[11400] <= 8'h00
            reg_file[11401] <= 8'h00
            reg_file[11402] <= 8'h00
            reg_file[11403] <= 8'h00
            reg_file[11404] <= 8'h00
            reg_file[11405] <= 8'h00
            reg_file[11406] <= 8'h00
            reg_file[11407] <= 8'h00
            reg_file[11408] <= 8'h00
            reg_file[11409] <= 8'h00
            reg_file[11410] <= 8'h00
            reg_file[11411] <= 8'h00
            reg_file[11412] <= 8'h00
            reg_file[11413] <= 8'h00
            reg_file[11414] <= 8'h00
            reg_file[11415] <= 8'h00
            reg_file[11416] <= 8'h00
            reg_file[11417] <= 8'h00
            reg_file[11418] <= 8'h00
            reg_file[11419] <= 8'h00
            reg_file[11420] <= 8'h00
            reg_file[11421] <= 8'h00
            reg_file[11422] <= 8'h00
            reg_file[11423] <= 8'h00
            reg_file[11424] <= 8'h00
            reg_file[11425] <= 8'h00
            reg_file[11426] <= 8'h00
            reg_file[11427] <= 8'h00
            reg_file[11428] <= 8'h00
            reg_file[11429] <= 8'h00
            reg_file[11430] <= 8'h00
            reg_file[11431] <= 8'h00
            reg_file[11432] <= 8'h00
            reg_file[11433] <= 8'h00
            reg_file[11434] <= 8'h00
            reg_file[11435] <= 8'h00
            reg_file[11436] <= 8'h00
            reg_file[11437] <= 8'h00
            reg_file[11438] <= 8'h00
            reg_file[11439] <= 8'h00
            reg_file[11440] <= 8'h00
            reg_file[11441] <= 8'h00
            reg_file[11442] <= 8'h00
            reg_file[11443] <= 8'h00
            reg_file[11444] <= 8'h00
            reg_file[11445] <= 8'h00
            reg_file[11446] <= 8'h00
            reg_file[11447] <= 8'h00
            reg_file[11448] <= 8'h00
            reg_file[11449] <= 8'h00
            reg_file[11450] <= 8'h00
            reg_file[11451] <= 8'h00
            reg_file[11452] <= 8'h00
            reg_file[11453] <= 8'h00
            reg_file[11454] <= 8'h00
            reg_file[11455] <= 8'h00
            reg_file[11456] <= 8'h00
            reg_file[11457] <= 8'h00
            reg_file[11458] <= 8'h00
            reg_file[11459] <= 8'h00
            reg_file[11460] <= 8'h00
            reg_file[11461] <= 8'h00
            reg_file[11462] <= 8'h00
            reg_file[11463] <= 8'h00
            reg_file[11464] <= 8'h00
            reg_file[11465] <= 8'h00
            reg_file[11466] <= 8'h00
            reg_file[11467] <= 8'h00
            reg_file[11468] <= 8'h00
            reg_file[11469] <= 8'h00
            reg_file[11470] <= 8'h00
            reg_file[11471] <= 8'h00
            reg_file[11472] <= 8'h00
            reg_file[11473] <= 8'h00
            reg_file[11474] <= 8'h00
            reg_file[11475] <= 8'h00
            reg_file[11476] <= 8'h00
            reg_file[11477] <= 8'h00
            reg_file[11478] <= 8'h00
            reg_file[11479] <= 8'h00
            reg_file[11480] <= 8'h00
            reg_file[11481] <= 8'h00
            reg_file[11482] <= 8'h00
            reg_file[11483] <= 8'h00
            reg_file[11484] <= 8'h00
            reg_file[11485] <= 8'h00
            reg_file[11486] <= 8'h00
            reg_file[11487] <= 8'h00
            reg_file[11488] <= 8'h00
            reg_file[11489] <= 8'h00
            reg_file[11490] <= 8'h00
            reg_file[11491] <= 8'h00
            reg_file[11492] <= 8'h00
            reg_file[11493] <= 8'h00
            reg_file[11494] <= 8'h00
            reg_file[11495] <= 8'h00
            reg_file[11496] <= 8'h00
            reg_file[11497] <= 8'h00
            reg_file[11498] <= 8'h00
            reg_file[11499] <= 8'h00
            reg_file[11500] <= 8'h00
            reg_file[11501] <= 8'h00
            reg_file[11502] <= 8'h00
            reg_file[11503] <= 8'h00
            reg_file[11504] <= 8'h00
            reg_file[11505] <= 8'h00
            reg_file[11506] <= 8'h00
            reg_file[11507] <= 8'h00
            reg_file[11508] <= 8'h00
            reg_file[11509] <= 8'h00
            reg_file[11510] <= 8'h00
            reg_file[11511] <= 8'h00
            reg_file[11512] <= 8'h00
            reg_file[11513] <= 8'h00
            reg_file[11514] <= 8'h00
            reg_file[11515] <= 8'h00
            reg_file[11516] <= 8'h00
            reg_file[11517] <= 8'h00
            reg_file[11518] <= 8'h00
            reg_file[11519] <= 8'h00
            reg_file[11520] <= 8'h00
            reg_file[11521] <= 8'h00
            reg_file[11522] <= 8'h00
            reg_file[11523] <= 8'h00
            reg_file[11524] <= 8'h00
            reg_file[11525] <= 8'h00
            reg_file[11526] <= 8'h00
            reg_file[11527] <= 8'h00
            reg_file[11528] <= 8'h00
            reg_file[11529] <= 8'h00
            reg_file[11530] <= 8'h00
            reg_file[11531] <= 8'h00
            reg_file[11532] <= 8'h00
            reg_file[11533] <= 8'h00
            reg_file[11534] <= 8'h00
            reg_file[11535] <= 8'h00
            reg_file[11536] <= 8'h00
            reg_file[11537] <= 8'h00
            reg_file[11538] <= 8'h00
            reg_file[11539] <= 8'h00
            reg_file[11540] <= 8'h00
            reg_file[11541] <= 8'h00
            reg_file[11542] <= 8'h00
            reg_file[11543] <= 8'h00
            reg_file[11544] <= 8'h00
            reg_file[11545] <= 8'h00
            reg_file[11546] <= 8'h00
            reg_file[11547] <= 8'h00
            reg_file[11548] <= 8'h00
            reg_file[11549] <= 8'h00
            reg_file[11550] <= 8'h00
            reg_file[11551] <= 8'h00
            reg_file[11552] <= 8'h00
            reg_file[11553] <= 8'h00
            reg_file[11554] <= 8'h00
            reg_file[11555] <= 8'h00
            reg_file[11556] <= 8'h00
            reg_file[11557] <= 8'h00
            reg_file[11558] <= 8'h00
            reg_file[11559] <= 8'h00
            reg_file[11560] <= 8'h00
            reg_file[11561] <= 8'h00
            reg_file[11562] <= 8'h00
            reg_file[11563] <= 8'h00
            reg_file[11564] <= 8'h00
            reg_file[11565] <= 8'h00
            reg_file[11566] <= 8'h00
            reg_file[11567] <= 8'h00
            reg_file[11568] <= 8'h00
            reg_file[11569] <= 8'h00
            reg_file[11570] <= 8'h00
            reg_file[11571] <= 8'h00
            reg_file[11572] <= 8'h00
            reg_file[11573] <= 8'h00
            reg_file[11574] <= 8'h00
            reg_file[11575] <= 8'h00
            reg_file[11576] <= 8'h00
            reg_file[11577] <= 8'h00
            reg_file[11578] <= 8'h00
            reg_file[11579] <= 8'h00
            reg_file[11580] <= 8'h00
            reg_file[11581] <= 8'h00
            reg_file[11582] <= 8'h00
            reg_file[11583] <= 8'h00
            reg_file[11584] <= 8'h00
            reg_file[11585] <= 8'h00
            reg_file[11586] <= 8'h00
            reg_file[11587] <= 8'h00
            reg_file[11588] <= 8'h00
            reg_file[11589] <= 8'h00
            reg_file[11590] <= 8'h00
            reg_file[11591] <= 8'h00
            reg_file[11592] <= 8'h00
            reg_file[11593] <= 8'h00
            reg_file[11594] <= 8'h00
            reg_file[11595] <= 8'h00
            reg_file[11596] <= 8'h00
            reg_file[11597] <= 8'h00
            reg_file[11598] <= 8'h00
            reg_file[11599] <= 8'h00
            reg_file[11600] <= 8'h00
            reg_file[11601] <= 8'h00
            reg_file[11602] <= 8'h00
            reg_file[11603] <= 8'h00
            reg_file[11604] <= 8'h00
            reg_file[11605] <= 8'h00
            reg_file[11606] <= 8'h00
            reg_file[11607] <= 8'h00
            reg_file[11608] <= 8'h00
            reg_file[11609] <= 8'h00
            reg_file[11610] <= 8'h00
            reg_file[11611] <= 8'h00
            reg_file[11612] <= 8'h00
            reg_file[11613] <= 8'h00
            reg_file[11614] <= 8'h00
            reg_file[11615] <= 8'h00
            reg_file[11616] <= 8'h00
            reg_file[11617] <= 8'h00
            reg_file[11618] <= 8'h00
            reg_file[11619] <= 8'h00
            reg_file[11620] <= 8'h00
            reg_file[11621] <= 8'h00
            reg_file[11622] <= 8'h00
            reg_file[11623] <= 8'h00
            reg_file[11624] <= 8'h00
            reg_file[11625] <= 8'h00
            reg_file[11626] <= 8'h00
            reg_file[11627] <= 8'h00
            reg_file[11628] <= 8'h00
            reg_file[11629] <= 8'h00
            reg_file[11630] <= 8'h00
            reg_file[11631] <= 8'h00
            reg_file[11632] <= 8'h00
            reg_file[11633] <= 8'h00
            reg_file[11634] <= 8'h00
            reg_file[11635] <= 8'h00
            reg_file[11636] <= 8'h00
            reg_file[11637] <= 8'h00
            reg_file[11638] <= 8'h00
            reg_file[11639] <= 8'h00
            reg_file[11640] <= 8'h00
            reg_file[11641] <= 8'h00
            reg_file[11642] <= 8'h00
            reg_file[11643] <= 8'h00
            reg_file[11644] <= 8'h00
            reg_file[11645] <= 8'h00
            reg_file[11646] <= 8'h00
            reg_file[11647] <= 8'h00
            reg_file[11648] <= 8'h00
            reg_file[11649] <= 8'h00
            reg_file[11650] <= 8'h00
            reg_file[11651] <= 8'h00
            reg_file[11652] <= 8'h00
            reg_file[11653] <= 8'h00
            reg_file[11654] <= 8'h00
            reg_file[11655] <= 8'h00
            reg_file[11656] <= 8'h00
            reg_file[11657] <= 8'h00
            reg_file[11658] <= 8'h00
            reg_file[11659] <= 8'h00
            reg_file[11660] <= 8'h00
            reg_file[11661] <= 8'h00
            reg_file[11662] <= 8'h00
            reg_file[11663] <= 8'h00
            reg_file[11664] <= 8'h00
            reg_file[11665] <= 8'h00
            reg_file[11666] <= 8'h00
            reg_file[11667] <= 8'h00
            reg_file[11668] <= 8'h00
            reg_file[11669] <= 8'h00
            reg_file[11670] <= 8'h00
            reg_file[11671] <= 8'h00
            reg_file[11672] <= 8'h00
            reg_file[11673] <= 8'h00
            reg_file[11674] <= 8'h00
            reg_file[11675] <= 8'h00
            reg_file[11676] <= 8'h00
            reg_file[11677] <= 8'h00
            reg_file[11678] <= 8'h00
            reg_file[11679] <= 8'h00
            reg_file[11680] <= 8'h00
            reg_file[11681] <= 8'h00
            reg_file[11682] <= 8'h00
            reg_file[11683] <= 8'h00
            reg_file[11684] <= 8'h00
            reg_file[11685] <= 8'h00
            reg_file[11686] <= 8'h00
            reg_file[11687] <= 8'h00
            reg_file[11688] <= 8'h00
            reg_file[11689] <= 8'h00
            reg_file[11690] <= 8'h00
            reg_file[11691] <= 8'h00
            reg_file[11692] <= 8'h00
            reg_file[11693] <= 8'h00
            reg_file[11694] <= 8'h00
            reg_file[11695] <= 8'h00
            reg_file[11696] <= 8'h00
            reg_file[11697] <= 8'h00
            reg_file[11698] <= 8'h00
            reg_file[11699] <= 8'h00
            reg_file[11700] <= 8'h00
            reg_file[11701] <= 8'h00
            reg_file[11702] <= 8'h00
            reg_file[11703] <= 8'h00
            reg_file[11704] <= 8'h00
            reg_file[11705] <= 8'h00
            reg_file[11706] <= 8'h00
            reg_file[11707] <= 8'h00
            reg_file[11708] <= 8'h00
            reg_file[11709] <= 8'h00
            reg_file[11710] <= 8'h00
            reg_file[11711] <= 8'h00
            reg_file[11712] <= 8'h00
            reg_file[11713] <= 8'h00
            reg_file[11714] <= 8'h00
            reg_file[11715] <= 8'h00
            reg_file[11716] <= 8'h00
            reg_file[11717] <= 8'h00
            reg_file[11718] <= 8'h00
            reg_file[11719] <= 8'h00
            reg_file[11720] <= 8'h00
            reg_file[11721] <= 8'h00
            reg_file[11722] <= 8'h00
            reg_file[11723] <= 8'h00
            reg_file[11724] <= 8'h00
            reg_file[11725] <= 8'h00
            reg_file[11726] <= 8'h00
            reg_file[11727] <= 8'h00
            reg_file[11728] <= 8'h00
            reg_file[11729] <= 8'h00
            reg_file[11730] <= 8'h00
            reg_file[11731] <= 8'h00
            reg_file[11732] <= 8'h00
            reg_file[11733] <= 8'h00
            reg_file[11734] <= 8'h00
            reg_file[11735] <= 8'h00
            reg_file[11736] <= 8'h00
            reg_file[11737] <= 8'h00
            reg_file[11738] <= 8'h00
            reg_file[11739] <= 8'h00
            reg_file[11740] <= 8'h00
            reg_file[11741] <= 8'h00
            reg_file[11742] <= 8'h00
            reg_file[11743] <= 8'h00
            reg_file[11744] <= 8'h00
            reg_file[11745] <= 8'h00
            reg_file[11746] <= 8'h00
            reg_file[11747] <= 8'h00
            reg_file[11748] <= 8'h00
            reg_file[11749] <= 8'h00
            reg_file[11750] <= 8'h00
            reg_file[11751] <= 8'h00
            reg_file[11752] <= 8'h00
            reg_file[11753] <= 8'h00
            reg_file[11754] <= 8'h00
            reg_file[11755] <= 8'h00
            reg_file[11756] <= 8'h00
            reg_file[11757] <= 8'h00
            reg_file[11758] <= 8'h00
            reg_file[11759] <= 8'h00
            reg_file[11760] <= 8'h00
            reg_file[11761] <= 8'h00
            reg_file[11762] <= 8'h00
            reg_file[11763] <= 8'h00
            reg_file[11764] <= 8'h00
            reg_file[11765] <= 8'h00
            reg_file[11766] <= 8'h00
            reg_file[11767] <= 8'h00
            reg_file[11768] <= 8'h00
            reg_file[11769] <= 8'h00
            reg_file[11770] <= 8'h00
            reg_file[11771] <= 8'h00
            reg_file[11772] <= 8'h00
            reg_file[11773] <= 8'h00
            reg_file[11774] <= 8'h00
            reg_file[11775] <= 8'h00
            reg_file[11776] <= 8'h00
            reg_file[11777] <= 8'h00
            reg_file[11778] <= 8'h00
            reg_file[11779] <= 8'h00
            reg_file[11780] <= 8'h00
            reg_file[11781] <= 8'h00
            reg_file[11782] <= 8'h00
            reg_file[11783] <= 8'h00
            reg_file[11784] <= 8'h00
            reg_file[11785] <= 8'h00
            reg_file[11786] <= 8'h00
            reg_file[11787] <= 8'h00
            reg_file[11788] <= 8'h00
            reg_file[11789] <= 8'h00
            reg_file[11790] <= 8'h00
            reg_file[11791] <= 8'h00
            reg_file[11792] <= 8'h00
            reg_file[11793] <= 8'h00
            reg_file[11794] <= 8'h00
            reg_file[11795] <= 8'h00
            reg_file[11796] <= 8'h00
            reg_file[11797] <= 8'h00
            reg_file[11798] <= 8'h00
            reg_file[11799] <= 8'h00
            reg_file[11800] <= 8'h00
            reg_file[11801] <= 8'h00
            reg_file[11802] <= 8'h00
            reg_file[11803] <= 8'h00
            reg_file[11804] <= 8'h00
            reg_file[11805] <= 8'h00
            reg_file[11806] <= 8'h00
            reg_file[11807] <= 8'h00
            reg_file[11808] <= 8'h00
            reg_file[11809] <= 8'h00
            reg_file[11810] <= 8'h00
            reg_file[11811] <= 8'h00
            reg_file[11812] <= 8'h00
            reg_file[11813] <= 8'h00
            reg_file[11814] <= 8'h00
            reg_file[11815] <= 8'h00
            reg_file[11816] <= 8'h00
            reg_file[11817] <= 8'h00
            reg_file[11818] <= 8'h00
            reg_file[11819] <= 8'h00
            reg_file[11820] <= 8'h00
            reg_file[11821] <= 8'h00
            reg_file[11822] <= 8'h00
            reg_file[11823] <= 8'h00
            reg_file[11824] <= 8'h00
            reg_file[11825] <= 8'h00
            reg_file[11826] <= 8'h00
            reg_file[11827] <= 8'h00
            reg_file[11828] <= 8'h00
            reg_file[11829] <= 8'h00
            reg_file[11830] <= 8'h00
            reg_file[11831] <= 8'h00
            reg_file[11832] <= 8'h00
            reg_file[11833] <= 8'h00
            reg_file[11834] <= 8'h00
            reg_file[11835] <= 8'h00
            reg_file[11836] <= 8'h00
            reg_file[11837] <= 8'h00
            reg_file[11838] <= 8'h00
            reg_file[11839] <= 8'h00
            reg_file[11840] <= 8'h00
            reg_file[11841] <= 8'h00
            reg_file[11842] <= 8'h00
            reg_file[11843] <= 8'h00
            reg_file[11844] <= 8'h00
            reg_file[11845] <= 8'h00
            reg_file[11846] <= 8'h00
            reg_file[11847] <= 8'h00
            reg_file[11848] <= 8'h00
            reg_file[11849] <= 8'h00
            reg_file[11850] <= 8'h00
            reg_file[11851] <= 8'h00
            reg_file[11852] <= 8'h00
            reg_file[11853] <= 8'h00
            reg_file[11854] <= 8'h00
            reg_file[11855] <= 8'h00
            reg_file[11856] <= 8'h00
            reg_file[11857] <= 8'h00
            reg_file[11858] <= 8'h00
            reg_file[11859] <= 8'h00
            reg_file[11860] <= 8'h00
            reg_file[11861] <= 8'h00
            reg_file[11862] <= 8'h00
            reg_file[11863] <= 8'h00
            reg_file[11864] <= 8'h00
            reg_file[11865] <= 8'h00
            reg_file[11866] <= 8'h00
            reg_file[11867] <= 8'h00
            reg_file[11868] <= 8'h00
            reg_file[11869] <= 8'h00
            reg_file[11870] <= 8'h00
            reg_file[11871] <= 8'h00
            reg_file[11872] <= 8'h00
            reg_file[11873] <= 8'h00
            reg_file[11874] <= 8'h00
            reg_file[11875] <= 8'h00
            reg_file[11876] <= 8'h00
            reg_file[11877] <= 8'h00
            reg_file[11878] <= 8'h00
            reg_file[11879] <= 8'h00
            reg_file[11880] <= 8'h00
            reg_file[11881] <= 8'h00
            reg_file[11882] <= 8'h00
            reg_file[11883] <= 8'h00
            reg_file[11884] <= 8'h00
            reg_file[11885] <= 8'h00
            reg_file[11886] <= 8'h00
            reg_file[11887] <= 8'h00
            reg_file[11888] <= 8'h00
            reg_file[11889] <= 8'h00
            reg_file[11890] <= 8'h00
            reg_file[11891] <= 8'h00
            reg_file[11892] <= 8'h00
            reg_file[11893] <= 8'h00
            reg_file[11894] <= 8'h00
            reg_file[11895] <= 8'h00
            reg_file[11896] <= 8'h00
            reg_file[11897] <= 8'h00
            reg_file[11898] <= 8'h00
            reg_file[11899] <= 8'h00
            reg_file[11900] <= 8'h00
            reg_file[11901] <= 8'h00
            reg_file[11902] <= 8'h00
            reg_file[11903] <= 8'h00
            reg_file[11904] <= 8'h00
            reg_file[11905] <= 8'h00
            reg_file[11906] <= 8'h00
            reg_file[11907] <= 8'h00
            reg_file[11908] <= 8'h00
            reg_file[11909] <= 8'h00
            reg_file[11910] <= 8'h00
            reg_file[11911] <= 8'h00
            reg_file[11912] <= 8'h00
            reg_file[11913] <= 8'h00
            reg_file[11914] <= 8'h00
            reg_file[11915] <= 8'h00
            reg_file[11916] <= 8'h00
            reg_file[11917] <= 8'h00
            reg_file[11918] <= 8'h00
            reg_file[11919] <= 8'h00
            reg_file[11920] <= 8'h00
            reg_file[11921] <= 8'h00
            reg_file[11922] <= 8'h00
            reg_file[11923] <= 8'h00
            reg_file[11924] <= 8'h00
            reg_file[11925] <= 8'h00
            reg_file[11926] <= 8'h00
            reg_file[11927] <= 8'h00
            reg_file[11928] <= 8'h00
            reg_file[11929] <= 8'h00
            reg_file[11930] <= 8'h00
            reg_file[11931] <= 8'h00
            reg_file[11932] <= 8'h00
            reg_file[11933] <= 8'h00
            reg_file[11934] <= 8'h00
            reg_file[11935] <= 8'h00
            reg_file[11936] <= 8'h00
            reg_file[11937] <= 8'h00
            reg_file[11938] <= 8'h00
            reg_file[11939] <= 8'h00
            reg_file[11940] <= 8'h00
            reg_file[11941] <= 8'h00
            reg_file[11942] <= 8'h00
            reg_file[11943] <= 8'h00
            reg_file[11944] <= 8'h00
            reg_file[11945] <= 8'h00
            reg_file[11946] <= 8'h00
            reg_file[11947] <= 8'h00
            reg_file[11948] <= 8'h00
            reg_file[11949] <= 8'h00
            reg_file[11950] <= 8'h00
            reg_file[11951] <= 8'h00
            reg_file[11952] <= 8'h00
            reg_file[11953] <= 8'h00
            reg_file[11954] <= 8'h00
            reg_file[11955] <= 8'h00
            reg_file[11956] <= 8'h00
            reg_file[11957] <= 8'h00
            reg_file[11958] <= 8'h00
            reg_file[11959] <= 8'h00
            reg_file[11960] <= 8'h00
            reg_file[11961] <= 8'h00
            reg_file[11962] <= 8'h00
            reg_file[11963] <= 8'h00
            reg_file[11964] <= 8'h00
            reg_file[11965] <= 8'h00
            reg_file[11966] <= 8'h00
            reg_file[11967] <= 8'h00
            reg_file[11968] <= 8'h00
            reg_file[11969] <= 8'h00
            reg_file[11970] <= 8'h00
            reg_file[11971] <= 8'h00
            reg_file[11972] <= 8'h00
            reg_file[11973] <= 8'h00
            reg_file[11974] <= 8'h00
            reg_file[11975] <= 8'h00
            reg_file[11976] <= 8'h00
            reg_file[11977] <= 8'h00
            reg_file[11978] <= 8'h00
            reg_file[11979] <= 8'h00
            reg_file[11980] <= 8'h00
            reg_file[11981] <= 8'h00
            reg_file[11982] <= 8'h00
            reg_file[11983] <= 8'h00
            reg_file[11984] <= 8'h00
            reg_file[11985] <= 8'h00
            reg_file[11986] <= 8'h00
            reg_file[11987] <= 8'h00
            reg_file[11988] <= 8'h00
            reg_file[11989] <= 8'h00
            reg_file[11990] <= 8'h00
            reg_file[11991] <= 8'h00
            reg_file[11992] <= 8'h00
            reg_file[11993] <= 8'h00
            reg_file[11994] <= 8'h00
            reg_file[11995] <= 8'h00
            reg_file[11996] <= 8'h00
            reg_file[11997] <= 8'h00
            reg_file[11998] <= 8'h00
            reg_file[11999] <= 8'h00
            reg_file[12000] <= 8'h00
            reg_file[12001] <= 8'h00
            reg_file[12002] <= 8'h00
            reg_file[12003] <= 8'h00
            reg_file[12004] <= 8'h00
            reg_file[12005] <= 8'h00
            reg_file[12006] <= 8'h00
            reg_file[12007] <= 8'h00
            reg_file[12008] <= 8'h00
            reg_file[12009] <= 8'h00
            reg_file[12010] <= 8'h00
            reg_file[12011] <= 8'h00
            reg_file[12012] <= 8'h00
            reg_file[12013] <= 8'h00
            reg_file[12014] <= 8'h00
            reg_file[12015] <= 8'h00
            reg_file[12016] <= 8'h00
            reg_file[12017] <= 8'h00
            reg_file[12018] <= 8'h00
            reg_file[12019] <= 8'h00
            reg_file[12020] <= 8'h00
            reg_file[12021] <= 8'h00
            reg_file[12022] <= 8'h00
            reg_file[12023] <= 8'h00
            reg_file[12024] <= 8'h00
            reg_file[12025] <= 8'h00
            reg_file[12026] <= 8'h00
            reg_file[12027] <= 8'h00
            reg_file[12028] <= 8'h00
            reg_file[12029] <= 8'h00
            reg_file[12030] <= 8'h00
            reg_file[12031] <= 8'h00
            reg_file[12032] <= 8'h00
            reg_file[12033] <= 8'h00
            reg_file[12034] <= 8'h00
            reg_file[12035] <= 8'h00
            reg_file[12036] <= 8'h00
            reg_file[12037] <= 8'h00
            reg_file[12038] <= 8'h00
            reg_file[12039] <= 8'h00
            reg_file[12040] <= 8'h00
            reg_file[12041] <= 8'h00
            reg_file[12042] <= 8'h00
            reg_file[12043] <= 8'h00
            reg_file[12044] <= 8'h00
            reg_file[12045] <= 8'h00
            reg_file[12046] <= 8'h00
            reg_file[12047] <= 8'h00
            reg_file[12048] <= 8'h00
            reg_file[12049] <= 8'h00
            reg_file[12050] <= 8'h00
            reg_file[12051] <= 8'h00
            reg_file[12052] <= 8'h00
            reg_file[12053] <= 8'h00
            reg_file[12054] <= 8'h00
            reg_file[12055] <= 8'h00
            reg_file[12056] <= 8'h00
            reg_file[12057] <= 8'h00
            reg_file[12058] <= 8'h00
            reg_file[12059] <= 8'h00
            reg_file[12060] <= 8'h00
            reg_file[12061] <= 8'h00
            reg_file[12062] <= 8'h00
            reg_file[12063] <= 8'h00
            reg_file[12064] <= 8'h00
            reg_file[12065] <= 8'h00
            reg_file[12066] <= 8'h00
            reg_file[12067] <= 8'h00
            reg_file[12068] <= 8'h00
            reg_file[12069] <= 8'h00
            reg_file[12070] <= 8'h00
            reg_file[12071] <= 8'h00
            reg_file[12072] <= 8'h00
            reg_file[12073] <= 8'h00
            reg_file[12074] <= 8'h00
            reg_file[12075] <= 8'h00
            reg_file[12076] <= 8'h00
            reg_file[12077] <= 8'h00
            reg_file[12078] <= 8'h00
            reg_file[12079] <= 8'h00
            reg_file[12080] <= 8'h00
            reg_file[12081] <= 8'h00
            reg_file[12082] <= 8'h00
            reg_file[12083] <= 8'h00
            reg_file[12084] <= 8'h00
            reg_file[12085] <= 8'h00
            reg_file[12086] <= 8'h00
            reg_file[12087] <= 8'h00
            reg_file[12088] <= 8'h00
            reg_file[12089] <= 8'h00
            reg_file[12090] <= 8'h00
            reg_file[12091] <= 8'h00
            reg_file[12092] <= 8'h00
            reg_file[12093] <= 8'h00
            reg_file[12094] <= 8'h00
            reg_file[12095] <= 8'h00
            reg_file[12096] <= 8'h00
            reg_file[12097] <= 8'h00
            reg_file[12098] <= 8'h00
            reg_file[12099] <= 8'h00
            reg_file[12100] <= 8'h00
            reg_file[12101] <= 8'h00
            reg_file[12102] <= 8'h00
            reg_file[12103] <= 8'h00
            reg_file[12104] <= 8'h00
            reg_file[12105] <= 8'h00
            reg_file[12106] <= 8'h00
            reg_file[12107] <= 8'h00
            reg_file[12108] <= 8'h00
            reg_file[12109] <= 8'h00
            reg_file[12110] <= 8'h00
            reg_file[12111] <= 8'h00
            reg_file[12112] <= 8'h00
            reg_file[12113] <= 8'h00
            reg_file[12114] <= 8'h00
            reg_file[12115] <= 8'h00
            reg_file[12116] <= 8'h00
            reg_file[12117] <= 8'h00
            reg_file[12118] <= 8'h00
            reg_file[12119] <= 8'h00
            reg_file[12120] <= 8'h00
            reg_file[12121] <= 8'h00
            reg_file[12122] <= 8'h00
            reg_file[12123] <= 8'h00
            reg_file[12124] <= 8'h00
            reg_file[12125] <= 8'h00
            reg_file[12126] <= 8'h00
            reg_file[12127] <= 8'h00
            reg_file[12128] <= 8'h00
            reg_file[12129] <= 8'h00
            reg_file[12130] <= 8'h00
            reg_file[12131] <= 8'h00
            reg_file[12132] <= 8'h00
            reg_file[12133] <= 8'h00
            reg_file[12134] <= 8'h00
            reg_file[12135] <= 8'h00
            reg_file[12136] <= 8'h00
            reg_file[12137] <= 8'h00
            reg_file[12138] <= 8'h00
            reg_file[12139] <= 8'h00
            reg_file[12140] <= 8'h00
            reg_file[12141] <= 8'h00
            reg_file[12142] <= 8'h00
            reg_file[12143] <= 8'h00
            reg_file[12144] <= 8'h00
            reg_file[12145] <= 8'h00
            reg_file[12146] <= 8'h00
            reg_file[12147] <= 8'h00
            reg_file[12148] <= 8'h00
            reg_file[12149] <= 8'h00
            reg_file[12150] <= 8'h00
            reg_file[12151] <= 8'h00
            reg_file[12152] <= 8'h00
            reg_file[12153] <= 8'h00
            reg_file[12154] <= 8'h00
            reg_file[12155] <= 8'h00
            reg_file[12156] <= 8'h00
            reg_file[12157] <= 8'h00
            reg_file[12158] <= 8'h00
            reg_file[12159] <= 8'h00
            reg_file[12160] <= 8'h00
            reg_file[12161] <= 8'h00
            reg_file[12162] <= 8'h00
            reg_file[12163] <= 8'h00
            reg_file[12164] <= 8'h00
            reg_file[12165] <= 8'h00
            reg_file[12166] <= 8'h00
            reg_file[12167] <= 8'h00
            reg_file[12168] <= 8'h00
            reg_file[12169] <= 8'h00
            reg_file[12170] <= 8'h00
            reg_file[12171] <= 8'h00
            reg_file[12172] <= 8'h00
            reg_file[12173] <= 8'h00
            reg_file[12174] <= 8'h00
            reg_file[12175] <= 8'h00
            reg_file[12176] <= 8'h00
            reg_file[12177] <= 8'h00
            reg_file[12178] <= 8'h00
            reg_file[12179] <= 8'h00
            reg_file[12180] <= 8'h00
            reg_file[12181] <= 8'h00
            reg_file[12182] <= 8'h00
            reg_file[12183] <= 8'h00
            reg_file[12184] <= 8'h00
            reg_file[12185] <= 8'h00
            reg_file[12186] <= 8'h00
            reg_file[12187] <= 8'h00
            reg_file[12188] <= 8'h00
            reg_file[12189] <= 8'h00
            reg_file[12190] <= 8'h00
            reg_file[12191] <= 8'h00
            reg_file[12192] <= 8'h00
            reg_file[12193] <= 8'h00
            reg_file[12194] <= 8'h00
            reg_file[12195] <= 8'h00
            reg_file[12196] <= 8'h00
            reg_file[12197] <= 8'h00
            reg_file[12198] <= 8'h00
            reg_file[12199] <= 8'h00
            reg_file[12200] <= 8'h00
            reg_file[12201] <= 8'h00
            reg_file[12202] <= 8'h00
            reg_file[12203] <= 8'h00
            reg_file[12204] <= 8'h00
            reg_file[12205] <= 8'h00
            reg_file[12206] <= 8'h00
            reg_file[12207] <= 8'h00
            reg_file[12208] <= 8'h00
            reg_file[12209] <= 8'h00
            reg_file[12210] <= 8'h00
            reg_file[12211] <= 8'h00
            reg_file[12212] <= 8'h00
            reg_file[12213] <= 8'h00
            reg_file[12214] <= 8'h00
            reg_file[12215] <= 8'h00
            reg_file[12216] <= 8'h00
            reg_file[12217] <= 8'h00
            reg_file[12218] <= 8'h00
            reg_file[12219] <= 8'h00
            reg_file[12220] <= 8'h00
            reg_file[12221] <= 8'h00
            reg_file[12222] <= 8'h00
            reg_file[12223] <= 8'h00
            reg_file[12224] <= 8'h00
            reg_file[12225] <= 8'h00
            reg_file[12226] <= 8'h00
            reg_file[12227] <= 8'h00
            reg_file[12228] <= 8'h00
            reg_file[12229] <= 8'h00
            reg_file[12230] <= 8'h00
            reg_file[12231] <= 8'h00
            reg_file[12232] <= 8'h00
            reg_file[12233] <= 8'h00
            reg_file[12234] <= 8'h00
            reg_file[12235] <= 8'h00
            reg_file[12236] <= 8'h00
            reg_file[12237] <= 8'h00
            reg_file[12238] <= 8'h00
            reg_file[12239] <= 8'h00
            reg_file[12240] <= 8'h00
            reg_file[12241] <= 8'h00
            reg_file[12242] <= 8'h00
            reg_file[12243] <= 8'h00
            reg_file[12244] <= 8'h00
            reg_file[12245] <= 8'h00
            reg_file[12246] <= 8'h00
            reg_file[12247] <= 8'h00
            reg_file[12248] <= 8'h00
            reg_file[12249] <= 8'h00
            reg_file[12250] <= 8'h00
            reg_file[12251] <= 8'h00
            reg_file[12252] <= 8'h00
            reg_file[12253] <= 8'h00
            reg_file[12254] <= 8'h00
            reg_file[12255] <= 8'h00
            reg_file[12256] <= 8'h00
            reg_file[12257] <= 8'h00
            reg_file[12258] <= 8'h00
            reg_file[12259] <= 8'h00
            reg_file[12260] <= 8'h00
            reg_file[12261] <= 8'h00
            reg_file[12262] <= 8'h00
            reg_file[12263] <= 8'h00
            reg_file[12264] <= 8'h00
            reg_file[12265] <= 8'h00
            reg_file[12266] <= 8'h00
            reg_file[12267] <= 8'h00
            reg_file[12268] <= 8'h00
            reg_file[12269] <= 8'h00
            reg_file[12270] <= 8'h00
            reg_file[12271] <= 8'h00
            reg_file[12272] <= 8'h00
            reg_file[12273] <= 8'h00
            reg_file[12274] <= 8'h00
            reg_file[12275] <= 8'h00
            reg_file[12276] <= 8'h00
            reg_file[12277] <= 8'h00
            reg_file[12278] <= 8'h00
            reg_file[12279] <= 8'h00
            reg_file[12280] <= 8'h00
            reg_file[12281] <= 8'h00
            reg_file[12282] <= 8'h00
            reg_file[12283] <= 8'h00
            reg_file[12284] <= 8'h00
            reg_file[12285] <= 8'h00
            reg_file[12286] <= 8'h00
            reg_file[12287] <= 8'h00
            reg_file[12288] <= 8'h00
            reg_file[12289] <= 8'h00
            reg_file[12290] <= 8'h00
            reg_file[12291] <= 8'h00
            reg_file[12292] <= 8'h00
            reg_file[12293] <= 8'h00
            reg_file[12294] <= 8'h00
            reg_file[12295] <= 8'h00
            reg_file[12296] <= 8'h00
            reg_file[12297] <= 8'h00
            reg_file[12298] <= 8'h00
            reg_file[12299] <= 8'h00
            reg_file[12300] <= 8'h00
            reg_file[12301] <= 8'h00
            reg_file[12302] <= 8'h00
            reg_file[12303] <= 8'h00
            reg_file[12304] <= 8'h00
            reg_file[12305] <= 8'h00
            reg_file[12306] <= 8'h00
            reg_file[12307] <= 8'h00
            reg_file[12308] <= 8'h00
            reg_file[12309] <= 8'h00
            reg_file[12310] <= 8'h00
            reg_file[12311] <= 8'h00
            reg_file[12312] <= 8'h00
            reg_file[12313] <= 8'h00
            reg_file[12314] <= 8'h00
            reg_file[12315] <= 8'h00
            reg_file[12316] <= 8'h00
            reg_file[12317] <= 8'h00
            reg_file[12318] <= 8'h00
            reg_file[12319] <= 8'h00
            reg_file[12320] <= 8'h00
            reg_file[12321] <= 8'h00
            reg_file[12322] <= 8'h00
            reg_file[12323] <= 8'h00
            reg_file[12324] <= 8'h00
            reg_file[12325] <= 8'h00
            reg_file[12326] <= 8'h00
            reg_file[12327] <= 8'h00
            reg_file[12328] <= 8'h00
            reg_file[12329] <= 8'h00
            reg_file[12330] <= 8'h00
            reg_file[12331] <= 8'h00
            reg_file[12332] <= 8'h00
            reg_file[12333] <= 8'h00
            reg_file[12334] <= 8'h00
            reg_file[12335] <= 8'h00
            reg_file[12336] <= 8'h00
            reg_file[12337] <= 8'h00
            reg_file[12338] <= 8'h00
            reg_file[12339] <= 8'h00
            reg_file[12340] <= 8'h00
            reg_file[12341] <= 8'h00
            reg_file[12342] <= 8'h00
            reg_file[12343] <= 8'h00
            reg_file[12344] <= 8'h00
            reg_file[12345] <= 8'h00
            reg_file[12346] <= 8'h00
            reg_file[12347] <= 8'h00
            reg_file[12348] <= 8'h00
            reg_file[12349] <= 8'h00
            reg_file[12350] <= 8'h00
            reg_file[12351] <= 8'h00
            reg_file[12352] <= 8'h00
            reg_file[12353] <= 8'h00
            reg_file[12354] <= 8'h00
            reg_file[12355] <= 8'h00
            reg_file[12356] <= 8'h00
            reg_file[12357] <= 8'h00
            reg_file[12358] <= 8'h00
            reg_file[12359] <= 8'h00
            reg_file[12360] <= 8'h00
            reg_file[12361] <= 8'h00
            reg_file[12362] <= 8'h00
            reg_file[12363] <= 8'h00
            reg_file[12364] <= 8'h00
            reg_file[12365] <= 8'h00
            reg_file[12366] <= 8'h00
            reg_file[12367] <= 8'h00
            reg_file[12368] <= 8'h00
            reg_file[12369] <= 8'h00
            reg_file[12370] <= 8'h00
            reg_file[12371] <= 8'h00
            reg_file[12372] <= 8'h00
            reg_file[12373] <= 8'h00
            reg_file[12374] <= 8'h00
            reg_file[12375] <= 8'h00
            reg_file[12376] <= 8'h00
            reg_file[12377] <= 8'h00
            reg_file[12378] <= 8'h00
            reg_file[12379] <= 8'h00
            reg_file[12380] <= 8'h00
            reg_file[12381] <= 8'h00
            reg_file[12382] <= 8'h00
            reg_file[12383] <= 8'h00
            reg_file[12384] <= 8'h00
            reg_file[12385] <= 8'h00
            reg_file[12386] <= 8'h00
            reg_file[12387] <= 8'h00
            reg_file[12388] <= 8'h00
            reg_file[12389] <= 8'h00
            reg_file[12390] <= 8'h00
            reg_file[12391] <= 8'h00
            reg_file[12392] <= 8'h00
            reg_file[12393] <= 8'h00
            reg_file[12394] <= 8'h00
            reg_file[12395] <= 8'h00
            reg_file[12396] <= 8'h00
            reg_file[12397] <= 8'h00
            reg_file[12398] <= 8'h00
            reg_file[12399] <= 8'h00
            reg_file[12400] <= 8'h00
            reg_file[12401] <= 8'h00
            reg_file[12402] <= 8'h00
            reg_file[12403] <= 8'h00
            reg_file[12404] <= 8'h00
            reg_file[12405] <= 8'h00
            reg_file[12406] <= 8'h00
            reg_file[12407] <= 8'h00
            reg_file[12408] <= 8'h00
            reg_file[12409] <= 8'h00
            reg_file[12410] <= 8'h00
            reg_file[12411] <= 8'h00
            reg_file[12412] <= 8'h00
            reg_file[12413] <= 8'h00
            reg_file[12414] <= 8'h00
            reg_file[12415] <= 8'h00
            reg_file[12416] <= 8'h00
            reg_file[12417] <= 8'h00
            reg_file[12418] <= 8'h00
            reg_file[12419] <= 8'h00
            reg_file[12420] <= 8'h00
            reg_file[12421] <= 8'h00
            reg_file[12422] <= 8'h00
            reg_file[12423] <= 8'h00
            reg_file[12424] <= 8'h00
            reg_file[12425] <= 8'h00
            reg_file[12426] <= 8'h00
            reg_file[12427] <= 8'h00
            reg_file[12428] <= 8'h00
            reg_file[12429] <= 8'h00
            reg_file[12430] <= 8'h00
            reg_file[12431] <= 8'h00
            reg_file[12432] <= 8'h00
            reg_file[12433] <= 8'h00
            reg_file[12434] <= 8'h00
            reg_file[12435] <= 8'h00
            reg_file[12436] <= 8'h00
            reg_file[12437] <= 8'h00
            reg_file[12438] <= 8'h00
            reg_file[12439] <= 8'h00
            reg_file[12440] <= 8'h00
            reg_file[12441] <= 8'h00
            reg_file[12442] <= 8'h00
            reg_file[12443] <= 8'h00
            reg_file[12444] <= 8'h00
            reg_file[12445] <= 8'h00
            reg_file[12446] <= 8'h00
            reg_file[12447] <= 8'h00
            reg_file[12448] <= 8'h00
            reg_file[12449] <= 8'h00
            reg_file[12450] <= 8'h00
            reg_file[12451] <= 8'h00
            reg_file[12452] <= 8'h00
            reg_file[12453] <= 8'h00
            reg_file[12454] <= 8'h00
            reg_file[12455] <= 8'h00
            reg_file[12456] <= 8'h00
            reg_file[12457] <= 8'h00
            reg_file[12458] <= 8'h00
            reg_file[12459] <= 8'h00
            reg_file[12460] <= 8'h00
            reg_file[12461] <= 8'h00
            reg_file[12462] <= 8'h00
            reg_file[12463] <= 8'h00
            reg_file[12464] <= 8'h00
            reg_file[12465] <= 8'h00
            reg_file[12466] <= 8'h00
            reg_file[12467] <= 8'h00
            reg_file[12468] <= 8'h00
            reg_file[12469] <= 8'h00
            reg_file[12470] <= 8'h00
            reg_file[12471] <= 8'h00
            reg_file[12472] <= 8'h00
            reg_file[12473] <= 8'h00
            reg_file[12474] <= 8'h00
            reg_file[12475] <= 8'h00
            reg_file[12476] <= 8'h00
            reg_file[12477] <= 8'h00
            reg_file[12478] <= 8'h00
            reg_file[12479] <= 8'h00
            reg_file[12480] <= 8'h00
            reg_file[12481] <= 8'h00
            reg_file[12482] <= 8'h00
            reg_file[12483] <= 8'h00
            reg_file[12484] <= 8'h00
            reg_file[12485] <= 8'h00
            reg_file[12486] <= 8'h00
            reg_file[12487] <= 8'h00
            reg_file[12488] <= 8'h00
            reg_file[12489] <= 8'h00
            reg_file[12490] <= 8'h00
            reg_file[12491] <= 8'h00
            reg_file[12492] <= 8'h00
            reg_file[12493] <= 8'h00
            reg_file[12494] <= 8'h00
            reg_file[12495] <= 8'h00
            reg_file[12496] <= 8'h00
            reg_file[12497] <= 8'h00
            reg_file[12498] <= 8'h00
            reg_file[12499] <= 8'h00
            reg_file[12500] <= 8'h00
            reg_file[12501] <= 8'h00
            reg_file[12502] <= 8'h00
            reg_file[12503] <= 8'h00
            reg_file[12504] <= 8'h00
            reg_file[12505] <= 8'h00
            reg_file[12506] <= 8'h00
            reg_file[12507] <= 8'h00
            reg_file[12508] <= 8'h00
            reg_file[12509] <= 8'h00
            reg_file[12510] <= 8'h00
            reg_file[12511] <= 8'h00
            reg_file[12512] <= 8'h00
            reg_file[12513] <= 8'h00
            reg_file[12514] <= 8'h00
            reg_file[12515] <= 8'h00
            reg_file[12516] <= 8'h00
            reg_file[12517] <= 8'h00
            reg_file[12518] <= 8'h00
            reg_file[12519] <= 8'h00
            reg_file[12520] <= 8'h00
            reg_file[12521] <= 8'h00
            reg_file[12522] <= 8'h00
            reg_file[12523] <= 8'h00
            reg_file[12524] <= 8'h00
            reg_file[12525] <= 8'h00
            reg_file[12526] <= 8'h00
            reg_file[12527] <= 8'h00
            reg_file[12528] <= 8'h00
            reg_file[12529] <= 8'h00
            reg_file[12530] <= 8'h00
            reg_file[12531] <= 8'h00
            reg_file[12532] <= 8'h00
            reg_file[12533] <= 8'h00
            reg_file[12534] <= 8'h00
            reg_file[12535] <= 8'h00
            reg_file[12536] <= 8'h00
            reg_file[12537] <= 8'h00
            reg_file[12538] <= 8'h00
            reg_file[12539] <= 8'h00
            reg_file[12540] <= 8'h00
            reg_file[12541] <= 8'h00
            reg_file[12542] <= 8'h00
            reg_file[12543] <= 8'h00
            reg_file[12544] <= 8'h00
            reg_file[12545] <= 8'h00
            reg_file[12546] <= 8'h00
            reg_file[12547] <= 8'h00
            reg_file[12548] <= 8'h00
            reg_file[12549] <= 8'h00
            reg_file[12550] <= 8'h00
            reg_file[12551] <= 8'h00
            reg_file[12552] <= 8'h00
            reg_file[12553] <= 8'h00
            reg_file[12554] <= 8'h00
            reg_file[12555] <= 8'h00
            reg_file[12556] <= 8'h00
            reg_file[12557] <= 8'h00
            reg_file[12558] <= 8'h00
            reg_file[12559] <= 8'h00
            reg_file[12560] <= 8'h00
            reg_file[12561] <= 8'h00
            reg_file[12562] <= 8'h00
            reg_file[12563] <= 8'h00
            reg_file[12564] <= 8'h00
            reg_file[12565] <= 8'h00
            reg_file[12566] <= 8'h00
            reg_file[12567] <= 8'h00
            reg_file[12568] <= 8'h00
            reg_file[12569] <= 8'h00
            reg_file[12570] <= 8'h00
            reg_file[12571] <= 8'h00
            reg_file[12572] <= 8'h00
            reg_file[12573] <= 8'h00
            reg_file[12574] <= 8'h00
            reg_file[12575] <= 8'h00
            reg_file[12576] <= 8'h00
            reg_file[12577] <= 8'h00
            reg_file[12578] <= 8'h00
            reg_file[12579] <= 8'h00
            reg_file[12580] <= 8'h00
            reg_file[12581] <= 8'h00
            reg_file[12582] <= 8'h00
            reg_file[12583] <= 8'h00
            reg_file[12584] <= 8'h00
            reg_file[12585] <= 8'h00
            reg_file[12586] <= 8'h00
            reg_file[12587] <= 8'h00
            reg_file[12588] <= 8'h00
            reg_file[12589] <= 8'h00
            reg_file[12590] <= 8'h00
            reg_file[12591] <= 8'h00
            reg_file[12592] <= 8'h00
            reg_file[12593] <= 8'h00
            reg_file[12594] <= 8'h00
            reg_file[12595] <= 8'h00
            reg_file[12596] <= 8'h00
            reg_file[12597] <= 8'h00
            reg_file[12598] <= 8'h00
            reg_file[12599] <= 8'h00
            reg_file[12600] <= 8'h00
            reg_file[12601] <= 8'h00
            reg_file[12602] <= 8'h00
            reg_file[12603] <= 8'h00
            reg_file[12604] <= 8'h00
            reg_file[12605] <= 8'h00
            reg_file[12606] <= 8'h00
            reg_file[12607] <= 8'h00
            reg_file[12608] <= 8'h00
            reg_file[12609] <= 8'h00
            reg_file[12610] <= 8'h00
            reg_file[12611] <= 8'h00
            reg_file[12612] <= 8'h00
            reg_file[12613] <= 8'h00
            reg_file[12614] <= 8'h00
            reg_file[12615] <= 8'h00
            reg_file[12616] <= 8'h00
            reg_file[12617] <= 8'h00
            reg_file[12618] <= 8'h00
            reg_file[12619] <= 8'h00
            reg_file[12620] <= 8'h00
            reg_file[12621] <= 8'h00
            reg_file[12622] <= 8'h00
            reg_file[12623] <= 8'h00
            reg_file[12624] <= 8'h00
            reg_file[12625] <= 8'h00
            reg_file[12626] <= 8'h00
            reg_file[12627] <= 8'h00
            reg_file[12628] <= 8'h00
            reg_file[12629] <= 8'h00
            reg_file[12630] <= 8'h00
            reg_file[12631] <= 8'h00
            reg_file[12632] <= 8'h00
            reg_file[12633] <= 8'h00
            reg_file[12634] <= 8'h00
            reg_file[12635] <= 8'h00
            reg_file[12636] <= 8'h00
            reg_file[12637] <= 8'h00
            reg_file[12638] <= 8'h00
            reg_file[12639] <= 8'h00
            reg_file[12640] <= 8'h00
            reg_file[12641] <= 8'h00
            reg_file[12642] <= 8'h00
            reg_file[12643] <= 8'h00
            reg_file[12644] <= 8'h00
            reg_file[12645] <= 8'h00
            reg_file[12646] <= 8'h00
            reg_file[12647] <= 8'h00
            reg_file[12648] <= 8'h00
            reg_file[12649] <= 8'h00
            reg_file[12650] <= 8'h00
            reg_file[12651] <= 8'h00
            reg_file[12652] <= 8'h00
            reg_file[12653] <= 8'h00
            reg_file[12654] <= 8'h00
            reg_file[12655] <= 8'h00
            reg_file[12656] <= 8'h00
            reg_file[12657] <= 8'h00
            reg_file[12658] <= 8'h00
            reg_file[12659] <= 8'h00
            reg_file[12660] <= 8'h00
            reg_file[12661] <= 8'h00
            reg_file[12662] <= 8'h00
            reg_file[12663] <= 8'h00
            reg_file[12664] <= 8'h00
            reg_file[12665] <= 8'h00
            reg_file[12666] <= 8'h00
            reg_file[12667] <= 8'h00
            reg_file[12668] <= 8'h00
            reg_file[12669] <= 8'h00
            reg_file[12670] <= 8'h00
            reg_file[12671] <= 8'h00
            reg_file[12672] <= 8'h00
            reg_file[12673] <= 8'h00
            reg_file[12674] <= 8'h00
            reg_file[12675] <= 8'h00
            reg_file[12676] <= 8'h00
            reg_file[12677] <= 8'h00
            reg_file[12678] <= 8'h00
            reg_file[12679] <= 8'h00
            reg_file[12680] <= 8'h00
            reg_file[12681] <= 8'h00
            reg_file[12682] <= 8'h00
            reg_file[12683] <= 8'h00
            reg_file[12684] <= 8'h00
            reg_file[12685] <= 8'h00
            reg_file[12686] <= 8'h00
            reg_file[12687] <= 8'h00
            reg_file[12688] <= 8'h00
            reg_file[12689] <= 8'h00
            reg_file[12690] <= 8'h00
            reg_file[12691] <= 8'h00
            reg_file[12692] <= 8'h00
            reg_file[12693] <= 8'h00
            reg_file[12694] <= 8'h00
            reg_file[12695] <= 8'h00
            reg_file[12696] <= 8'h00
            reg_file[12697] <= 8'h00
            reg_file[12698] <= 8'h00
            reg_file[12699] <= 8'h00
            reg_file[12700] <= 8'h00
            reg_file[12701] <= 8'h00
            reg_file[12702] <= 8'h00
            reg_file[12703] <= 8'h00
            reg_file[12704] <= 8'h00
            reg_file[12705] <= 8'h00
            reg_file[12706] <= 8'h00
            reg_file[12707] <= 8'h00
            reg_file[12708] <= 8'h00
            reg_file[12709] <= 8'h00
            reg_file[12710] <= 8'h00
            reg_file[12711] <= 8'h00
            reg_file[12712] <= 8'h00
            reg_file[12713] <= 8'h00
            reg_file[12714] <= 8'h00
            reg_file[12715] <= 8'h00
            reg_file[12716] <= 8'h00
            reg_file[12717] <= 8'h00
            reg_file[12718] <= 8'h00
            reg_file[12719] <= 8'h00
            reg_file[12720] <= 8'h00
            reg_file[12721] <= 8'h00
            reg_file[12722] <= 8'h00
            reg_file[12723] <= 8'h00
            reg_file[12724] <= 8'h00
            reg_file[12725] <= 8'h00
            reg_file[12726] <= 8'h00
            reg_file[12727] <= 8'h00
            reg_file[12728] <= 8'h00
            reg_file[12729] <= 8'h00
            reg_file[12730] <= 8'h00
            reg_file[12731] <= 8'h00
            reg_file[12732] <= 8'h00
            reg_file[12733] <= 8'h00
            reg_file[12734] <= 8'h00
            reg_file[12735] <= 8'h00
            reg_file[12736] <= 8'h00
            reg_file[12737] <= 8'h00
            reg_file[12738] <= 8'h00
            reg_file[12739] <= 8'h00
            reg_file[12740] <= 8'h00
            reg_file[12741] <= 8'h00
            reg_file[12742] <= 8'h00
            reg_file[12743] <= 8'h00
            reg_file[12744] <= 8'h00
            reg_file[12745] <= 8'h00
            reg_file[12746] <= 8'h00
            reg_file[12747] <= 8'h00
            reg_file[12748] <= 8'h00
            reg_file[12749] <= 8'h00
            reg_file[12750] <= 8'h00
            reg_file[12751] <= 8'h00
            reg_file[12752] <= 8'h00
            reg_file[12753] <= 8'h00
            reg_file[12754] <= 8'h00
            reg_file[12755] <= 8'h00
            reg_file[12756] <= 8'h00
            reg_file[12757] <= 8'h00
            reg_file[12758] <= 8'h00
            reg_file[12759] <= 8'h00
            reg_file[12760] <= 8'h00
            reg_file[12761] <= 8'h00
            reg_file[12762] <= 8'h00
            reg_file[12763] <= 8'h00
            reg_file[12764] <= 8'h00
            reg_file[12765] <= 8'h00
            reg_file[12766] <= 8'h00
            reg_file[12767] <= 8'h00
            reg_file[12768] <= 8'h00
            reg_file[12769] <= 8'h00
            reg_file[12770] <= 8'h00
            reg_file[12771] <= 8'h00
            reg_file[12772] <= 8'h00
            reg_file[12773] <= 8'h00
            reg_file[12774] <= 8'h00
            reg_file[12775] <= 8'h00
            reg_file[12776] <= 8'h00
            reg_file[12777] <= 8'h00
            reg_file[12778] <= 8'h00
            reg_file[12779] <= 8'h00
            reg_file[12780] <= 8'h00
            reg_file[12781] <= 8'h00
            reg_file[12782] <= 8'h00
            reg_file[12783] <= 8'h00
            reg_file[12784] <= 8'h00
            reg_file[12785] <= 8'h00
            reg_file[12786] <= 8'h00
            reg_file[12787] <= 8'h00
            reg_file[12788] <= 8'h00
            reg_file[12789] <= 8'h00
            reg_file[12790] <= 8'h00
            reg_file[12791] <= 8'h00
            reg_file[12792] <= 8'h00
            reg_file[12793] <= 8'h00
            reg_file[12794] <= 8'h00
            reg_file[12795] <= 8'h00
            reg_file[12796] <= 8'h00
            reg_file[12797] <= 8'h00
            reg_file[12798] <= 8'h00
            reg_file[12799] <= 8'h00
            reg_file[12800] <= 8'h00
            reg_file[12801] <= 8'h00
            reg_file[12802] <= 8'h00
            reg_file[12803] <= 8'h00
            reg_file[12804] <= 8'h00
            reg_file[12805] <= 8'h00
            reg_file[12806] <= 8'h00
            reg_file[12807] <= 8'h00
            reg_file[12808] <= 8'h00
            reg_file[12809] <= 8'h00
            reg_file[12810] <= 8'h00
            reg_file[12811] <= 8'h00
            reg_file[12812] <= 8'h00
            reg_file[12813] <= 8'h00
            reg_file[12814] <= 8'h00
            reg_file[12815] <= 8'h00
            reg_file[12816] <= 8'h00
            reg_file[12817] <= 8'h00
            reg_file[12818] <= 8'h00
            reg_file[12819] <= 8'h00
            reg_file[12820] <= 8'h00
            reg_file[12821] <= 8'h00
            reg_file[12822] <= 8'h00
            reg_file[12823] <= 8'h00
            reg_file[12824] <= 8'h00
            reg_file[12825] <= 8'h00
            reg_file[12826] <= 8'h00
            reg_file[12827] <= 8'h00
            reg_file[12828] <= 8'h00
            reg_file[12829] <= 8'h00
            reg_file[12830] <= 8'h00
            reg_file[12831] <= 8'h00
            reg_file[12832] <= 8'h00
            reg_file[12833] <= 8'h00
            reg_file[12834] <= 8'h00
            reg_file[12835] <= 8'h00
            reg_file[12836] <= 8'h00
            reg_file[12837] <= 8'h00
            reg_file[12838] <= 8'h00
            reg_file[12839] <= 8'h00
            reg_file[12840] <= 8'h00
            reg_file[12841] <= 8'h00
            reg_file[12842] <= 8'h00
            reg_file[12843] <= 8'h00
            reg_file[12844] <= 8'h00
            reg_file[12845] <= 8'h00
            reg_file[12846] <= 8'h00
            reg_file[12847] <= 8'h00
            reg_file[12848] <= 8'h00
            reg_file[12849] <= 8'h00
            reg_file[12850] <= 8'h00
            reg_file[12851] <= 8'h00
            reg_file[12852] <= 8'h00
            reg_file[12853] <= 8'h00
            reg_file[12854] <= 8'h00
            reg_file[12855] <= 8'h00
            reg_file[12856] <= 8'h00
            reg_file[12857] <= 8'h00
            reg_file[12858] <= 8'h00
            reg_file[12859] <= 8'h00
            reg_file[12860] <= 8'h00
            reg_file[12861] <= 8'h00
            reg_file[12862] <= 8'h00
            reg_file[12863] <= 8'h00
            reg_file[12864] <= 8'h00
            reg_file[12865] <= 8'h00
            reg_file[12866] <= 8'h00
            reg_file[12867] <= 8'h00
            reg_file[12868] <= 8'h00
            reg_file[12869] <= 8'h00
            reg_file[12870] <= 8'h00
            reg_file[12871] <= 8'h00
            reg_file[12872] <= 8'h00
            reg_file[12873] <= 8'h00
            reg_file[12874] <= 8'h00
            reg_file[12875] <= 8'h00
            reg_file[12876] <= 8'h00
            reg_file[12877] <= 8'h00
            reg_file[12878] <= 8'h00
            reg_file[12879] <= 8'h00
            reg_file[12880] <= 8'h00
            reg_file[12881] <= 8'h00
            reg_file[12882] <= 8'h00
            reg_file[12883] <= 8'h00
            reg_file[12884] <= 8'h00
            reg_file[12885] <= 8'h00
            reg_file[12886] <= 8'h00
            reg_file[12887] <= 8'h00
            reg_file[12888] <= 8'h00
            reg_file[12889] <= 8'h00
            reg_file[12890] <= 8'h00
            reg_file[12891] <= 8'h00
            reg_file[12892] <= 8'h00
            reg_file[12893] <= 8'h00
            reg_file[12894] <= 8'h00
            reg_file[12895] <= 8'h00
            reg_file[12896] <= 8'h00
            reg_file[12897] <= 8'h00
            reg_file[12898] <= 8'h00
            reg_file[12899] <= 8'h00
            reg_file[12900] <= 8'h00
            reg_file[12901] <= 8'h00
            reg_file[12902] <= 8'h00
            reg_file[12903] <= 8'h00
            reg_file[12904] <= 8'h00
            reg_file[12905] <= 8'h00
            reg_file[12906] <= 8'h00
            reg_file[12907] <= 8'h00
            reg_file[12908] <= 8'h00
            reg_file[12909] <= 8'h00
            reg_file[12910] <= 8'h00
            reg_file[12911] <= 8'h00
            reg_file[12912] <= 8'h00
            reg_file[12913] <= 8'h00
            reg_file[12914] <= 8'h00
            reg_file[12915] <= 8'h00
            reg_file[12916] <= 8'h00
            reg_file[12917] <= 8'h00
            reg_file[12918] <= 8'h00
            reg_file[12919] <= 8'h00
            reg_file[12920] <= 8'h00
            reg_file[12921] <= 8'h00
            reg_file[12922] <= 8'h00
            reg_file[12923] <= 8'h00
            reg_file[12924] <= 8'h00
            reg_file[12925] <= 8'h00
            reg_file[12926] <= 8'h00
            reg_file[12927] <= 8'h00
            reg_file[12928] <= 8'h00
            reg_file[12929] <= 8'h00
            reg_file[12930] <= 8'h00
            reg_file[12931] <= 8'h00
            reg_file[12932] <= 8'h00
            reg_file[12933] <= 8'h00
            reg_file[12934] <= 8'h00
            reg_file[12935] <= 8'h00
            reg_file[12936] <= 8'h00
            reg_file[12937] <= 8'h00
            reg_file[12938] <= 8'h00
            reg_file[12939] <= 8'h00
            reg_file[12940] <= 8'h00
            reg_file[12941] <= 8'h00
            reg_file[12942] <= 8'h00
            reg_file[12943] <= 8'h00
            reg_file[12944] <= 8'h00
            reg_file[12945] <= 8'h00
            reg_file[12946] <= 8'h00
            reg_file[12947] <= 8'h00
            reg_file[12948] <= 8'h00
            reg_file[12949] <= 8'h00
            reg_file[12950] <= 8'h00
            reg_file[12951] <= 8'h00
            reg_file[12952] <= 8'h00
            reg_file[12953] <= 8'h00
            reg_file[12954] <= 8'h00
            reg_file[12955] <= 8'h00
            reg_file[12956] <= 8'h00
            reg_file[12957] <= 8'h00
            reg_file[12958] <= 8'h00
            reg_file[12959] <= 8'h00
            reg_file[12960] <= 8'h00
            reg_file[12961] <= 8'h00
            reg_file[12962] <= 8'h00
            reg_file[12963] <= 8'h00
            reg_file[12964] <= 8'h00
            reg_file[12965] <= 8'h00
            reg_file[12966] <= 8'h00
            reg_file[12967] <= 8'h00
            reg_file[12968] <= 8'h00
            reg_file[12969] <= 8'h00
            reg_file[12970] <= 8'h00
            reg_file[12971] <= 8'h00
            reg_file[12972] <= 8'h00
            reg_file[12973] <= 8'h00
            reg_file[12974] <= 8'h00
            reg_file[12975] <= 8'h00
            reg_file[12976] <= 8'h00
            reg_file[12977] <= 8'h00
            reg_file[12978] <= 8'h00
            reg_file[12979] <= 8'h00
            reg_file[12980] <= 8'h00
            reg_file[12981] <= 8'h00
            reg_file[12982] <= 8'h00
            reg_file[12983] <= 8'h00
            reg_file[12984] <= 8'h00
            reg_file[12985] <= 8'h00
            reg_file[12986] <= 8'h00
            reg_file[12987] <= 8'h00
            reg_file[12988] <= 8'h00
            reg_file[12989] <= 8'h00
            reg_file[12990] <= 8'h00
            reg_file[12991] <= 8'h00
            reg_file[12992] <= 8'h00
            reg_file[12993] <= 8'h00
            reg_file[12994] <= 8'h00
            reg_file[12995] <= 8'h00
            reg_file[12996] <= 8'h00
            reg_file[12997] <= 8'h00
            reg_file[12998] <= 8'h00
            reg_file[12999] <= 8'h00
            reg_file[13000] <= 8'h00
            reg_file[13001] <= 8'h00
            reg_file[13002] <= 8'h00
            reg_file[13003] <= 8'h00
            reg_file[13004] <= 8'h00
            reg_file[13005] <= 8'h00
            reg_file[13006] <= 8'h00
            reg_file[13007] <= 8'h00
            reg_file[13008] <= 8'h00
            reg_file[13009] <= 8'h00
            reg_file[13010] <= 8'h00
            reg_file[13011] <= 8'h00
            reg_file[13012] <= 8'h00
            reg_file[13013] <= 8'h00
            reg_file[13014] <= 8'h00
            reg_file[13015] <= 8'h00
            reg_file[13016] <= 8'h00
            reg_file[13017] <= 8'h00
            reg_file[13018] <= 8'h00
            reg_file[13019] <= 8'h00
            reg_file[13020] <= 8'h00
            reg_file[13021] <= 8'h00
            reg_file[13022] <= 8'h00
            reg_file[13023] <= 8'h00
            reg_file[13024] <= 8'h00
            reg_file[13025] <= 8'h00
            reg_file[13026] <= 8'h00
            reg_file[13027] <= 8'h00
            reg_file[13028] <= 8'h00
            reg_file[13029] <= 8'h00
            reg_file[13030] <= 8'h00
            reg_file[13031] <= 8'h00
            reg_file[13032] <= 8'h00
            reg_file[13033] <= 8'h00
            reg_file[13034] <= 8'h00
            reg_file[13035] <= 8'h00
            reg_file[13036] <= 8'h00
            reg_file[13037] <= 8'h00
            reg_file[13038] <= 8'h00
            reg_file[13039] <= 8'h00
            reg_file[13040] <= 8'h00
            reg_file[13041] <= 8'h00
            reg_file[13042] <= 8'h00
            reg_file[13043] <= 8'h00
            reg_file[13044] <= 8'h00
            reg_file[13045] <= 8'h00
            reg_file[13046] <= 8'h00
            reg_file[13047] <= 8'h00
            reg_file[13048] <= 8'h00
            reg_file[13049] <= 8'h00
            reg_file[13050] <= 8'h00
            reg_file[13051] <= 8'h00
            reg_file[13052] <= 8'h00
            reg_file[13053] <= 8'h00
            reg_file[13054] <= 8'h00
            reg_file[13055] <= 8'h00
            reg_file[13056] <= 8'h00
            reg_file[13057] <= 8'h00
            reg_file[13058] <= 8'h00
            reg_file[13059] <= 8'h00
            reg_file[13060] <= 8'h00
            reg_file[13061] <= 8'h00
            reg_file[13062] <= 8'h00
            reg_file[13063] <= 8'h00
            reg_file[13064] <= 8'h00
            reg_file[13065] <= 8'h00
            reg_file[13066] <= 8'h00
            reg_file[13067] <= 8'h00
            reg_file[13068] <= 8'h00
            reg_file[13069] <= 8'h00
            reg_file[13070] <= 8'h00
            reg_file[13071] <= 8'h00
            reg_file[13072] <= 8'h00
            reg_file[13073] <= 8'h00
            reg_file[13074] <= 8'h00
            reg_file[13075] <= 8'h00
            reg_file[13076] <= 8'h00
            reg_file[13077] <= 8'h00
            reg_file[13078] <= 8'h00
            reg_file[13079] <= 8'h00
            reg_file[13080] <= 8'h00
            reg_file[13081] <= 8'h00
            reg_file[13082] <= 8'h00
            reg_file[13083] <= 8'h00
            reg_file[13084] <= 8'h00
            reg_file[13085] <= 8'h00
            reg_file[13086] <= 8'h00
            reg_file[13087] <= 8'h00
            reg_file[13088] <= 8'h00
            reg_file[13089] <= 8'h00
            reg_file[13090] <= 8'h00
            reg_file[13091] <= 8'h00
            reg_file[13092] <= 8'h00
            reg_file[13093] <= 8'h00
            reg_file[13094] <= 8'h00
            reg_file[13095] <= 8'h00
            reg_file[13096] <= 8'h00
            reg_file[13097] <= 8'h00
            reg_file[13098] <= 8'h00
            reg_file[13099] <= 8'h00
            reg_file[13100] <= 8'h00
            reg_file[13101] <= 8'h00
            reg_file[13102] <= 8'h00
            reg_file[13103] <= 8'h00
            reg_file[13104] <= 8'h00
            reg_file[13105] <= 8'h00
            reg_file[13106] <= 8'h00
            reg_file[13107] <= 8'h00
            reg_file[13108] <= 8'h00
            reg_file[13109] <= 8'h00
            reg_file[13110] <= 8'h00
            reg_file[13111] <= 8'h00
            reg_file[13112] <= 8'h00
            reg_file[13113] <= 8'h00
            reg_file[13114] <= 8'h00
            reg_file[13115] <= 8'h00
            reg_file[13116] <= 8'h00
            reg_file[13117] <= 8'h00
            reg_file[13118] <= 8'h00
            reg_file[13119] <= 8'h00
            reg_file[13120] <= 8'h00
            reg_file[13121] <= 8'h00
            reg_file[13122] <= 8'h00
            reg_file[13123] <= 8'h00
            reg_file[13124] <= 8'h00
            reg_file[13125] <= 8'h00
            reg_file[13126] <= 8'h00
            reg_file[13127] <= 8'h00
            reg_file[13128] <= 8'h00
            reg_file[13129] <= 8'h00
            reg_file[13130] <= 8'h00
            reg_file[13131] <= 8'h00
            reg_file[13132] <= 8'h00
            reg_file[13133] <= 8'h00
            reg_file[13134] <= 8'h00
            reg_file[13135] <= 8'h00
            reg_file[13136] <= 8'h00
            reg_file[13137] <= 8'h00
            reg_file[13138] <= 8'h00
            reg_file[13139] <= 8'h00
            reg_file[13140] <= 8'h00
            reg_file[13141] <= 8'h00
            reg_file[13142] <= 8'h00
            reg_file[13143] <= 8'h00
            reg_file[13144] <= 8'h00
            reg_file[13145] <= 8'h00
            reg_file[13146] <= 8'h00
            reg_file[13147] <= 8'h00
            reg_file[13148] <= 8'h00
            reg_file[13149] <= 8'h00
            reg_file[13150] <= 8'h00
            reg_file[13151] <= 8'h00
            reg_file[13152] <= 8'h00
            reg_file[13153] <= 8'h00
            reg_file[13154] <= 8'h00
            reg_file[13155] <= 8'h00
            reg_file[13156] <= 8'h00
            reg_file[13157] <= 8'h00
            reg_file[13158] <= 8'h00
            reg_file[13159] <= 8'h00
            reg_file[13160] <= 8'h00
            reg_file[13161] <= 8'h00
            reg_file[13162] <= 8'h00
            reg_file[13163] <= 8'h00
            reg_file[13164] <= 8'h00
            reg_file[13165] <= 8'h00
            reg_file[13166] <= 8'h00
            reg_file[13167] <= 8'h00
            reg_file[13168] <= 8'h00
            reg_file[13169] <= 8'h00
            reg_file[13170] <= 8'h00
            reg_file[13171] <= 8'h00
            reg_file[13172] <= 8'h00
            reg_file[13173] <= 8'h00
            reg_file[13174] <= 8'h00
            reg_file[13175] <= 8'h00
            reg_file[13176] <= 8'h00
            reg_file[13177] <= 8'h00
            reg_file[13178] <= 8'h00
            reg_file[13179] <= 8'h00
            reg_file[13180] <= 8'h00
            reg_file[13181] <= 8'h00
            reg_file[13182] <= 8'h00
            reg_file[13183] <= 8'h00
            reg_file[13184] <= 8'h00
            reg_file[13185] <= 8'h00
            reg_file[13186] <= 8'h00
            reg_file[13187] <= 8'h00
            reg_file[13188] <= 8'h00
            reg_file[13189] <= 8'h00
            reg_file[13190] <= 8'h00
            reg_file[13191] <= 8'h00
            reg_file[13192] <= 8'h00
            reg_file[13193] <= 8'h00
            reg_file[13194] <= 8'h00
            reg_file[13195] <= 8'h00
            reg_file[13196] <= 8'h00
            reg_file[13197] <= 8'h00
            reg_file[13198] <= 8'h00
            reg_file[13199] <= 8'h00
            reg_file[13200] <= 8'h00
            reg_file[13201] <= 8'h00
            reg_file[13202] <= 8'h00
            reg_file[13203] <= 8'h00
            reg_file[13204] <= 8'h00
            reg_file[13205] <= 8'h00
            reg_file[13206] <= 8'h00
            reg_file[13207] <= 8'h00
            reg_file[13208] <= 8'h00
            reg_file[13209] <= 8'h00
            reg_file[13210] <= 8'h00
            reg_file[13211] <= 8'h00
            reg_file[13212] <= 8'h00
            reg_file[13213] <= 8'h00
            reg_file[13214] <= 8'h00
            reg_file[13215] <= 8'h00
            reg_file[13216] <= 8'h00
            reg_file[13217] <= 8'h00
            reg_file[13218] <= 8'h00
            reg_file[13219] <= 8'h00
            reg_file[13220] <= 8'h00
            reg_file[13221] <= 8'h00
            reg_file[13222] <= 8'h00
            reg_file[13223] <= 8'h00
            reg_file[13224] <= 8'h00
            reg_file[13225] <= 8'h00
            reg_file[13226] <= 8'h00
            reg_file[13227] <= 8'h00
            reg_file[13228] <= 8'h00
            reg_file[13229] <= 8'h00
            reg_file[13230] <= 8'h00
            reg_file[13231] <= 8'h00
            reg_file[13232] <= 8'h00
            reg_file[13233] <= 8'h00
            reg_file[13234] <= 8'h00
            reg_file[13235] <= 8'h00
            reg_file[13236] <= 8'h00
            reg_file[13237] <= 8'h00
            reg_file[13238] <= 8'h00
            reg_file[13239] <= 8'h00
            reg_file[13240] <= 8'h00
            reg_file[13241] <= 8'h00
            reg_file[13242] <= 8'h00
            reg_file[13243] <= 8'h00
            reg_file[13244] <= 8'h00
            reg_file[13245] <= 8'h00
            reg_file[13246] <= 8'h00
            reg_file[13247] <= 8'h00
            reg_file[13248] <= 8'h00
            reg_file[13249] <= 8'h00
            reg_file[13250] <= 8'h00
            reg_file[13251] <= 8'h00
            reg_file[13252] <= 8'h00
            reg_file[13253] <= 8'h00
            reg_file[13254] <= 8'h00
            reg_file[13255] <= 8'h00
            reg_file[13256] <= 8'h00
            reg_file[13257] <= 8'h00
            reg_file[13258] <= 8'h00
            reg_file[13259] <= 8'h00
            reg_file[13260] <= 8'h00
            reg_file[13261] <= 8'h00
            reg_file[13262] <= 8'h00
            reg_file[13263] <= 8'h00
            reg_file[13264] <= 8'h00
            reg_file[13265] <= 8'h00
            reg_file[13266] <= 8'h00
            reg_file[13267] <= 8'h00
            reg_file[13268] <= 8'h00
            reg_file[13269] <= 8'h00
            reg_file[13270] <= 8'h00
            reg_file[13271] <= 8'h00
            reg_file[13272] <= 8'h00
            reg_file[13273] <= 8'h00
            reg_file[13274] <= 8'h00
            reg_file[13275] <= 8'h00
            reg_file[13276] <= 8'h00
            reg_file[13277] <= 8'h00
            reg_file[13278] <= 8'h00
            reg_file[13279] <= 8'h00
            reg_file[13280] <= 8'h00
            reg_file[13281] <= 8'h00
            reg_file[13282] <= 8'h00
            reg_file[13283] <= 8'h00
            reg_file[13284] <= 8'h00
            reg_file[13285] <= 8'h00
            reg_file[13286] <= 8'h00
            reg_file[13287] <= 8'h00
            reg_file[13288] <= 8'h00
            reg_file[13289] <= 8'h00
            reg_file[13290] <= 8'h00
            reg_file[13291] <= 8'h00
            reg_file[13292] <= 8'h00
            reg_file[13293] <= 8'h00
            reg_file[13294] <= 8'h00
            reg_file[13295] <= 8'h00
            reg_file[13296] <= 8'h00
            reg_file[13297] <= 8'h00
            reg_file[13298] <= 8'h00
            reg_file[13299] <= 8'h00
            reg_file[13300] <= 8'h00
            reg_file[13301] <= 8'h00
            reg_file[13302] <= 8'h00
            reg_file[13303] <= 8'h00
            reg_file[13304] <= 8'h00
            reg_file[13305] <= 8'h00
            reg_file[13306] <= 8'h00
            reg_file[13307] <= 8'h00
            reg_file[13308] <= 8'h00
            reg_file[13309] <= 8'h00
            reg_file[13310] <= 8'h00
            reg_file[13311] <= 8'h00
            reg_file[13312] <= 8'h00
            reg_file[13313] <= 8'h00
            reg_file[13314] <= 8'h00
            reg_file[13315] <= 8'h00
            reg_file[13316] <= 8'h00
            reg_file[13317] <= 8'h00
            reg_file[13318] <= 8'h00
            reg_file[13319] <= 8'h00
            reg_file[13320] <= 8'h00
            reg_file[13321] <= 8'h00
            reg_file[13322] <= 8'h00
            reg_file[13323] <= 8'h00
            reg_file[13324] <= 8'h00
            reg_file[13325] <= 8'h00
            reg_file[13326] <= 8'h00
            reg_file[13327] <= 8'h00
            reg_file[13328] <= 8'h00
            reg_file[13329] <= 8'h00
            reg_file[13330] <= 8'h00
            reg_file[13331] <= 8'h00
            reg_file[13332] <= 8'h00
            reg_file[13333] <= 8'h00
            reg_file[13334] <= 8'h00
            reg_file[13335] <= 8'h00
            reg_file[13336] <= 8'h00
            reg_file[13337] <= 8'h00
            reg_file[13338] <= 8'h00
            reg_file[13339] <= 8'h00
            reg_file[13340] <= 8'h00
            reg_file[13341] <= 8'h00
            reg_file[13342] <= 8'h00
            reg_file[13343] <= 8'h00
            reg_file[13344] <= 8'h00
            reg_file[13345] <= 8'h00
            reg_file[13346] <= 8'h00
            reg_file[13347] <= 8'h00
            reg_file[13348] <= 8'h00
            reg_file[13349] <= 8'h00
            reg_file[13350] <= 8'h00
            reg_file[13351] <= 8'h00
            reg_file[13352] <= 8'h00
            reg_file[13353] <= 8'h00
            reg_file[13354] <= 8'h00
            reg_file[13355] <= 8'h00
            reg_file[13356] <= 8'h00
            reg_file[13357] <= 8'h00
            reg_file[13358] <= 8'h00
            reg_file[13359] <= 8'h00
            reg_file[13360] <= 8'h00
            reg_file[13361] <= 8'h00
            reg_file[13362] <= 8'h00
            reg_file[13363] <= 8'h00
            reg_file[13364] <= 8'h00
            reg_file[13365] <= 8'h00
            reg_file[13366] <= 8'h00
            reg_file[13367] <= 8'h00
            reg_file[13368] <= 8'h00
            reg_file[13369] <= 8'h00
            reg_file[13370] <= 8'h00
            reg_file[13371] <= 8'h00
            reg_file[13372] <= 8'h00
            reg_file[13373] <= 8'h00
            reg_file[13374] <= 8'h00
            reg_file[13375] <= 8'h00
            reg_file[13376] <= 8'h00
            reg_file[13377] <= 8'h00
            reg_file[13378] <= 8'h00
            reg_file[13379] <= 8'h00
            reg_file[13380] <= 8'h00
            reg_file[13381] <= 8'h00
            reg_file[13382] <= 8'h00
            reg_file[13383] <= 8'h00
            reg_file[13384] <= 8'h00
            reg_file[13385] <= 8'h00
            reg_file[13386] <= 8'h00
            reg_file[13387] <= 8'h00
            reg_file[13388] <= 8'h00
            reg_file[13389] <= 8'h00
            reg_file[13390] <= 8'h00
            reg_file[13391] <= 8'h00
            reg_file[13392] <= 8'h00
            reg_file[13393] <= 8'h00
            reg_file[13394] <= 8'h00
            reg_file[13395] <= 8'h00
            reg_file[13396] <= 8'h00
            reg_file[13397] <= 8'h00
            reg_file[13398] <= 8'h00
            reg_file[13399] <= 8'h00
            reg_file[13400] <= 8'h00
            reg_file[13401] <= 8'h00
            reg_file[13402] <= 8'h00
            reg_file[13403] <= 8'h00
            reg_file[13404] <= 8'h00
            reg_file[13405] <= 8'h00
            reg_file[13406] <= 8'h00
            reg_file[13407] <= 8'h00
            reg_file[13408] <= 8'h00
            reg_file[13409] <= 8'h00
            reg_file[13410] <= 8'h00
            reg_file[13411] <= 8'h00
            reg_file[13412] <= 8'h00
            reg_file[13413] <= 8'h00
            reg_file[13414] <= 8'h00
            reg_file[13415] <= 8'h00
            reg_file[13416] <= 8'h00
            reg_file[13417] <= 8'h00
            reg_file[13418] <= 8'h00
            reg_file[13419] <= 8'h00
            reg_file[13420] <= 8'h00
            reg_file[13421] <= 8'h00
            reg_file[13422] <= 8'h00
            reg_file[13423] <= 8'h00
            reg_file[13424] <= 8'h00
            reg_file[13425] <= 8'h00
            reg_file[13426] <= 8'h00
            reg_file[13427] <= 8'h00
            reg_file[13428] <= 8'h00
            reg_file[13429] <= 8'h00
            reg_file[13430] <= 8'h00
            reg_file[13431] <= 8'h00
            reg_file[13432] <= 8'h00
            reg_file[13433] <= 8'h00
            reg_file[13434] <= 8'h00
            reg_file[13435] <= 8'h00
            reg_file[13436] <= 8'h00
            reg_file[13437] <= 8'h00
            reg_file[13438] <= 8'h00
            reg_file[13439] <= 8'h00
            reg_file[13440] <= 8'h00
            reg_file[13441] <= 8'h00
            reg_file[13442] <= 8'h00
            reg_file[13443] <= 8'h00
            reg_file[13444] <= 8'h00
            reg_file[13445] <= 8'h00
            reg_file[13446] <= 8'h00
            reg_file[13447] <= 8'h00
            reg_file[13448] <= 8'h00
            reg_file[13449] <= 8'h00
            reg_file[13450] <= 8'h00
            reg_file[13451] <= 8'h00
            reg_file[13452] <= 8'h00
            reg_file[13453] <= 8'h00
            reg_file[13454] <= 8'h00
            reg_file[13455] <= 8'h00
            reg_file[13456] <= 8'h00
            reg_file[13457] <= 8'h00
            reg_file[13458] <= 8'h00
            reg_file[13459] <= 8'h00
            reg_file[13460] <= 8'h00
            reg_file[13461] <= 8'h00
            reg_file[13462] <= 8'h00
            reg_file[13463] <= 8'h00
            reg_file[13464] <= 8'h00
            reg_file[13465] <= 8'h00
            reg_file[13466] <= 8'h00
            reg_file[13467] <= 8'h00
            reg_file[13468] <= 8'h00
            reg_file[13469] <= 8'h00
            reg_file[13470] <= 8'h00
            reg_file[13471] <= 8'h00
            reg_file[13472] <= 8'h00
            reg_file[13473] <= 8'h00
            reg_file[13474] <= 8'h00
            reg_file[13475] <= 8'h00
            reg_file[13476] <= 8'h00
            reg_file[13477] <= 8'h00
            reg_file[13478] <= 8'h00
            reg_file[13479] <= 8'h00
            reg_file[13480] <= 8'h00
            reg_file[13481] <= 8'h00
            reg_file[13482] <= 8'h00
            reg_file[13483] <= 8'h00
            reg_file[13484] <= 8'h00
            reg_file[13485] <= 8'h00
            reg_file[13486] <= 8'h00
            reg_file[13487] <= 8'h00
            reg_file[13488] <= 8'h00
            reg_file[13489] <= 8'h00
            reg_file[13490] <= 8'h00
            reg_file[13491] <= 8'h00
            reg_file[13492] <= 8'h00
            reg_file[13493] <= 8'h00
            reg_file[13494] <= 8'h00
            reg_file[13495] <= 8'h00
            reg_file[13496] <= 8'h00
            reg_file[13497] <= 8'h00
            reg_file[13498] <= 8'h00
            reg_file[13499] <= 8'h00
            reg_file[13500] <= 8'h00
            reg_file[13501] <= 8'h00
            reg_file[13502] <= 8'h00
            reg_file[13503] <= 8'h00
            reg_file[13504] <= 8'h00
            reg_file[13505] <= 8'h00
            reg_file[13506] <= 8'h00
            reg_file[13507] <= 8'h00
            reg_file[13508] <= 8'h00
            reg_file[13509] <= 8'h00
            reg_file[13510] <= 8'h00
            reg_file[13511] <= 8'h00
            reg_file[13512] <= 8'h00
            reg_file[13513] <= 8'h00
            reg_file[13514] <= 8'h00
            reg_file[13515] <= 8'h00
            reg_file[13516] <= 8'h00
            reg_file[13517] <= 8'h00
            reg_file[13518] <= 8'h00
            reg_file[13519] <= 8'h00
            reg_file[13520] <= 8'h00
            reg_file[13521] <= 8'h00
            reg_file[13522] <= 8'h00
            reg_file[13523] <= 8'h00
            reg_file[13524] <= 8'h00
            reg_file[13525] <= 8'h00
            reg_file[13526] <= 8'h00
            reg_file[13527] <= 8'h00
            reg_file[13528] <= 8'h00
            reg_file[13529] <= 8'h00
            reg_file[13530] <= 8'h00
            reg_file[13531] <= 8'h00
            reg_file[13532] <= 8'h00
            reg_file[13533] <= 8'h00
            reg_file[13534] <= 8'h00
            reg_file[13535] <= 8'h00
            reg_file[13536] <= 8'h00
            reg_file[13537] <= 8'h00
            reg_file[13538] <= 8'h00
            reg_file[13539] <= 8'h00
            reg_file[13540] <= 8'h00
            reg_file[13541] <= 8'h00
            reg_file[13542] <= 8'h00
            reg_file[13543] <= 8'h00
            reg_file[13544] <= 8'h00
            reg_file[13545] <= 8'h00
            reg_file[13546] <= 8'h00
            reg_file[13547] <= 8'h00
            reg_file[13548] <= 8'h00
            reg_file[13549] <= 8'h00
            reg_file[13550] <= 8'h00
            reg_file[13551] <= 8'h00
            reg_file[13552] <= 8'h00
            reg_file[13553] <= 8'h00
            reg_file[13554] <= 8'h00
            reg_file[13555] <= 8'h00
            reg_file[13556] <= 8'h00
            reg_file[13557] <= 8'h00
            reg_file[13558] <= 8'h00
            reg_file[13559] <= 8'h00
            reg_file[13560] <= 8'h00
            reg_file[13561] <= 8'h00
            reg_file[13562] <= 8'h00
            reg_file[13563] <= 8'h00
            reg_file[13564] <= 8'h00
            reg_file[13565] <= 8'h00
            reg_file[13566] <= 8'h00
            reg_file[13567] <= 8'h00
            reg_file[13568] <= 8'h00
            reg_file[13569] <= 8'h00
            reg_file[13570] <= 8'h00
            reg_file[13571] <= 8'h00
            reg_file[13572] <= 8'h00
            reg_file[13573] <= 8'h00
            reg_file[13574] <= 8'h00
            reg_file[13575] <= 8'h00
            reg_file[13576] <= 8'h00
            reg_file[13577] <= 8'h00
            reg_file[13578] <= 8'h00
            reg_file[13579] <= 8'h00
            reg_file[13580] <= 8'h00
            reg_file[13581] <= 8'h00
            reg_file[13582] <= 8'h00
            reg_file[13583] <= 8'h00
            reg_file[13584] <= 8'h00
            reg_file[13585] <= 8'h00
            reg_file[13586] <= 8'h00
            reg_file[13587] <= 8'h00
            reg_file[13588] <= 8'h00
            reg_file[13589] <= 8'h00
            reg_file[13590] <= 8'h00
            reg_file[13591] <= 8'h00
            reg_file[13592] <= 8'h00
            reg_file[13593] <= 8'h00
            reg_file[13594] <= 8'h00
            reg_file[13595] <= 8'h00
            reg_file[13596] <= 8'h00
            reg_file[13597] <= 8'h00
            reg_file[13598] <= 8'h00
            reg_file[13599] <= 8'h00
            reg_file[13600] <= 8'h00
            reg_file[13601] <= 8'h00
            reg_file[13602] <= 8'h00
            reg_file[13603] <= 8'h00
            reg_file[13604] <= 8'h00
            reg_file[13605] <= 8'h00
            reg_file[13606] <= 8'h00
            reg_file[13607] <= 8'h00
            reg_file[13608] <= 8'h00
            reg_file[13609] <= 8'h00
            reg_file[13610] <= 8'h00
            reg_file[13611] <= 8'h00
            reg_file[13612] <= 8'h00
            reg_file[13613] <= 8'h00
            reg_file[13614] <= 8'h00
            reg_file[13615] <= 8'h00
            reg_file[13616] <= 8'h00
            reg_file[13617] <= 8'h00
            reg_file[13618] <= 8'h00
            reg_file[13619] <= 8'h00
            reg_file[13620] <= 8'h00
            reg_file[13621] <= 8'h00
            reg_file[13622] <= 8'h00
            reg_file[13623] <= 8'h00
            reg_file[13624] <= 8'h00
            reg_file[13625] <= 8'h00
            reg_file[13626] <= 8'h00
            reg_file[13627] <= 8'h00
            reg_file[13628] <= 8'h00
            reg_file[13629] <= 8'h00
            reg_file[13630] <= 8'h00
            reg_file[13631] <= 8'h00
            reg_file[13632] <= 8'h00
            reg_file[13633] <= 8'h00
            reg_file[13634] <= 8'h00
            reg_file[13635] <= 8'h00
            reg_file[13636] <= 8'h00
            reg_file[13637] <= 8'h00
            reg_file[13638] <= 8'h00
            reg_file[13639] <= 8'h00
            reg_file[13640] <= 8'h00
            reg_file[13641] <= 8'h00
            reg_file[13642] <= 8'h00
            reg_file[13643] <= 8'h00
            reg_file[13644] <= 8'h00
            reg_file[13645] <= 8'h00
            reg_file[13646] <= 8'h00
            reg_file[13647] <= 8'h00
            reg_file[13648] <= 8'h00
            reg_file[13649] <= 8'h00
            reg_file[13650] <= 8'h00
            reg_file[13651] <= 8'h00
            reg_file[13652] <= 8'h00
            reg_file[13653] <= 8'h00
            reg_file[13654] <= 8'h00
            reg_file[13655] <= 8'h00
            reg_file[13656] <= 8'h00
            reg_file[13657] <= 8'h00
            reg_file[13658] <= 8'h00
            reg_file[13659] <= 8'h00
            reg_file[13660] <= 8'h00
            reg_file[13661] <= 8'h00
            reg_file[13662] <= 8'h00
            reg_file[13663] <= 8'h00
            reg_file[13664] <= 8'h00
            reg_file[13665] <= 8'h00
            reg_file[13666] <= 8'h00
            reg_file[13667] <= 8'h00
            reg_file[13668] <= 8'h00
            reg_file[13669] <= 8'h00
            reg_file[13670] <= 8'h00
            reg_file[13671] <= 8'h00
            reg_file[13672] <= 8'h00
            reg_file[13673] <= 8'h00
            reg_file[13674] <= 8'h00
            reg_file[13675] <= 8'h00
            reg_file[13676] <= 8'h00
            reg_file[13677] <= 8'h00
            reg_file[13678] <= 8'h00
            reg_file[13679] <= 8'h00
            reg_file[13680] <= 8'h00
            reg_file[13681] <= 8'h00
            reg_file[13682] <= 8'h00
            reg_file[13683] <= 8'h00
            reg_file[13684] <= 8'h00
            reg_file[13685] <= 8'h00
            reg_file[13686] <= 8'h00
            reg_file[13687] <= 8'h00
            reg_file[13688] <= 8'h00
            reg_file[13689] <= 8'h00
            reg_file[13690] <= 8'h00
            reg_file[13691] <= 8'h00
            reg_file[13692] <= 8'h00
            reg_file[13693] <= 8'h00
            reg_file[13694] <= 8'h00
            reg_file[13695] <= 8'h00
            reg_file[13696] <= 8'h00
            reg_file[13697] <= 8'h00
            reg_file[13698] <= 8'h00
            reg_file[13699] <= 8'h00
            reg_file[13700] <= 8'h00
            reg_file[13701] <= 8'h00
            reg_file[13702] <= 8'h00
            reg_file[13703] <= 8'h00
            reg_file[13704] <= 8'h00
            reg_file[13705] <= 8'h00
            reg_file[13706] <= 8'h00
            reg_file[13707] <= 8'h00
            reg_file[13708] <= 8'h00
            reg_file[13709] <= 8'h00
            reg_file[13710] <= 8'h00
            reg_file[13711] <= 8'h00
            reg_file[13712] <= 8'h00
            reg_file[13713] <= 8'h00
            reg_file[13714] <= 8'h00
            reg_file[13715] <= 8'h00
            reg_file[13716] <= 8'h00
            reg_file[13717] <= 8'h00
            reg_file[13718] <= 8'h00
            reg_file[13719] <= 8'h00
            reg_file[13720] <= 8'h00
            reg_file[13721] <= 8'h00
            reg_file[13722] <= 8'h00
            reg_file[13723] <= 8'h00
            reg_file[13724] <= 8'h00
            reg_file[13725] <= 8'h00
            reg_file[13726] <= 8'h00
            reg_file[13727] <= 8'h00
            reg_file[13728] <= 8'h00
            reg_file[13729] <= 8'h00
            reg_file[13730] <= 8'h00
            reg_file[13731] <= 8'h00
            reg_file[13732] <= 8'h00
            reg_file[13733] <= 8'h00
            reg_file[13734] <= 8'h00
            reg_file[13735] <= 8'h00
            reg_file[13736] <= 8'h00
            reg_file[13737] <= 8'h00
            reg_file[13738] <= 8'h00
            reg_file[13739] <= 8'h00
            reg_file[13740] <= 8'h00
            reg_file[13741] <= 8'h00
            reg_file[13742] <= 8'h00
            reg_file[13743] <= 8'h00
            reg_file[13744] <= 8'h00
            reg_file[13745] <= 8'h00
            reg_file[13746] <= 8'h00
            reg_file[13747] <= 8'h00
            reg_file[13748] <= 8'h00
            reg_file[13749] <= 8'h00
            reg_file[13750] <= 8'h00
            reg_file[13751] <= 8'h00
            reg_file[13752] <= 8'h00
            reg_file[13753] <= 8'h00
            reg_file[13754] <= 8'h00
            reg_file[13755] <= 8'h00
            reg_file[13756] <= 8'h00
            reg_file[13757] <= 8'h00
            reg_file[13758] <= 8'h00
            reg_file[13759] <= 8'h00
            reg_file[13760] <= 8'h00
            reg_file[13761] <= 8'h00
            reg_file[13762] <= 8'h00
            reg_file[13763] <= 8'h00
            reg_file[13764] <= 8'h00
            reg_file[13765] <= 8'h00
            reg_file[13766] <= 8'h00
            reg_file[13767] <= 8'h00
            reg_file[13768] <= 8'h00
            reg_file[13769] <= 8'h00
            reg_file[13770] <= 8'h00
            reg_file[13771] <= 8'h00
            reg_file[13772] <= 8'h00
            reg_file[13773] <= 8'h00
            reg_file[13774] <= 8'h00
            reg_file[13775] <= 8'h00
            reg_file[13776] <= 8'h00
            reg_file[13777] <= 8'h00
            reg_file[13778] <= 8'h00
            reg_file[13779] <= 8'h00
            reg_file[13780] <= 8'h00
            reg_file[13781] <= 8'h00
            reg_file[13782] <= 8'h00
            reg_file[13783] <= 8'h00
            reg_file[13784] <= 8'h00
            reg_file[13785] <= 8'h00
            reg_file[13786] <= 8'h00
            reg_file[13787] <= 8'h00
            reg_file[13788] <= 8'h00
            reg_file[13789] <= 8'h00
            reg_file[13790] <= 8'h00
            reg_file[13791] <= 8'h00
            reg_file[13792] <= 8'h00
            reg_file[13793] <= 8'h00
            reg_file[13794] <= 8'h00
            reg_file[13795] <= 8'h00
            reg_file[13796] <= 8'h00
            reg_file[13797] <= 8'h00
            reg_file[13798] <= 8'h00
            reg_file[13799] <= 8'h00
            reg_file[13800] <= 8'h00
            reg_file[13801] <= 8'h00
            reg_file[13802] <= 8'h00
            reg_file[13803] <= 8'h00
            reg_file[13804] <= 8'h00
            reg_file[13805] <= 8'h00
            reg_file[13806] <= 8'h00
            reg_file[13807] <= 8'h00
            reg_file[13808] <= 8'h00
            reg_file[13809] <= 8'h00
            reg_file[13810] <= 8'h00
            reg_file[13811] <= 8'h00
            reg_file[13812] <= 8'h00
            reg_file[13813] <= 8'h00
            reg_file[13814] <= 8'h00
            reg_file[13815] <= 8'h00
            reg_file[13816] <= 8'h00
            reg_file[13817] <= 8'h00
            reg_file[13818] <= 8'h00
            reg_file[13819] <= 8'h00
            reg_file[13820] <= 8'h00
            reg_file[13821] <= 8'h00
            reg_file[13822] <= 8'h00
            reg_file[13823] <= 8'h00
            reg_file[13824] <= 8'h00
            reg_file[13825] <= 8'h00
            reg_file[13826] <= 8'h00
            reg_file[13827] <= 8'h00
            reg_file[13828] <= 8'h00
            reg_file[13829] <= 8'h00
            reg_file[13830] <= 8'h00
            reg_file[13831] <= 8'h00
            reg_file[13832] <= 8'h00
            reg_file[13833] <= 8'h00
            reg_file[13834] <= 8'h00
            reg_file[13835] <= 8'h00
            reg_file[13836] <= 8'h00
            reg_file[13837] <= 8'h00
            reg_file[13838] <= 8'h00
            reg_file[13839] <= 8'h00
            reg_file[13840] <= 8'h00
            reg_file[13841] <= 8'h00
            reg_file[13842] <= 8'h00
            reg_file[13843] <= 8'h00
            reg_file[13844] <= 8'h00
            reg_file[13845] <= 8'h00
            reg_file[13846] <= 8'h00
            reg_file[13847] <= 8'h00
            reg_file[13848] <= 8'h00
            reg_file[13849] <= 8'h00
            reg_file[13850] <= 8'h00
            reg_file[13851] <= 8'h00
            reg_file[13852] <= 8'h00
            reg_file[13853] <= 8'h00
            reg_file[13854] <= 8'h00
            reg_file[13855] <= 8'h00
            reg_file[13856] <= 8'h00
            reg_file[13857] <= 8'h00
            reg_file[13858] <= 8'h00
            reg_file[13859] <= 8'h00
            reg_file[13860] <= 8'h00
            reg_file[13861] <= 8'h00
            reg_file[13862] <= 8'h00
            reg_file[13863] <= 8'h00
            reg_file[13864] <= 8'h00
            reg_file[13865] <= 8'h00
            reg_file[13866] <= 8'h00
            reg_file[13867] <= 8'h00
            reg_file[13868] <= 8'h00
            reg_file[13869] <= 8'h00
            reg_file[13870] <= 8'h00
            reg_file[13871] <= 8'h00
            reg_file[13872] <= 8'h00
            reg_file[13873] <= 8'h00
            reg_file[13874] <= 8'h00
            reg_file[13875] <= 8'h00
            reg_file[13876] <= 8'h00
            reg_file[13877] <= 8'h00
            reg_file[13878] <= 8'h00
            reg_file[13879] <= 8'h00
            reg_file[13880] <= 8'h00
            reg_file[13881] <= 8'h00
            reg_file[13882] <= 8'h00
            reg_file[13883] <= 8'h00
            reg_file[13884] <= 8'h00
            reg_file[13885] <= 8'h00
            reg_file[13886] <= 8'h00
            reg_file[13887] <= 8'h00
            reg_file[13888] <= 8'h00
            reg_file[13889] <= 8'h00
            reg_file[13890] <= 8'h00
            reg_file[13891] <= 8'h00
            reg_file[13892] <= 8'h00
            reg_file[13893] <= 8'h00
            reg_file[13894] <= 8'h00
            reg_file[13895] <= 8'h00
            reg_file[13896] <= 8'h00
            reg_file[13897] <= 8'h00
            reg_file[13898] <= 8'h00
            reg_file[13899] <= 8'h00
            reg_file[13900] <= 8'h00
            reg_file[13901] <= 8'h00
            reg_file[13902] <= 8'h00
            reg_file[13903] <= 8'h00
            reg_file[13904] <= 8'h00
            reg_file[13905] <= 8'h00
            reg_file[13906] <= 8'h00
            reg_file[13907] <= 8'h00
            reg_file[13908] <= 8'h00
            reg_file[13909] <= 8'h00
            reg_file[13910] <= 8'h00
            reg_file[13911] <= 8'h00
            reg_file[13912] <= 8'h00
            reg_file[13913] <= 8'h00
            reg_file[13914] <= 8'h00
            reg_file[13915] <= 8'h00
            reg_file[13916] <= 8'h00
            reg_file[13917] <= 8'h00
            reg_file[13918] <= 8'h00
            reg_file[13919] <= 8'h00
            reg_file[13920] <= 8'h00
            reg_file[13921] <= 8'h00
            reg_file[13922] <= 8'h00
            reg_file[13923] <= 8'h00
            reg_file[13924] <= 8'h00
            reg_file[13925] <= 8'h00
            reg_file[13926] <= 8'h00
            reg_file[13927] <= 8'h00
            reg_file[13928] <= 8'h00
            reg_file[13929] <= 8'h00
            reg_file[13930] <= 8'h00
            reg_file[13931] <= 8'h00
            reg_file[13932] <= 8'h00
            reg_file[13933] <= 8'h00
            reg_file[13934] <= 8'h00
            reg_file[13935] <= 8'h00
            reg_file[13936] <= 8'h00
            reg_file[13937] <= 8'h00
            reg_file[13938] <= 8'h00
            reg_file[13939] <= 8'h00
            reg_file[13940] <= 8'h00
            reg_file[13941] <= 8'h00
            reg_file[13942] <= 8'h00
            reg_file[13943] <= 8'h00
            reg_file[13944] <= 8'h00
            reg_file[13945] <= 8'h00
            reg_file[13946] <= 8'h00
            reg_file[13947] <= 8'h00
            reg_file[13948] <= 8'h00
            reg_file[13949] <= 8'h00
            reg_file[13950] <= 8'h00
            reg_file[13951] <= 8'h00
            reg_file[13952] <= 8'h00
            reg_file[13953] <= 8'h00
            reg_file[13954] <= 8'h00
            reg_file[13955] <= 8'h00
            reg_file[13956] <= 8'h00
            reg_file[13957] <= 8'h00
            reg_file[13958] <= 8'h00
            reg_file[13959] <= 8'h00
            reg_file[13960] <= 8'h00
            reg_file[13961] <= 8'h00
            reg_file[13962] <= 8'h00
            reg_file[13963] <= 8'h00
            reg_file[13964] <= 8'h00
            reg_file[13965] <= 8'h00
            reg_file[13966] <= 8'h00
            reg_file[13967] <= 8'h00
            reg_file[13968] <= 8'h00
            reg_file[13969] <= 8'h00
            reg_file[13970] <= 8'h00
            reg_file[13971] <= 8'h00
            reg_file[13972] <= 8'h00
            reg_file[13973] <= 8'h00
            reg_file[13974] <= 8'h00
            reg_file[13975] <= 8'h00
            reg_file[13976] <= 8'h00
            reg_file[13977] <= 8'h00
            reg_file[13978] <= 8'h00
            reg_file[13979] <= 8'h00
            reg_file[13980] <= 8'h00
            reg_file[13981] <= 8'h00
            reg_file[13982] <= 8'h00
            reg_file[13983] <= 8'h00
            reg_file[13984] <= 8'h00
            reg_file[13985] <= 8'h00
            reg_file[13986] <= 8'h00
            reg_file[13987] <= 8'h00
            reg_file[13988] <= 8'h00
            reg_file[13989] <= 8'h00
            reg_file[13990] <= 8'h00
            reg_file[13991] <= 8'h00
            reg_file[13992] <= 8'h00
            reg_file[13993] <= 8'h00
            reg_file[13994] <= 8'h00
            reg_file[13995] <= 8'h00
            reg_file[13996] <= 8'h00
            reg_file[13997] <= 8'h00
            reg_file[13998] <= 8'h00
            reg_file[13999] <= 8'h00
            reg_file[14000] <= 8'h00
            reg_file[14001] <= 8'h00
            reg_file[14002] <= 8'h00
            reg_file[14003] <= 8'h00
            reg_file[14004] <= 8'h00
            reg_file[14005] <= 8'h00
            reg_file[14006] <= 8'h00
            reg_file[14007] <= 8'h00
            reg_file[14008] <= 8'h00
            reg_file[14009] <= 8'h00
            reg_file[14010] <= 8'h00
            reg_file[14011] <= 8'h00
            reg_file[14012] <= 8'h00
            reg_file[14013] <= 8'h00
            reg_file[14014] <= 8'h00
            reg_file[14015] <= 8'h00
            reg_file[14016] <= 8'h00
            reg_file[14017] <= 8'h00
            reg_file[14018] <= 8'h00
            reg_file[14019] <= 8'h00
            reg_file[14020] <= 8'h00
            reg_file[14021] <= 8'h00
            reg_file[14022] <= 8'h00
            reg_file[14023] <= 8'h00
            reg_file[14024] <= 8'h00
            reg_file[14025] <= 8'h00
            reg_file[14026] <= 8'h00
            reg_file[14027] <= 8'h00
            reg_file[14028] <= 8'h00
            reg_file[14029] <= 8'h00
            reg_file[14030] <= 8'h00
            reg_file[14031] <= 8'h00
            reg_file[14032] <= 8'h00
            reg_file[14033] <= 8'h00
            reg_file[14034] <= 8'h00
            reg_file[14035] <= 8'h00
            reg_file[14036] <= 8'h00
            reg_file[14037] <= 8'h00
            reg_file[14038] <= 8'h00
            reg_file[14039] <= 8'h00
            reg_file[14040] <= 8'h00
            reg_file[14041] <= 8'h00
            reg_file[14042] <= 8'h00
            reg_file[14043] <= 8'h00
            reg_file[14044] <= 8'h00
            reg_file[14045] <= 8'h00
            reg_file[14046] <= 8'h00
            reg_file[14047] <= 8'h00
            reg_file[14048] <= 8'h00
            reg_file[14049] <= 8'h00
            reg_file[14050] <= 8'h00
            reg_file[14051] <= 8'h00
            reg_file[14052] <= 8'h00
            reg_file[14053] <= 8'h00
            reg_file[14054] <= 8'h00
            reg_file[14055] <= 8'h00
            reg_file[14056] <= 8'h00
            reg_file[14057] <= 8'h00
            reg_file[14058] <= 8'h00
            reg_file[14059] <= 8'h00
            reg_file[14060] <= 8'h00
            reg_file[14061] <= 8'h00
            reg_file[14062] <= 8'h00
            reg_file[14063] <= 8'h00
            reg_file[14064] <= 8'h00
            reg_file[14065] <= 8'h00
            reg_file[14066] <= 8'h00
            reg_file[14067] <= 8'h00
            reg_file[14068] <= 8'h00
            reg_file[14069] <= 8'h00
            reg_file[14070] <= 8'h00
            reg_file[14071] <= 8'h00
            reg_file[14072] <= 8'h00
            reg_file[14073] <= 8'h00
            reg_file[14074] <= 8'h00
            reg_file[14075] <= 8'h00
            reg_file[14076] <= 8'h00
            reg_file[14077] <= 8'h00
            reg_file[14078] <= 8'h00
            reg_file[14079] <= 8'h00
            reg_file[14080] <= 8'h00
            reg_file[14081] <= 8'h00
            reg_file[14082] <= 8'h00
            reg_file[14083] <= 8'h00
            reg_file[14084] <= 8'h00
            reg_file[14085] <= 8'h00
            reg_file[14086] <= 8'h00
            reg_file[14087] <= 8'h00
            reg_file[14088] <= 8'h00
            reg_file[14089] <= 8'h00
            reg_file[14090] <= 8'h00
            reg_file[14091] <= 8'h00
            reg_file[14092] <= 8'h00
            reg_file[14093] <= 8'h00
            reg_file[14094] <= 8'h00
            reg_file[14095] <= 8'h00
            reg_file[14096] <= 8'h00
            reg_file[14097] <= 8'h00
            reg_file[14098] <= 8'h00
            reg_file[14099] <= 8'h00
            reg_file[14100] <= 8'h00
            reg_file[14101] <= 8'h00
            reg_file[14102] <= 8'h00
            reg_file[14103] <= 8'h00
            reg_file[14104] <= 8'h00
            reg_file[14105] <= 8'h00
            reg_file[14106] <= 8'h00
            reg_file[14107] <= 8'h00
            reg_file[14108] <= 8'h00
            reg_file[14109] <= 8'h00
            reg_file[14110] <= 8'h00
            reg_file[14111] <= 8'h00
            reg_file[14112] <= 8'h00
            reg_file[14113] <= 8'h00
            reg_file[14114] <= 8'h00
            reg_file[14115] <= 8'h00
            reg_file[14116] <= 8'h00
            reg_file[14117] <= 8'h00
            reg_file[14118] <= 8'h00
            reg_file[14119] <= 8'h00
            reg_file[14120] <= 8'h00
            reg_file[14121] <= 8'h00
            reg_file[14122] <= 8'h00
            reg_file[14123] <= 8'h00
            reg_file[14124] <= 8'h00
            reg_file[14125] <= 8'h00
            reg_file[14126] <= 8'h00
            reg_file[14127] <= 8'h00
            reg_file[14128] <= 8'h00
            reg_file[14129] <= 8'h00
            reg_file[14130] <= 8'h00
            reg_file[14131] <= 8'h00
            reg_file[14132] <= 8'h00
            reg_file[14133] <= 8'h00
            reg_file[14134] <= 8'h00
            reg_file[14135] <= 8'h00
            reg_file[14136] <= 8'h00
            reg_file[14137] <= 8'h00
            reg_file[14138] <= 8'h00
            reg_file[14139] <= 8'h00
            reg_file[14140] <= 8'h00
            reg_file[14141] <= 8'h00
            reg_file[14142] <= 8'h00
            reg_file[14143] <= 8'h00
            reg_file[14144] <= 8'h00
            reg_file[14145] <= 8'h00
            reg_file[14146] <= 8'h00
            reg_file[14147] <= 8'h00
            reg_file[14148] <= 8'h00
            reg_file[14149] <= 8'h00
            reg_file[14150] <= 8'h00
            reg_file[14151] <= 8'h00
            reg_file[14152] <= 8'h00
            reg_file[14153] <= 8'h00
            reg_file[14154] <= 8'h00
            reg_file[14155] <= 8'h00
            reg_file[14156] <= 8'h00
            reg_file[14157] <= 8'h00
            reg_file[14158] <= 8'h00
            reg_file[14159] <= 8'h00
            reg_file[14160] <= 8'h00
            reg_file[14161] <= 8'h00
            reg_file[14162] <= 8'h00
            reg_file[14163] <= 8'h00
            reg_file[14164] <= 8'h00
            reg_file[14165] <= 8'h00
            reg_file[14166] <= 8'h00
            reg_file[14167] <= 8'h00
            reg_file[14168] <= 8'h00
            reg_file[14169] <= 8'h00
            reg_file[14170] <= 8'h00
            reg_file[14171] <= 8'h00
            reg_file[14172] <= 8'h00
            reg_file[14173] <= 8'h00
            reg_file[14174] <= 8'h00
            reg_file[14175] <= 8'h00
            reg_file[14176] <= 8'h00
            reg_file[14177] <= 8'h00
            reg_file[14178] <= 8'h00
            reg_file[14179] <= 8'h00
            reg_file[14180] <= 8'h00
            reg_file[14181] <= 8'h00
            reg_file[14182] <= 8'h00
            reg_file[14183] <= 8'h00
            reg_file[14184] <= 8'h00
            reg_file[14185] <= 8'h00
            reg_file[14186] <= 8'h00
            reg_file[14187] <= 8'h00
            reg_file[14188] <= 8'h00
            reg_file[14189] <= 8'h00
            reg_file[14190] <= 8'h00
            reg_file[14191] <= 8'h00
            reg_file[14192] <= 8'h00
            reg_file[14193] <= 8'h00
            reg_file[14194] <= 8'h00
            reg_file[14195] <= 8'h00
            reg_file[14196] <= 8'h00
            reg_file[14197] <= 8'h00
            reg_file[14198] <= 8'h00
            reg_file[14199] <= 8'h00
            reg_file[14200] <= 8'h00
            reg_file[14201] <= 8'h00
            reg_file[14202] <= 8'h00
            reg_file[14203] <= 8'h00
            reg_file[14204] <= 8'h00
            reg_file[14205] <= 8'h00
            reg_file[14206] <= 8'h00
            reg_file[14207] <= 8'h00
            reg_file[14208] <= 8'h00
            reg_file[14209] <= 8'h00
            reg_file[14210] <= 8'h00
            reg_file[14211] <= 8'h00
            reg_file[14212] <= 8'h00
            reg_file[14213] <= 8'h00
            reg_file[14214] <= 8'h00
            reg_file[14215] <= 8'h00
            reg_file[14216] <= 8'h00
            reg_file[14217] <= 8'h00
            reg_file[14218] <= 8'h00
            reg_file[14219] <= 8'h00
            reg_file[14220] <= 8'h00
            reg_file[14221] <= 8'h00
            reg_file[14222] <= 8'h00
            reg_file[14223] <= 8'h00
            reg_file[14224] <= 8'h00
            reg_file[14225] <= 8'h00
            reg_file[14226] <= 8'h00
            reg_file[14227] <= 8'h00
            reg_file[14228] <= 8'h00
            reg_file[14229] <= 8'h00
            reg_file[14230] <= 8'h00
            reg_file[14231] <= 8'h00
            reg_file[14232] <= 8'h00
            reg_file[14233] <= 8'h00
            reg_file[14234] <= 8'h00
            reg_file[14235] <= 8'h00
            reg_file[14236] <= 8'h00
            reg_file[14237] <= 8'h00
            reg_file[14238] <= 8'h00
            reg_file[14239] <= 8'h00
            reg_file[14240] <= 8'h00
            reg_file[14241] <= 8'h00
            reg_file[14242] <= 8'h00
            reg_file[14243] <= 8'h00
            reg_file[14244] <= 8'h00
            reg_file[14245] <= 8'h00
            reg_file[14246] <= 8'h00
            reg_file[14247] <= 8'h00
            reg_file[14248] <= 8'h00
            reg_file[14249] <= 8'h00
            reg_file[14250] <= 8'h00
            reg_file[14251] <= 8'h00
            reg_file[14252] <= 8'h00
            reg_file[14253] <= 8'h00
            reg_file[14254] <= 8'h00
            reg_file[14255] <= 8'h00
            reg_file[14256] <= 8'h00
            reg_file[14257] <= 8'h00
            reg_file[14258] <= 8'h00
            reg_file[14259] <= 8'h00
            reg_file[14260] <= 8'h00
            reg_file[14261] <= 8'h00
            reg_file[14262] <= 8'h00
            reg_file[14263] <= 8'h00
            reg_file[14264] <= 8'h00
            reg_file[14265] <= 8'h00
            reg_file[14266] <= 8'h00
            reg_file[14267] <= 8'h00
            reg_file[14268] <= 8'h00
            reg_file[14269] <= 8'h00
            reg_file[14270] <= 8'h00
            reg_file[14271] <= 8'h00
            reg_file[14272] <= 8'h00
            reg_file[14273] <= 8'h00
            reg_file[14274] <= 8'h00
            reg_file[14275] <= 8'h00
            reg_file[14276] <= 8'h00
            reg_file[14277] <= 8'h00
            reg_file[14278] <= 8'h00
            reg_file[14279] <= 8'h00
            reg_file[14280] <= 8'h00
            reg_file[14281] <= 8'h00
            reg_file[14282] <= 8'h00
            reg_file[14283] <= 8'h00
            reg_file[14284] <= 8'h00
            reg_file[14285] <= 8'h00
            reg_file[14286] <= 8'h00
            reg_file[14287] <= 8'h00
            reg_file[14288] <= 8'h00
            reg_file[14289] <= 8'h00
            reg_file[14290] <= 8'h00
            reg_file[14291] <= 8'h00
            reg_file[14292] <= 8'h00
            reg_file[14293] <= 8'h00
            reg_file[14294] <= 8'h00
            reg_file[14295] <= 8'h00
            reg_file[14296] <= 8'h00
            reg_file[14297] <= 8'h00
            reg_file[14298] <= 8'h00
            reg_file[14299] <= 8'h00
            reg_file[14300] <= 8'h00
            reg_file[14301] <= 8'h00
            reg_file[14302] <= 8'h00
            reg_file[14303] <= 8'h00
            reg_file[14304] <= 8'h00
            reg_file[14305] <= 8'h00
            reg_file[14306] <= 8'h00
            reg_file[14307] <= 8'h00
            reg_file[14308] <= 8'h00
            reg_file[14309] <= 8'h00
            reg_file[14310] <= 8'h00
            reg_file[14311] <= 8'h00
            reg_file[14312] <= 8'h00
            reg_file[14313] <= 8'h00
            reg_file[14314] <= 8'h00
            reg_file[14315] <= 8'h00
            reg_file[14316] <= 8'h00
            reg_file[14317] <= 8'h00
            reg_file[14318] <= 8'h00
            reg_file[14319] <= 8'h00
            reg_file[14320] <= 8'h00
            reg_file[14321] <= 8'h00
            reg_file[14322] <= 8'h00
            reg_file[14323] <= 8'h00
            reg_file[14324] <= 8'h00
            reg_file[14325] <= 8'h00
            reg_file[14326] <= 8'h00
            reg_file[14327] <= 8'h00
            reg_file[14328] <= 8'h00
            reg_file[14329] <= 8'h00
            reg_file[14330] <= 8'h00
            reg_file[14331] <= 8'h00
            reg_file[14332] <= 8'h00
            reg_file[14333] <= 8'h00
            reg_file[14334] <= 8'h00
            reg_file[14335] <= 8'h00
            reg_file[14336] <= 8'h00
            reg_file[14337] <= 8'h00
            reg_file[14338] <= 8'h00
            reg_file[14339] <= 8'h00
            reg_file[14340] <= 8'h00
            reg_file[14341] <= 8'h00
            reg_file[14342] <= 8'h00
            reg_file[14343] <= 8'h00
            reg_file[14344] <= 8'h00
            reg_file[14345] <= 8'h00
            reg_file[14346] <= 8'h00
            reg_file[14347] <= 8'h00
            reg_file[14348] <= 8'h00
            reg_file[14349] <= 8'h00
            reg_file[14350] <= 8'h00
            reg_file[14351] <= 8'h00
            reg_file[14352] <= 8'h00
            reg_file[14353] <= 8'h00
            reg_file[14354] <= 8'h00
            reg_file[14355] <= 8'h00
            reg_file[14356] <= 8'h00
            reg_file[14357] <= 8'h00
            reg_file[14358] <= 8'h00
            reg_file[14359] <= 8'h00
            reg_file[14360] <= 8'h00
            reg_file[14361] <= 8'h00
            reg_file[14362] <= 8'h00
            reg_file[14363] <= 8'h00
            reg_file[14364] <= 8'h00
            reg_file[14365] <= 8'h00
            reg_file[14366] <= 8'h00
            reg_file[14367] <= 8'h00
            reg_file[14368] <= 8'h00
            reg_file[14369] <= 8'h00
            reg_file[14370] <= 8'h00
            reg_file[14371] <= 8'h00
            reg_file[14372] <= 8'h00
            reg_file[14373] <= 8'h00
            reg_file[14374] <= 8'h00
            reg_file[14375] <= 8'h00
            reg_file[14376] <= 8'h00
            reg_file[14377] <= 8'h00
            reg_file[14378] <= 8'h00
            reg_file[14379] <= 8'h00
            reg_file[14380] <= 8'h00
            reg_file[14381] <= 8'h00
            reg_file[14382] <= 8'h00
            reg_file[14383] <= 8'h00
            reg_file[14384] <= 8'h00
            reg_file[14385] <= 8'h00
            reg_file[14386] <= 8'h00
            reg_file[14387] <= 8'h00
            reg_file[14388] <= 8'h00
            reg_file[14389] <= 8'h00
            reg_file[14390] <= 8'h00
            reg_file[14391] <= 8'h00
            reg_file[14392] <= 8'h00
            reg_file[14393] <= 8'h00
            reg_file[14394] <= 8'h00
            reg_file[14395] <= 8'h00
            reg_file[14396] <= 8'h00
            reg_file[14397] <= 8'h00
            reg_file[14398] <= 8'h00
            reg_file[14399] <= 8'h00
            reg_file[14400] <= 8'h00
            reg_file[14401] <= 8'h00
            reg_file[14402] <= 8'h00
            reg_file[14403] <= 8'h00
            reg_file[14404] <= 8'h00
            reg_file[14405] <= 8'h00
            reg_file[14406] <= 8'h00
            reg_file[14407] <= 8'h00
            reg_file[14408] <= 8'h00
            reg_file[14409] <= 8'h00
            reg_file[14410] <= 8'h00
            reg_file[14411] <= 8'h00
            reg_file[14412] <= 8'h00
            reg_file[14413] <= 8'h00
            reg_file[14414] <= 8'h00
            reg_file[14415] <= 8'h00
            reg_file[14416] <= 8'h00
            reg_file[14417] <= 8'h00
            reg_file[14418] <= 8'h00
            reg_file[14419] <= 8'h00
            reg_file[14420] <= 8'h00
            reg_file[14421] <= 8'h00
            reg_file[14422] <= 8'h00
            reg_file[14423] <= 8'h00
            reg_file[14424] <= 8'h00
            reg_file[14425] <= 8'h00
            reg_file[14426] <= 8'h00
            reg_file[14427] <= 8'h00
            reg_file[14428] <= 8'h00
            reg_file[14429] <= 8'h00
            reg_file[14430] <= 8'h00
            reg_file[14431] <= 8'h00
            reg_file[14432] <= 8'h00
            reg_file[14433] <= 8'h00
            reg_file[14434] <= 8'h00
            reg_file[14435] <= 8'h00
            reg_file[14436] <= 8'h00
            reg_file[14437] <= 8'h00
            reg_file[14438] <= 8'h00
            reg_file[14439] <= 8'h00
            reg_file[14440] <= 8'h00
            reg_file[14441] <= 8'h00
            reg_file[14442] <= 8'h00
            reg_file[14443] <= 8'h00
            reg_file[14444] <= 8'h00
            reg_file[14445] <= 8'h00
            reg_file[14446] <= 8'h00
            reg_file[14447] <= 8'h00
            reg_file[14448] <= 8'h00
            reg_file[14449] <= 8'h00
            reg_file[14450] <= 8'h00
            reg_file[14451] <= 8'h00
            reg_file[14452] <= 8'h00
            reg_file[14453] <= 8'h00
            reg_file[14454] <= 8'h00
            reg_file[14455] <= 8'h00
            reg_file[14456] <= 8'h00
            reg_file[14457] <= 8'h00
            reg_file[14458] <= 8'h00
            reg_file[14459] <= 8'h00
            reg_file[14460] <= 8'h00
            reg_file[14461] <= 8'h00
            reg_file[14462] <= 8'h00
            reg_file[14463] <= 8'h00
            reg_file[14464] <= 8'h00
            reg_file[14465] <= 8'h00
            reg_file[14466] <= 8'h00
            reg_file[14467] <= 8'h00
            reg_file[14468] <= 8'h00
            reg_file[14469] <= 8'h00
            reg_file[14470] <= 8'h00
            reg_file[14471] <= 8'h00
            reg_file[14472] <= 8'h00
            reg_file[14473] <= 8'h00
            reg_file[14474] <= 8'h00
            reg_file[14475] <= 8'h00
            reg_file[14476] <= 8'h00
            reg_file[14477] <= 8'h00
            reg_file[14478] <= 8'h00
            reg_file[14479] <= 8'h00
            reg_file[14480] <= 8'h00
            reg_file[14481] <= 8'h00
            reg_file[14482] <= 8'h00
            reg_file[14483] <= 8'h00
            reg_file[14484] <= 8'h00
            reg_file[14485] <= 8'h00
            reg_file[14486] <= 8'h00
            reg_file[14487] <= 8'h00
            reg_file[14488] <= 8'h00
            reg_file[14489] <= 8'h00
            reg_file[14490] <= 8'h00
            reg_file[14491] <= 8'h00
            reg_file[14492] <= 8'h00
            reg_file[14493] <= 8'h00
            reg_file[14494] <= 8'h00
            reg_file[14495] <= 8'h00
            reg_file[14496] <= 8'h00
            reg_file[14497] <= 8'h00
            reg_file[14498] <= 8'h00
            reg_file[14499] <= 8'h00
            reg_file[14500] <= 8'h00
            reg_file[14501] <= 8'h00
            reg_file[14502] <= 8'h00
            reg_file[14503] <= 8'h00
            reg_file[14504] <= 8'h00
            reg_file[14505] <= 8'h00
            reg_file[14506] <= 8'h00
            reg_file[14507] <= 8'h00
            reg_file[14508] <= 8'h00
            reg_file[14509] <= 8'h00
            reg_file[14510] <= 8'h00
            reg_file[14511] <= 8'h00
            reg_file[14512] <= 8'h00
            reg_file[14513] <= 8'h00
            reg_file[14514] <= 8'h00
            reg_file[14515] <= 8'h00
            reg_file[14516] <= 8'h00
            reg_file[14517] <= 8'h00
            reg_file[14518] <= 8'h00
            reg_file[14519] <= 8'h00
            reg_file[14520] <= 8'h00
            reg_file[14521] <= 8'h00
            reg_file[14522] <= 8'h00
            reg_file[14523] <= 8'h00
            reg_file[14524] <= 8'h00
            reg_file[14525] <= 8'h00
            reg_file[14526] <= 8'h00
            reg_file[14527] <= 8'h00
            reg_file[14528] <= 8'h00
            reg_file[14529] <= 8'h00
            reg_file[14530] <= 8'h00
            reg_file[14531] <= 8'h00
            reg_file[14532] <= 8'h00
            reg_file[14533] <= 8'h00
            reg_file[14534] <= 8'h00
            reg_file[14535] <= 8'h00
            reg_file[14536] <= 8'h00
            reg_file[14537] <= 8'h00
            reg_file[14538] <= 8'h00
            reg_file[14539] <= 8'h00
            reg_file[14540] <= 8'h00
            reg_file[14541] <= 8'h00
            reg_file[14542] <= 8'h00
            reg_file[14543] <= 8'h00
            reg_file[14544] <= 8'h00
            reg_file[14545] <= 8'h00
            reg_file[14546] <= 8'h00
            reg_file[14547] <= 8'h00
            reg_file[14548] <= 8'h00
            reg_file[14549] <= 8'h00
            reg_file[14550] <= 8'h00
            reg_file[14551] <= 8'h00
            reg_file[14552] <= 8'h00
            reg_file[14553] <= 8'h00
            reg_file[14554] <= 8'h00
            reg_file[14555] <= 8'h00
            reg_file[14556] <= 8'h00
            reg_file[14557] <= 8'h00
            reg_file[14558] <= 8'h00
            reg_file[14559] <= 8'h00
            reg_file[14560] <= 8'h00
            reg_file[14561] <= 8'h00
            reg_file[14562] <= 8'h00
            reg_file[14563] <= 8'h00
            reg_file[14564] <= 8'h00
            reg_file[14565] <= 8'h00
            reg_file[14566] <= 8'h00
            reg_file[14567] <= 8'h00
            reg_file[14568] <= 8'h00
            reg_file[14569] <= 8'h00
            reg_file[14570] <= 8'h00
            reg_file[14571] <= 8'h00
            reg_file[14572] <= 8'h00
            reg_file[14573] <= 8'h00
            reg_file[14574] <= 8'h00
            reg_file[14575] <= 8'h00
            reg_file[14576] <= 8'h00
            reg_file[14577] <= 8'h00
            reg_file[14578] <= 8'h00
            reg_file[14579] <= 8'h00
            reg_file[14580] <= 8'h00
            reg_file[14581] <= 8'h00
            reg_file[14582] <= 8'h00
            reg_file[14583] <= 8'h00
            reg_file[14584] <= 8'h00
            reg_file[14585] <= 8'h00
            reg_file[14586] <= 8'h00
            reg_file[14587] <= 8'h00
            reg_file[14588] <= 8'h00
            reg_file[14589] <= 8'h00
            reg_file[14590] <= 8'h00
            reg_file[14591] <= 8'h00
            reg_file[14592] <= 8'h00
            reg_file[14593] <= 8'h00
            reg_file[14594] <= 8'h00
            reg_file[14595] <= 8'h00
            reg_file[14596] <= 8'h00
            reg_file[14597] <= 8'h00
            reg_file[14598] <= 8'h00
            reg_file[14599] <= 8'h00
            reg_file[14600] <= 8'h00
            reg_file[14601] <= 8'h00
            reg_file[14602] <= 8'h00
            reg_file[14603] <= 8'h00
            reg_file[14604] <= 8'h00
            reg_file[14605] <= 8'h00
            reg_file[14606] <= 8'h00
            reg_file[14607] <= 8'h00
            reg_file[14608] <= 8'h00
            reg_file[14609] <= 8'h00
            reg_file[14610] <= 8'h00
            reg_file[14611] <= 8'h00
            reg_file[14612] <= 8'h00
            reg_file[14613] <= 8'h00
            reg_file[14614] <= 8'h00
            reg_file[14615] <= 8'h00
            reg_file[14616] <= 8'h00
            reg_file[14617] <= 8'h00
            reg_file[14618] <= 8'h00
            reg_file[14619] <= 8'h00
            reg_file[14620] <= 8'h00
            reg_file[14621] <= 8'h00
            reg_file[14622] <= 8'h00
            reg_file[14623] <= 8'h00
            reg_file[14624] <= 8'h00
            reg_file[14625] <= 8'h00
            reg_file[14626] <= 8'h00
            reg_file[14627] <= 8'h00
            reg_file[14628] <= 8'h00
            reg_file[14629] <= 8'h00
            reg_file[14630] <= 8'h00
            reg_file[14631] <= 8'h00
            reg_file[14632] <= 8'h00
            reg_file[14633] <= 8'h00
            reg_file[14634] <= 8'h00
            reg_file[14635] <= 8'h00
            reg_file[14636] <= 8'h00
            reg_file[14637] <= 8'h00
            reg_file[14638] <= 8'h00
            reg_file[14639] <= 8'h00
            reg_file[14640] <= 8'h00
            reg_file[14641] <= 8'h00
            reg_file[14642] <= 8'h00
            reg_file[14643] <= 8'h00
            reg_file[14644] <= 8'h00
            reg_file[14645] <= 8'h00
            reg_file[14646] <= 8'h00
            reg_file[14647] <= 8'h00
            reg_file[14648] <= 8'h00
            reg_file[14649] <= 8'h00
            reg_file[14650] <= 8'h00
            reg_file[14651] <= 8'h00
            reg_file[14652] <= 8'h00
            reg_file[14653] <= 8'h00
            reg_file[14654] <= 8'h00
            reg_file[14655] <= 8'h00
            reg_file[14656] <= 8'h00
            reg_file[14657] <= 8'h00
            reg_file[14658] <= 8'h00
            reg_file[14659] <= 8'h00
            reg_file[14660] <= 8'h00
            reg_file[14661] <= 8'h00
            reg_file[14662] <= 8'h00
            reg_file[14663] <= 8'h00
            reg_file[14664] <= 8'h00
            reg_file[14665] <= 8'h00
            reg_file[14666] <= 8'h00
            reg_file[14667] <= 8'h00
            reg_file[14668] <= 8'h00
            reg_file[14669] <= 8'h00
            reg_file[14670] <= 8'h00
            reg_file[14671] <= 8'h00
            reg_file[14672] <= 8'h00
            reg_file[14673] <= 8'h00
            reg_file[14674] <= 8'h00
            reg_file[14675] <= 8'h00
            reg_file[14676] <= 8'h00
            reg_file[14677] <= 8'h00
            reg_file[14678] <= 8'h00
            reg_file[14679] <= 8'h00
            reg_file[14680] <= 8'h00
            reg_file[14681] <= 8'h00
            reg_file[14682] <= 8'h00
            reg_file[14683] <= 8'h00
            reg_file[14684] <= 8'h00
            reg_file[14685] <= 8'h00
            reg_file[14686] <= 8'h00
            reg_file[14687] <= 8'h00
            reg_file[14688] <= 8'h00
            reg_file[14689] <= 8'h00
            reg_file[14690] <= 8'h00
            reg_file[14691] <= 8'h00
            reg_file[14692] <= 8'h00
            reg_file[14693] <= 8'h00
            reg_file[14694] <= 8'h00
            reg_file[14695] <= 8'h00
            reg_file[14696] <= 8'h00
            reg_file[14697] <= 8'h00
            reg_file[14698] <= 8'h00
            reg_file[14699] <= 8'h00
            reg_file[14700] <= 8'h00
            reg_file[14701] <= 8'h00
            reg_file[14702] <= 8'h00
            reg_file[14703] <= 8'h00
            reg_file[14704] <= 8'h00
            reg_file[14705] <= 8'h00
            reg_file[14706] <= 8'h00
            reg_file[14707] <= 8'h00
            reg_file[14708] <= 8'h00
            reg_file[14709] <= 8'h00
            reg_file[14710] <= 8'h00
            reg_file[14711] <= 8'h00
            reg_file[14712] <= 8'h00
            reg_file[14713] <= 8'h00
            reg_file[14714] <= 8'h00
            reg_file[14715] <= 8'h00
            reg_file[14716] <= 8'h00
            reg_file[14717] <= 8'h00
            reg_file[14718] <= 8'h00
            reg_file[14719] <= 8'h00
            reg_file[14720] <= 8'h00
            reg_file[14721] <= 8'h00
            reg_file[14722] <= 8'h00
            reg_file[14723] <= 8'h00
            reg_file[14724] <= 8'h00
            reg_file[14725] <= 8'h00
            reg_file[14726] <= 8'h00
            reg_file[14727] <= 8'h00
            reg_file[14728] <= 8'h00
            reg_file[14729] <= 8'h00
            reg_file[14730] <= 8'h00
            reg_file[14731] <= 8'h00
            reg_file[14732] <= 8'h00
            reg_file[14733] <= 8'h00
            reg_file[14734] <= 8'h00
            reg_file[14735] <= 8'h00
            reg_file[14736] <= 8'h00
            reg_file[14737] <= 8'h00
            reg_file[14738] <= 8'h00
            reg_file[14739] <= 8'h00
            reg_file[14740] <= 8'h00
            reg_file[14741] <= 8'h00
            reg_file[14742] <= 8'h00
            reg_file[14743] <= 8'h00
            reg_file[14744] <= 8'h00
            reg_file[14745] <= 8'h00
            reg_file[14746] <= 8'h00
            reg_file[14747] <= 8'h00
            reg_file[14748] <= 8'h00
            reg_file[14749] <= 8'h00
            reg_file[14750] <= 8'h00
            reg_file[14751] <= 8'h00
            reg_file[14752] <= 8'h00
            reg_file[14753] <= 8'h00
            reg_file[14754] <= 8'h00
            reg_file[14755] <= 8'h00
            reg_file[14756] <= 8'h00
            reg_file[14757] <= 8'h00
            reg_file[14758] <= 8'h00
            reg_file[14759] <= 8'h00
            reg_file[14760] <= 8'h00
            reg_file[14761] <= 8'h00
            reg_file[14762] <= 8'h00
            reg_file[14763] <= 8'h00
            reg_file[14764] <= 8'h00
            reg_file[14765] <= 8'h00
            reg_file[14766] <= 8'h00
            reg_file[14767] <= 8'h00
            reg_file[14768] <= 8'h00
            reg_file[14769] <= 8'h00
            reg_file[14770] <= 8'h00
            reg_file[14771] <= 8'h00
            reg_file[14772] <= 8'h00
            reg_file[14773] <= 8'h00
            reg_file[14774] <= 8'h00
            reg_file[14775] <= 8'h00
            reg_file[14776] <= 8'h00
            reg_file[14777] <= 8'h00
            reg_file[14778] <= 8'h00
            reg_file[14779] <= 8'h00
            reg_file[14780] <= 8'h00
            reg_file[14781] <= 8'h00
            reg_file[14782] <= 8'h00
            reg_file[14783] <= 8'h00
            reg_file[14784] <= 8'h00
            reg_file[14785] <= 8'h00
            reg_file[14786] <= 8'h00
            reg_file[14787] <= 8'h00
            reg_file[14788] <= 8'h00
            reg_file[14789] <= 8'h00
            reg_file[14790] <= 8'h00
            reg_file[14791] <= 8'h00
            reg_file[14792] <= 8'h00
            reg_file[14793] <= 8'h00
            reg_file[14794] <= 8'h00
            reg_file[14795] <= 8'h00
            reg_file[14796] <= 8'h00
            reg_file[14797] <= 8'h00
            reg_file[14798] <= 8'h00
            reg_file[14799] <= 8'h00
            reg_file[14800] <= 8'h00
            reg_file[14801] <= 8'h00
            reg_file[14802] <= 8'h00
            reg_file[14803] <= 8'h00
            reg_file[14804] <= 8'h00
            reg_file[14805] <= 8'h00
            reg_file[14806] <= 8'h00
            reg_file[14807] <= 8'h00
            reg_file[14808] <= 8'h00
            reg_file[14809] <= 8'h00
            reg_file[14810] <= 8'h00
            reg_file[14811] <= 8'h00
            reg_file[14812] <= 8'h00
            reg_file[14813] <= 8'h00
            reg_file[14814] <= 8'h00
            reg_file[14815] <= 8'h00
            reg_file[14816] <= 8'h00
            reg_file[14817] <= 8'h00
            reg_file[14818] <= 8'h00
            reg_file[14819] <= 8'h00
            reg_file[14820] <= 8'h00
            reg_file[14821] <= 8'h00
            reg_file[14822] <= 8'h00
            reg_file[14823] <= 8'h00
            reg_file[14824] <= 8'h00
            reg_file[14825] <= 8'h00
            reg_file[14826] <= 8'h00
            reg_file[14827] <= 8'h00
            reg_file[14828] <= 8'h00
            reg_file[14829] <= 8'h00
            reg_file[14830] <= 8'h00
            reg_file[14831] <= 8'h00
            reg_file[14832] <= 8'h00
            reg_file[14833] <= 8'h00
            reg_file[14834] <= 8'h00
            reg_file[14835] <= 8'h00
            reg_file[14836] <= 8'h00
            reg_file[14837] <= 8'h00
            reg_file[14838] <= 8'h00
            reg_file[14839] <= 8'h00
            reg_file[14840] <= 8'h00
            reg_file[14841] <= 8'h00
            reg_file[14842] <= 8'h00
            reg_file[14843] <= 8'h00
            reg_file[14844] <= 8'h00
            reg_file[14845] <= 8'h00
            reg_file[14846] <= 8'h00
            reg_file[14847] <= 8'h00
            reg_file[14848] <= 8'h00
            reg_file[14849] <= 8'h00
            reg_file[14850] <= 8'h00
            reg_file[14851] <= 8'h00
            reg_file[14852] <= 8'h00
            reg_file[14853] <= 8'h00
            reg_file[14854] <= 8'h00
            reg_file[14855] <= 8'h00
            reg_file[14856] <= 8'h00
            reg_file[14857] <= 8'h00
            reg_file[14858] <= 8'h00
            reg_file[14859] <= 8'h00
            reg_file[14860] <= 8'h00
            reg_file[14861] <= 8'h00
            reg_file[14862] <= 8'h00
            reg_file[14863] <= 8'h00
            reg_file[14864] <= 8'h00
            reg_file[14865] <= 8'h00
            reg_file[14866] <= 8'h00
            reg_file[14867] <= 8'h00
            reg_file[14868] <= 8'h00
            reg_file[14869] <= 8'h00
            reg_file[14870] <= 8'h00
            reg_file[14871] <= 8'h00
            reg_file[14872] <= 8'h00
            reg_file[14873] <= 8'h00
            reg_file[14874] <= 8'h00
            reg_file[14875] <= 8'h00
            reg_file[14876] <= 8'h00
            reg_file[14877] <= 8'h00
            reg_file[14878] <= 8'h00
            reg_file[14879] <= 8'h00
            reg_file[14880] <= 8'h00
            reg_file[14881] <= 8'h00
            reg_file[14882] <= 8'h00
            reg_file[14883] <= 8'h00
            reg_file[14884] <= 8'h00
            reg_file[14885] <= 8'h00
            reg_file[14886] <= 8'h00
            reg_file[14887] <= 8'h00
            reg_file[14888] <= 8'h00
            reg_file[14889] <= 8'h00
            reg_file[14890] <= 8'h00
            reg_file[14891] <= 8'h00
            reg_file[14892] <= 8'h00
            reg_file[14893] <= 8'h00
            reg_file[14894] <= 8'h00
            reg_file[14895] <= 8'h00
            reg_file[14896] <= 8'h00
            reg_file[14897] <= 8'h00
            reg_file[14898] <= 8'h00
            reg_file[14899] <= 8'h00
            reg_file[14900] <= 8'h00
            reg_file[14901] <= 8'h00
            reg_file[14902] <= 8'h00
            reg_file[14903] <= 8'h00
            reg_file[14904] <= 8'h00
            reg_file[14905] <= 8'h00
            reg_file[14906] <= 8'h00
            reg_file[14907] <= 8'h00
            reg_file[14908] <= 8'h00
            reg_file[14909] <= 8'h00
            reg_file[14910] <= 8'h00
            reg_file[14911] <= 8'h00
            reg_file[14912] <= 8'h00
            reg_file[14913] <= 8'h00
            reg_file[14914] <= 8'h00
            reg_file[14915] <= 8'h00
            reg_file[14916] <= 8'h00
            reg_file[14917] <= 8'h00
            reg_file[14918] <= 8'h00
            reg_file[14919] <= 8'h00
            reg_file[14920] <= 8'h00
            reg_file[14921] <= 8'h00
            reg_file[14922] <= 8'h00
            reg_file[14923] <= 8'h00
            reg_file[14924] <= 8'h00
            reg_file[14925] <= 8'h00
            reg_file[14926] <= 8'h00
            reg_file[14927] <= 8'h00
            reg_file[14928] <= 8'h00
            reg_file[14929] <= 8'h00
            reg_file[14930] <= 8'h00
            reg_file[14931] <= 8'h00
            reg_file[14932] <= 8'h00
            reg_file[14933] <= 8'h00
            reg_file[14934] <= 8'h00
            reg_file[14935] <= 8'h00
            reg_file[14936] <= 8'h00
            reg_file[14937] <= 8'h00
            reg_file[14938] <= 8'h00
            reg_file[14939] <= 8'h00
            reg_file[14940] <= 8'h00
            reg_file[14941] <= 8'h00
            reg_file[14942] <= 8'h00
            reg_file[14943] <= 8'h00
            reg_file[14944] <= 8'h00
            reg_file[14945] <= 8'h00
            reg_file[14946] <= 8'h00
            reg_file[14947] <= 8'h00
            reg_file[14948] <= 8'h00
            reg_file[14949] <= 8'h00
            reg_file[14950] <= 8'h00
            reg_file[14951] <= 8'h00
            reg_file[14952] <= 8'h00
            reg_file[14953] <= 8'h00
            reg_file[14954] <= 8'h00
            reg_file[14955] <= 8'h00
            reg_file[14956] <= 8'h00
            reg_file[14957] <= 8'h00
            reg_file[14958] <= 8'h00
            reg_file[14959] <= 8'h00
            reg_file[14960] <= 8'h00
            reg_file[14961] <= 8'h00
            reg_file[14962] <= 8'h00
            reg_file[14963] <= 8'h00
            reg_file[14964] <= 8'h00
            reg_file[14965] <= 8'h00
            reg_file[14966] <= 8'h00
            reg_file[14967] <= 8'h00
            reg_file[14968] <= 8'h00
            reg_file[14969] <= 8'h00
            reg_file[14970] <= 8'h00
            reg_file[14971] <= 8'h00
            reg_file[14972] <= 8'h00
            reg_file[14973] <= 8'h00
            reg_file[14974] <= 8'h00
            reg_file[14975] <= 8'h00
            reg_file[14976] <= 8'h00
            reg_file[14977] <= 8'h00
            reg_file[14978] <= 8'h00
            reg_file[14979] <= 8'h00
            reg_file[14980] <= 8'h00
            reg_file[14981] <= 8'h00
            reg_file[14982] <= 8'h00
            reg_file[14983] <= 8'h00
            reg_file[14984] <= 8'h00
            reg_file[14985] <= 8'h00
            reg_file[14986] <= 8'h00
            reg_file[14987] <= 8'h00
            reg_file[14988] <= 8'h00
            reg_file[14989] <= 8'h00
            reg_file[14990] <= 8'h00
            reg_file[14991] <= 8'h00
            reg_file[14992] <= 8'h00
            reg_file[14993] <= 8'h00
            reg_file[14994] <= 8'h00
            reg_file[14995] <= 8'h00
            reg_file[14996] <= 8'h00
            reg_file[14997] <= 8'h00
            reg_file[14998] <= 8'h00
            reg_file[14999] <= 8'h00
            reg_file[15000] <= 8'h00
            reg_file[15001] <= 8'h00
            reg_file[15002] <= 8'h00
            reg_file[15003] <= 8'h00
            reg_file[15004] <= 8'h00
            reg_file[15005] <= 8'h00
            reg_file[15006] <= 8'h00
            reg_file[15007] <= 8'h00
            reg_file[15008] <= 8'h00
            reg_file[15009] <= 8'h00
            reg_file[15010] <= 8'h00
            reg_file[15011] <= 8'h00
            reg_file[15012] <= 8'h00
            reg_file[15013] <= 8'h00
            reg_file[15014] <= 8'h00
            reg_file[15015] <= 8'h00
            reg_file[15016] <= 8'h00
            reg_file[15017] <= 8'h00
            reg_file[15018] <= 8'h00
            reg_file[15019] <= 8'h00
            reg_file[15020] <= 8'h00
            reg_file[15021] <= 8'h00
            reg_file[15022] <= 8'h00
            reg_file[15023] <= 8'h00
            reg_file[15024] <= 8'h00
            reg_file[15025] <= 8'h00
            reg_file[15026] <= 8'h00
            reg_file[15027] <= 8'h00
            reg_file[15028] <= 8'h00
            reg_file[15029] <= 8'h00
            reg_file[15030] <= 8'h00
            reg_file[15031] <= 8'h00
            reg_file[15032] <= 8'h00
            reg_file[15033] <= 8'h00
            reg_file[15034] <= 8'h00
            reg_file[15035] <= 8'h00
            reg_file[15036] <= 8'h00
            reg_file[15037] <= 8'h00
            reg_file[15038] <= 8'h00
            reg_file[15039] <= 8'h00
            reg_file[15040] <= 8'h00
            reg_file[15041] <= 8'h00
            reg_file[15042] <= 8'h00
            reg_file[15043] <= 8'h00
            reg_file[15044] <= 8'h00
            reg_file[15045] <= 8'h00
            reg_file[15046] <= 8'h00
            reg_file[15047] <= 8'h00
            reg_file[15048] <= 8'h00
            reg_file[15049] <= 8'h00
            reg_file[15050] <= 8'h00
            reg_file[15051] <= 8'h00
            reg_file[15052] <= 8'h00
            reg_file[15053] <= 8'h00
            reg_file[15054] <= 8'h00
            reg_file[15055] <= 8'h00
            reg_file[15056] <= 8'h00
            reg_file[15057] <= 8'h00
            reg_file[15058] <= 8'h00
            reg_file[15059] <= 8'h00
            reg_file[15060] <= 8'h00
            reg_file[15061] <= 8'h00
            reg_file[15062] <= 8'h00
            reg_file[15063] <= 8'h00
            reg_file[15064] <= 8'h00
            reg_file[15065] <= 8'h00
            reg_file[15066] <= 8'h00
            reg_file[15067] <= 8'h00
            reg_file[15068] <= 8'h00
            reg_file[15069] <= 8'h00
            reg_file[15070] <= 8'h00
            reg_file[15071] <= 8'h00
            reg_file[15072] <= 8'h00
            reg_file[15073] <= 8'h00
            reg_file[15074] <= 8'h00
            reg_file[15075] <= 8'h00
            reg_file[15076] <= 8'h00
            reg_file[15077] <= 8'h00
            reg_file[15078] <= 8'h00
            reg_file[15079] <= 8'h00
            reg_file[15080] <= 8'h00
            reg_file[15081] <= 8'h00
            reg_file[15082] <= 8'h00
            reg_file[15083] <= 8'h00
            reg_file[15084] <= 8'h00
            reg_file[15085] <= 8'h00
            reg_file[15086] <= 8'h00
            reg_file[15087] <= 8'h00
            reg_file[15088] <= 8'h00
            reg_file[15089] <= 8'h00
            reg_file[15090] <= 8'h00
            reg_file[15091] <= 8'h00
            reg_file[15092] <= 8'h00
            reg_file[15093] <= 8'h00
            reg_file[15094] <= 8'h00
            reg_file[15095] <= 8'h00
            reg_file[15096] <= 8'h00
            reg_file[15097] <= 8'h00
            reg_file[15098] <= 8'h00
            reg_file[15099] <= 8'h00
            reg_file[15100] <= 8'h00
            reg_file[15101] <= 8'h00
            reg_file[15102] <= 8'h00
            reg_file[15103] <= 8'h00
            reg_file[15104] <= 8'h00
            reg_file[15105] <= 8'h00
            reg_file[15106] <= 8'h00
            reg_file[15107] <= 8'h00
            reg_file[15108] <= 8'h00
            reg_file[15109] <= 8'h00
            reg_file[15110] <= 8'h00
            reg_file[15111] <= 8'h00
            reg_file[15112] <= 8'h00
            reg_file[15113] <= 8'h00
            reg_file[15114] <= 8'h00
            reg_file[15115] <= 8'h00
            reg_file[15116] <= 8'h00
            reg_file[15117] <= 8'h00
            reg_file[15118] <= 8'h00
            reg_file[15119] <= 8'h00
            reg_file[15120] <= 8'h00
            reg_file[15121] <= 8'h00
            reg_file[15122] <= 8'h00
            reg_file[15123] <= 8'h00
            reg_file[15124] <= 8'h00
            reg_file[15125] <= 8'h00
            reg_file[15126] <= 8'h00
            reg_file[15127] <= 8'h00
            reg_file[15128] <= 8'h00
            reg_file[15129] <= 8'h00
            reg_file[15130] <= 8'h00
            reg_file[15131] <= 8'h00
            reg_file[15132] <= 8'h00
            reg_file[15133] <= 8'h00
            reg_file[15134] <= 8'h00
            reg_file[15135] <= 8'h00
            reg_file[15136] <= 8'h00
            reg_file[15137] <= 8'h00
            reg_file[15138] <= 8'h00
            reg_file[15139] <= 8'h00
            reg_file[15140] <= 8'h00
            reg_file[15141] <= 8'h00
            reg_file[15142] <= 8'h00
            reg_file[15143] <= 8'h00
            reg_file[15144] <= 8'h00
            reg_file[15145] <= 8'h00
            reg_file[15146] <= 8'h00
            reg_file[15147] <= 8'h00
            reg_file[15148] <= 8'h00
            reg_file[15149] <= 8'h00
            reg_file[15150] <= 8'h00
            reg_file[15151] <= 8'h00
            reg_file[15152] <= 8'h00
            reg_file[15153] <= 8'h00
            reg_file[15154] <= 8'h00
            reg_file[15155] <= 8'h00
            reg_file[15156] <= 8'h00
            reg_file[15157] <= 8'h00
            reg_file[15158] <= 8'h00
            reg_file[15159] <= 8'h00
            reg_file[15160] <= 8'h00
            reg_file[15161] <= 8'h00
            reg_file[15162] <= 8'h00
            reg_file[15163] <= 8'h00
            reg_file[15164] <= 8'h00
            reg_file[15165] <= 8'h00
            reg_file[15166] <= 8'h00
            reg_file[15167] <= 8'h00
            reg_file[15168] <= 8'h00
            reg_file[15169] <= 8'h00
            reg_file[15170] <= 8'h00
            reg_file[15171] <= 8'h00
            reg_file[15172] <= 8'h00
            reg_file[15173] <= 8'h00
            reg_file[15174] <= 8'h00
            reg_file[15175] <= 8'h00
            reg_file[15176] <= 8'h00
            reg_file[15177] <= 8'h00
            reg_file[15178] <= 8'h00
            reg_file[15179] <= 8'h00
            reg_file[15180] <= 8'h00
            reg_file[15181] <= 8'h00
            reg_file[15182] <= 8'h00
            reg_file[15183] <= 8'h00
            reg_file[15184] <= 8'h00
            reg_file[15185] <= 8'h00
            reg_file[15186] <= 8'h00
            reg_file[15187] <= 8'h00
            reg_file[15188] <= 8'h00
            reg_file[15189] <= 8'h00
            reg_file[15190] <= 8'h00
            reg_file[15191] <= 8'h00
            reg_file[15192] <= 8'h00
            reg_file[15193] <= 8'h00
            reg_file[15194] <= 8'h00
            reg_file[15195] <= 8'h00
            reg_file[15196] <= 8'h00
            reg_file[15197] <= 8'h00
            reg_file[15198] <= 8'h00
            reg_file[15199] <= 8'h00
            reg_file[15200] <= 8'h00
            reg_file[15201] <= 8'h00
            reg_file[15202] <= 8'h00
            reg_file[15203] <= 8'h00
            reg_file[15204] <= 8'h00
            reg_file[15205] <= 8'h00
            reg_file[15206] <= 8'h00
            reg_file[15207] <= 8'h00
            reg_file[15208] <= 8'h00
            reg_file[15209] <= 8'h00
            reg_file[15210] <= 8'h00
            reg_file[15211] <= 8'h00
            reg_file[15212] <= 8'h00
            reg_file[15213] <= 8'h00
            reg_file[15214] <= 8'h00
            reg_file[15215] <= 8'h00
            reg_file[15216] <= 8'h00
            reg_file[15217] <= 8'h00
            reg_file[15218] <= 8'h00
            reg_file[15219] <= 8'h00
            reg_file[15220] <= 8'h00
            reg_file[15221] <= 8'h00
            reg_file[15222] <= 8'h00
            reg_file[15223] <= 8'h00
            reg_file[15224] <= 8'h00
            reg_file[15225] <= 8'h00
            reg_file[15226] <= 8'h00
            reg_file[15227] <= 8'h00
            reg_file[15228] <= 8'h00
            reg_file[15229] <= 8'h00
            reg_file[15230] <= 8'h00
            reg_file[15231] <= 8'h00
            reg_file[15232] <= 8'h00
            reg_file[15233] <= 8'h00
            reg_file[15234] <= 8'h00
            reg_file[15235] <= 8'h00
            reg_file[15236] <= 8'h00
            reg_file[15237] <= 8'h00
            reg_file[15238] <= 8'h00
            reg_file[15239] <= 8'h00
            reg_file[15240] <= 8'h00
            reg_file[15241] <= 8'h00
            reg_file[15242] <= 8'h00
            reg_file[15243] <= 8'h00
            reg_file[15244] <= 8'h00
            reg_file[15245] <= 8'h00
            reg_file[15246] <= 8'h00
            reg_file[15247] <= 8'h00
            reg_file[15248] <= 8'h00
            reg_file[15249] <= 8'h00
            reg_file[15250] <= 8'h00
            reg_file[15251] <= 8'h00
            reg_file[15252] <= 8'h00
            reg_file[15253] <= 8'h00
            reg_file[15254] <= 8'h00
            reg_file[15255] <= 8'h00
            reg_file[15256] <= 8'h00
            reg_file[15257] <= 8'h00
            reg_file[15258] <= 8'h00
            reg_file[15259] <= 8'h00
            reg_file[15260] <= 8'h00
            reg_file[15261] <= 8'h00
            reg_file[15262] <= 8'h00
            reg_file[15263] <= 8'h00
            reg_file[15264] <= 8'h00
            reg_file[15265] <= 8'h00
            reg_file[15266] <= 8'h00
            reg_file[15267] <= 8'h00
            reg_file[15268] <= 8'h00
            reg_file[15269] <= 8'h00
            reg_file[15270] <= 8'h00
            reg_file[15271] <= 8'h00
            reg_file[15272] <= 8'h00
            reg_file[15273] <= 8'h00
            reg_file[15274] <= 8'h00
            reg_file[15275] <= 8'h00
            reg_file[15276] <= 8'h00
            reg_file[15277] <= 8'h00
            reg_file[15278] <= 8'h00
            reg_file[15279] <= 8'h00
            reg_file[15280] <= 8'h00
            reg_file[15281] <= 8'h00
            reg_file[15282] <= 8'h00
            reg_file[15283] <= 8'h00
            reg_file[15284] <= 8'h00
            reg_file[15285] <= 8'h00
            reg_file[15286] <= 8'h00
            reg_file[15287] <= 8'h00
            reg_file[15288] <= 8'h00
            reg_file[15289] <= 8'h00
            reg_file[15290] <= 8'h00
            reg_file[15291] <= 8'h00
            reg_file[15292] <= 8'h00
            reg_file[15293] <= 8'h00
            reg_file[15294] <= 8'h00
            reg_file[15295] <= 8'h00
            reg_file[15296] <= 8'h00
            reg_file[15297] <= 8'h00
            reg_file[15298] <= 8'h00
            reg_file[15299] <= 8'h00
            reg_file[15300] <= 8'h00
            reg_file[15301] <= 8'h00
            reg_file[15302] <= 8'h00
            reg_file[15303] <= 8'h00
            reg_file[15304] <= 8'h00
            reg_file[15305] <= 8'h00
            reg_file[15306] <= 8'h00
            reg_file[15307] <= 8'h00
            reg_file[15308] <= 8'h00
            reg_file[15309] <= 8'h00
            reg_file[15310] <= 8'h00
            reg_file[15311] <= 8'h00
            reg_file[15312] <= 8'h00
            reg_file[15313] <= 8'h00
            reg_file[15314] <= 8'h00
            reg_file[15315] <= 8'h00
            reg_file[15316] <= 8'h00
            reg_file[15317] <= 8'h00
            reg_file[15318] <= 8'h00
            reg_file[15319] <= 8'h00
            reg_file[15320] <= 8'h00
            reg_file[15321] <= 8'h00
            reg_file[15322] <= 8'h00
            reg_file[15323] <= 8'h00
            reg_file[15324] <= 8'h00
            reg_file[15325] <= 8'h00
            reg_file[15326] <= 8'h00
            reg_file[15327] <= 8'h00
            reg_file[15328] <= 8'h00
            reg_file[15329] <= 8'h00
            reg_file[15330] <= 8'h00
            reg_file[15331] <= 8'h00
            reg_file[15332] <= 8'h00
            reg_file[15333] <= 8'h00
            reg_file[15334] <= 8'h00
            reg_file[15335] <= 8'h00
            reg_file[15336] <= 8'h00
            reg_file[15337] <= 8'h00
            reg_file[15338] <= 8'h00
            reg_file[15339] <= 8'h00
            reg_file[15340] <= 8'h00
            reg_file[15341] <= 8'h00
            reg_file[15342] <= 8'h00
            reg_file[15343] <= 8'h00
            reg_file[15344] <= 8'h00
            reg_file[15345] <= 8'h00
            reg_file[15346] <= 8'h00
            reg_file[15347] <= 8'h00
            reg_file[15348] <= 8'h00
            reg_file[15349] <= 8'h00
            reg_file[15350] <= 8'h00
            reg_file[15351] <= 8'h00
            reg_file[15352] <= 8'h00
            reg_file[15353] <= 8'h00
            reg_file[15354] <= 8'h00
            reg_file[15355] <= 8'h00
            reg_file[15356] <= 8'h00
            reg_file[15357] <= 8'h00
            reg_file[15358] <= 8'h00
            reg_file[15359] <= 8'h00
            reg_file[15360] <= 8'h00
            reg_file[15361] <= 8'h00
            reg_file[15362] <= 8'h00
            reg_file[15363] <= 8'h00
            reg_file[15364] <= 8'h00
            reg_file[15365] <= 8'h00
            reg_file[15366] <= 8'h00
            reg_file[15367] <= 8'h00
            reg_file[15368] <= 8'h00
            reg_file[15369] <= 8'h00
            reg_file[15370] <= 8'h00
            reg_file[15371] <= 8'h00
            reg_file[15372] <= 8'h00
            reg_file[15373] <= 8'h00
            reg_file[15374] <= 8'h00
            reg_file[15375] <= 8'h00
            reg_file[15376] <= 8'h00
            reg_file[15377] <= 8'h00
            reg_file[15378] <= 8'h00
            reg_file[15379] <= 8'h00
            reg_file[15380] <= 8'h00
            reg_file[15381] <= 8'h00
            reg_file[15382] <= 8'h00
            reg_file[15383] <= 8'h00
            reg_file[15384] <= 8'h00
            reg_file[15385] <= 8'h00
            reg_file[15386] <= 8'h00
            reg_file[15387] <= 8'h00
            reg_file[15388] <= 8'h00
            reg_file[15389] <= 8'h00
            reg_file[15390] <= 8'h00
            reg_file[15391] <= 8'h00
            reg_file[15392] <= 8'h00
            reg_file[15393] <= 8'h00
            reg_file[15394] <= 8'h00
            reg_file[15395] <= 8'h00
            reg_file[15396] <= 8'h00
            reg_file[15397] <= 8'h00
            reg_file[15398] <= 8'h00
            reg_file[15399] <= 8'h00
            reg_file[15400] <= 8'h00
            reg_file[15401] <= 8'h00
            reg_file[15402] <= 8'h00
            reg_file[15403] <= 8'h00
            reg_file[15404] <= 8'h00
            reg_file[15405] <= 8'h00
            reg_file[15406] <= 8'h00
            reg_file[15407] <= 8'h00
            reg_file[15408] <= 8'h00
            reg_file[15409] <= 8'h00
            reg_file[15410] <= 8'h00
            reg_file[15411] <= 8'h00
            reg_file[15412] <= 8'h00
            reg_file[15413] <= 8'h00
            reg_file[15414] <= 8'h00
            reg_file[15415] <= 8'h00
            reg_file[15416] <= 8'h00
            reg_file[15417] <= 8'h00
            reg_file[15418] <= 8'h00
            reg_file[15419] <= 8'h00
            reg_file[15420] <= 8'h00
            reg_file[15421] <= 8'h00
            reg_file[15422] <= 8'h00
            reg_file[15423] <= 8'h00
            reg_file[15424] <= 8'h00
            reg_file[15425] <= 8'h00
            reg_file[15426] <= 8'h00
            reg_file[15427] <= 8'h00
            reg_file[15428] <= 8'h00
            reg_file[15429] <= 8'h00
            reg_file[15430] <= 8'h00
            reg_file[15431] <= 8'h00
            reg_file[15432] <= 8'h00
            reg_file[15433] <= 8'h00
            reg_file[15434] <= 8'h00
            reg_file[15435] <= 8'h00
            reg_file[15436] <= 8'h00
            reg_file[15437] <= 8'h00
            reg_file[15438] <= 8'h00
            reg_file[15439] <= 8'h00
            reg_file[15440] <= 8'h00
            reg_file[15441] <= 8'h00
            reg_file[15442] <= 8'h00
            reg_file[15443] <= 8'h00
            reg_file[15444] <= 8'h00
            reg_file[15445] <= 8'h00
            reg_file[15446] <= 8'h00
            reg_file[15447] <= 8'h00
            reg_file[15448] <= 8'h00
            reg_file[15449] <= 8'h00
            reg_file[15450] <= 8'h00
            reg_file[15451] <= 8'h00
            reg_file[15452] <= 8'h00
            reg_file[15453] <= 8'h00
            reg_file[15454] <= 8'h00
            reg_file[15455] <= 8'h00
            reg_file[15456] <= 8'h00
            reg_file[15457] <= 8'h00
            reg_file[15458] <= 8'h00
            reg_file[15459] <= 8'h00
            reg_file[15460] <= 8'h00
            reg_file[15461] <= 8'h00
            reg_file[15462] <= 8'h00
            reg_file[15463] <= 8'h00
            reg_file[15464] <= 8'h00
            reg_file[15465] <= 8'h00
            reg_file[15466] <= 8'h00
            reg_file[15467] <= 8'h00
            reg_file[15468] <= 8'h00
            reg_file[15469] <= 8'h00
            reg_file[15470] <= 8'h00
            reg_file[15471] <= 8'h00
            reg_file[15472] <= 8'h00
            reg_file[15473] <= 8'h00
            reg_file[15474] <= 8'h00
            reg_file[15475] <= 8'h00
            reg_file[15476] <= 8'h00
            reg_file[15477] <= 8'h00
            reg_file[15478] <= 8'h00
            reg_file[15479] <= 8'h00
            reg_file[15480] <= 8'h00
            reg_file[15481] <= 8'h00
            reg_file[15482] <= 8'h00
            reg_file[15483] <= 8'h00
            reg_file[15484] <= 8'h00
            reg_file[15485] <= 8'h00
            reg_file[15486] <= 8'h00
            reg_file[15487] <= 8'h00
            reg_file[15488] <= 8'h00
            reg_file[15489] <= 8'h00
            reg_file[15490] <= 8'h00
            reg_file[15491] <= 8'h00
            reg_file[15492] <= 8'h00
            reg_file[15493] <= 8'h00
            reg_file[15494] <= 8'h00
            reg_file[15495] <= 8'h00
            reg_file[15496] <= 8'h00
            reg_file[15497] <= 8'h00
            reg_file[15498] <= 8'h00
            reg_file[15499] <= 8'h00
            reg_file[15500] <= 8'h00
            reg_file[15501] <= 8'h00
            reg_file[15502] <= 8'h00
            reg_file[15503] <= 8'h00
            reg_file[15504] <= 8'h00
            reg_file[15505] <= 8'h00
            reg_file[15506] <= 8'h00
            reg_file[15507] <= 8'h00
            reg_file[15508] <= 8'h00
            reg_file[15509] <= 8'h00
            reg_file[15510] <= 8'h00
            reg_file[15511] <= 8'h00
            reg_file[15512] <= 8'h00
            reg_file[15513] <= 8'h00
            reg_file[15514] <= 8'h00
            reg_file[15515] <= 8'h00
            reg_file[15516] <= 8'h00
            reg_file[15517] <= 8'h00
            reg_file[15518] <= 8'h00
            reg_file[15519] <= 8'h00
            reg_file[15520] <= 8'h00
            reg_file[15521] <= 8'h00
            reg_file[15522] <= 8'h00
            reg_file[15523] <= 8'h00
            reg_file[15524] <= 8'h00
            reg_file[15525] <= 8'h00
            reg_file[15526] <= 8'h00
            reg_file[15527] <= 8'h00
            reg_file[15528] <= 8'h00
            reg_file[15529] <= 8'h00
            reg_file[15530] <= 8'h00
            reg_file[15531] <= 8'h00
            reg_file[15532] <= 8'h00
            reg_file[15533] <= 8'h00
            reg_file[15534] <= 8'h00
            reg_file[15535] <= 8'h00
            reg_file[15536] <= 8'h00
            reg_file[15537] <= 8'h00
            reg_file[15538] <= 8'h00
            reg_file[15539] <= 8'h00
            reg_file[15540] <= 8'h00
            reg_file[15541] <= 8'h00
            reg_file[15542] <= 8'h00
            reg_file[15543] <= 8'h00
            reg_file[15544] <= 8'h00
            reg_file[15545] <= 8'h00
            reg_file[15546] <= 8'h00
            reg_file[15547] <= 8'h00
            reg_file[15548] <= 8'h00
            reg_file[15549] <= 8'h00
            reg_file[15550] <= 8'h00
            reg_file[15551] <= 8'h00
            reg_file[15552] <= 8'h00
            reg_file[15553] <= 8'h00
            reg_file[15554] <= 8'h00
            reg_file[15555] <= 8'h00
            reg_file[15556] <= 8'h00
            reg_file[15557] <= 8'h00
            reg_file[15558] <= 8'h00
            reg_file[15559] <= 8'h00
            reg_file[15560] <= 8'h00
            reg_file[15561] <= 8'h00
            reg_file[15562] <= 8'h00
            reg_file[15563] <= 8'h00
            reg_file[15564] <= 8'h00
            reg_file[15565] <= 8'h00
            reg_file[15566] <= 8'h00
            reg_file[15567] <= 8'h00
            reg_file[15568] <= 8'h00
            reg_file[15569] <= 8'h00
            reg_file[15570] <= 8'h00
            reg_file[15571] <= 8'h00
            reg_file[15572] <= 8'h00
            reg_file[15573] <= 8'h00
            reg_file[15574] <= 8'h00
            reg_file[15575] <= 8'h00
            reg_file[15576] <= 8'h00
            reg_file[15577] <= 8'h00
            reg_file[15578] <= 8'h00
            reg_file[15579] <= 8'h00
            reg_file[15580] <= 8'h00
            reg_file[15581] <= 8'h00
            reg_file[15582] <= 8'h00
            reg_file[15583] <= 8'h00
            reg_file[15584] <= 8'h00
            reg_file[15585] <= 8'h00
            reg_file[15586] <= 8'h00
            reg_file[15587] <= 8'h00
            reg_file[15588] <= 8'h00
            reg_file[15589] <= 8'h00
            reg_file[15590] <= 8'h00
            reg_file[15591] <= 8'h00
            reg_file[15592] <= 8'h00
            reg_file[15593] <= 8'h00
            reg_file[15594] <= 8'h00
            reg_file[15595] <= 8'h00
            reg_file[15596] <= 8'h00
            reg_file[15597] <= 8'h00
            reg_file[15598] <= 8'h00
            reg_file[15599] <= 8'h00
            reg_file[15600] <= 8'h00
            reg_file[15601] <= 8'h00
            reg_file[15602] <= 8'h00
            reg_file[15603] <= 8'h00
            reg_file[15604] <= 8'h00
            reg_file[15605] <= 8'h00
            reg_file[15606] <= 8'h00
            reg_file[15607] <= 8'h00
            reg_file[15608] <= 8'h00
            reg_file[15609] <= 8'h00
            reg_file[15610] <= 8'h00
            reg_file[15611] <= 8'h00
            reg_file[15612] <= 8'h00
            reg_file[15613] <= 8'h00
            reg_file[15614] <= 8'h00
            reg_file[15615] <= 8'h00
            reg_file[15616] <= 8'h00
            reg_file[15617] <= 8'h00
            reg_file[15618] <= 8'h00
            reg_file[15619] <= 8'h00
            reg_file[15620] <= 8'h00
            reg_file[15621] <= 8'h00
            reg_file[15622] <= 8'h00
            reg_file[15623] <= 8'h00
            reg_file[15624] <= 8'h00
            reg_file[15625] <= 8'h00
            reg_file[15626] <= 8'h00
            reg_file[15627] <= 8'h00
            reg_file[15628] <= 8'h00
            reg_file[15629] <= 8'h00
            reg_file[15630] <= 8'h00
            reg_file[15631] <= 8'h00
            reg_file[15632] <= 8'h00
            reg_file[15633] <= 8'h00
            reg_file[15634] <= 8'h00
            reg_file[15635] <= 8'h00
            reg_file[15636] <= 8'h00
            reg_file[15637] <= 8'h00
            reg_file[15638] <= 8'h00
            reg_file[15639] <= 8'h00
            reg_file[15640] <= 8'h00
            reg_file[15641] <= 8'h00
            reg_file[15642] <= 8'h00
            reg_file[15643] <= 8'h00
            reg_file[15644] <= 8'h00
            reg_file[15645] <= 8'h00
            reg_file[15646] <= 8'h00
            reg_file[15647] <= 8'h00
            reg_file[15648] <= 8'h00
            reg_file[15649] <= 8'h00
            reg_file[15650] <= 8'h00
            reg_file[15651] <= 8'h00
            reg_file[15652] <= 8'h00
            reg_file[15653] <= 8'h00
            reg_file[15654] <= 8'h00
            reg_file[15655] <= 8'h00
            reg_file[15656] <= 8'h00
            reg_file[15657] <= 8'h00
            reg_file[15658] <= 8'h00
            reg_file[15659] <= 8'h00
            reg_file[15660] <= 8'h00
            reg_file[15661] <= 8'h00
            reg_file[15662] <= 8'h00
            reg_file[15663] <= 8'h00
            reg_file[15664] <= 8'h00
            reg_file[15665] <= 8'h00
            reg_file[15666] <= 8'h00
            reg_file[15667] <= 8'h00
            reg_file[15668] <= 8'h00
            reg_file[15669] <= 8'h00
            reg_file[15670] <= 8'h00
            reg_file[15671] <= 8'h00
            reg_file[15672] <= 8'h00
            reg_file[15673] <= 8'h00
            reg_file[15674] <= 8'h00
            reg_file[15675] <= 8'h00
            reg_file[15676] <= 8'h00
            reg_file[15677] <= 8'h00
            reg_file[15678] <= 8'h00
            reg_file[15679] <= 8'h00
            reg_file[15680] <= 8'h00
            reg_file[15681] <= 8'h00
            reg_file[15682] <= 8'h00
            reg_file[15683] <= 8'h00
            reg_file[15684] <= 8'h00
            reg_file[15685] <= 8'h00
            reg_file[15686] <= 8'h00
            reg_file[15687] <= 8'h00
            reg_file[15688] <= 8'h00
            reg_file[15689] <= 8'h00
            reg_file[15690] <= 8'h00
            reg_file[15691] <= 8'h00
            reg_file[15692] <= 8'h00
            reg_file[15693] <= 8'h00
            reg_file[15694] <= 8'h00
            reg_file[15695] <= 8'h00
            reg_file[15696] <= 8'h00
            reg_file[15697] <= 8'h00
            reg_file[15698] <= 8'h00
            reg_file[15699] <= 8'h00
            reg_file[15700] <= 8'h00
            reg_file[15701] <= 8'h00
            reg_file[15702] <= 8'h00
            reg_file[15703] <= 8'h00
            reg_file[15704] <= 8'h00
            reg_file[15705] <= 8'h00
            reg_file[15706] <= 8'h00
            reg_file[15707] <= 8'h00
            reg_file[15708] <= 8'h00
            reg_file[15709] <= 8'h00
            reg_file[15710] <= 8'h00
            reg_file[15711] <= 8'h00
            reg_file[15712] <= 8'h00
            reg_file[15713] <= 8'h00
            reg_file[15714] <= 8'h00
            reg_file[15715] <= 8'h00
            reg_file[15716] <= 8'h00
            reg_file[15717] <= 8'h00
            reg_file[15718] <= 8'h00
            reg_file[15719] <= 8'h00
            reg_file[15720] <= 8'h00
            reg_file[15721] <= 8'h00
            reg_file[15722] <= 8'h00
            reg_file[15723] <= 8'h00
            reg_file[15724] <= 8'h00
            reg_file[15725] <= 8'h00
            reg_file[15726] <= 8'h00
            reg_file[15727] <= 8'h00
            reg_file[15728] <= 8'h00
            reg_file[15729] <= 8'h00
            reg_file[15730] <= 8'h00
            reg_file[15731] <= 8'h00
            reg_file[15732] <= 8'h00
            reg_file[15733] <= 8'h00
            reg_file[15734] <= 8'h00
            reg_file[15735] <= 8'h00
            reg_file[15736] <= 8'h00
            reg_file[15737] <= 8'h00
            reg_file[15738] <= 8'h00
            reg_file[15739] <= 8'h00
            reg_file[15740] <= 8'h00
            reg_file[15741] <= 8'h00
            reg_file[15742] <= 8'h00
            reg_file[15743] <= 8'h00
            reg_file[15744] <= 8'h00
            reg_file[15745] <= 8'h00
            reg_file[15746] <= 8'h00
            reg_file[15747] <= 8'h00
            reg_file[15748] <= 8'h00
            reg_file[15749] <= 8'h00
            reg_file[15750] <= 8'h00
            reg_file[15751] <= 8'h00
            reg_file[15752] <= 8'h00
            reg_file[15753] <= 8'h00
            reg_file[15754] <= 8'h00
            reg_file[15755] <= 8'h00
            reg_file[15756] <= 8'h00
            reg_file[15757] <= 8'h00
            reg_file[15758] <= 8'h00
            reg_file[15759] <= 8'h00
            reg_file[15760] <= 8'h00
            reg_file[15761] <= 8'h00
            reg_file[15762] <= 8'h00
            reg_file[15763] <= 8'h00
            reg_file[15764] <= 8'h00
            reg_file[15765] <= 8'h00
            reg_file[15766] <= 8'h00
            reg_file[15767] <= 8'h00
            reg_file[15768] <= 8'h00
            reg_file[15769] <= 8'h00
            reg_file[15770] <= 8'h00
            reg_file[15771] <= 8'h00
            reg_file[15772] <= 8'h00
            reg_file[15773] <= 8'h00
            reg_file[15774] <= 8'h00
            reg_file[15775] <= 8'h00
            reg_file[15776] <= 8'h00
            reg_file[15777] <= 8'h00
            reg_file[15778] <= 8'h00
            reg_file[15779] <= 8'h00
            reg_file[15780] <= 8'h00
            reg_file[15781] <= 8'h00
            reg_file[15782] <= 8'h00
            reg_file[15783] <= 8'h00
            reg_file[15784] <= 8'h00
            reg_file[15785] <= 8'h00
            reg_file[15786] <= 8'h00
            reg_file[15787] <= 8'h00
            reg_file[15788] <= 8'h00
            reg_file[15789] <= 8'h00
            reg_file[15790] <= 8'h00
            reg_file[15791] <= 8'h00
            reg_file[15792] <= 8'h00
            reg_file[15793] <= 8'h00
            reg_file[15794] <= 8'h00
            reg_file[15795] <= 8'h00
            reg_file[15796] <= 8'h00
            reg_file[15797] <= 8'h00
            reg_file[15798] <= 8'h00
            reg_file[15799] <= 8'h00
            reg_file[15800] <= 8'h00
            reg_file[15801] <= 8'h00
            reg_file[15802] <= 8'h00
            reg_file[15803] <= 8'h00
            reg_file[15804] <= 8'h00
            reg_file[15805] <= 8'h00
            reg_file[15806] <= 8'h00
            reg_file[15807] <= 8'h00
            reg_file[15808] <= 8'h00
            reg_file[15809] <= 8'h00
            reg_file[15810] <= 8'h00
            reg_file[15811] <= 8'h00
            reg_file[15812] <= 8'h00
            reg_file[15813] <= 8'h00
            reg_file[15814] <= 8'h00
            reg_file[15815] <= 8'h00
            reg_file[15816] <= 8'h00
            reg_file[15817] <= 8'h00
            reg_file[15818] <= 8'h00
            reg_file[15819] <= 8'h00
            reg_file[15820] <= 8'h00
            reg_file[15821] <= 8'h00
            reg_file[15822] <= 8'h00
            reg_file[15823] <= 8'h00
            reg_file[15824] <= 8'h00
            reg_file[15825] <= 8'h00
            reg_file[15826] <= 8'h00
            reg_file[15827] <= 8'h00
            reg_file[15828] <= 8'h00
            reg_file[15829] <= 8'h00
            reg_file[15830] <= 8'h00
            reg_file[15831] <= 8'h00
            reg_file[15832] <= 8'h00
            reg_file[15833] <= 8'h00
            reg_file[15834] <= 8'h00
            reg_file[15835] <= 8'h00
            reg_file[15836] <= 8'h00
            reg_file[15837] <= 8'h00
            reg_file[15838] <= 8'h00
            reg_file[15839] <= 8'h00
            reg_file[15840] <= 8'h00
            reg_file[15841] <= 8'h00
            reg_file[15842] <= 8'h00
            reg_file[15843] <= 8'h00
            reg_file[15844] <= 8'h00
            reg_file[15845] <= 8'h00
            reg_file[15846] <= 8'h00
            reg_file[15847] <= 8'h00
            reg_file[15848] <= 8'h00
            reg_file[15849] <= 8'h00
            reg_file[15850] <= 8'h00
            reg_file[15851] <= 8'h00
            reg_file[15852] <= 8'h00
            reg_file[15853] <= 8'h00
            reg_file[15854] <= 8'h00
            reg_file[15855] <= 8'h00
            reg_file[15856] <= 8'h00
            reg_file[15857] <= 8'h00
            reg_file[15858] <= 8'h00
            reg_file[15859] <= 8'h00
            reg_file[15860] <= 8'h00
            reg_file[15861] <= 8'h00
            reg_file[15862] <= 8'h00
            reg_file[15863] <= 8'h00
            reg_file[15864] <= 8'h00
            reg_file[15865] <= 8'h00
            reg_file[15866] <= 8'h00
            reg_file[15867] <= 8'h00
            reg_file[15868] <= 8'h00
            reg_file[15869] <= 8'h00
            reg_file[15870] <= 8'h00
            reg_file[15871] <= 8'h00
            reg_file[15872] <= 8'h00
            reg_file[15873] <= 8'h00
            reg_file[15874] <= 8'h00
            reg_file[15875] <= 8'h00
            reg_file[15876] <= 8'h00
            reg_file[15877] <= 8'h00
            reg_file[15878] <= 8'h00
            reg_file[15879] <= 8'h00
            reg_file[15880] <= 8'h00
            reg_file[15881] <= 8'h00
            reg_file[15882] <= 8'h00
            reg_file[15883] <= 8'h00
            reg_file[15884] <= 8'h00
            reg_file[15885] <= 8'h00
            reg_file[15886] <= 8'h00
            reg_file[15887] <= 8'h00
            reg_file[15888] <= 8'h00
            reg_file[15889] <= 8'h00
            reg_file[15890] <= 8'h00
            reg_file[15891] <= 8'h00
            reg_file[15892] <= 8'h00
            reg_file[15893] <= 8'h00
            reg_file[15894] <= 8'h00
            reg_file[15895] <= 8'h00
            reg_file[15896] <= 8'h00
            reg_file[15897] <= 8'h00
            reg_file[15898] <= 8'h00
            reg_file[15899] <= 8'h00
            reg_file[15900] <= 8'h00
            reg_file[15901] <= 8'h00
            reg_file[15902] <= 8'h00
            reg_file[15903] <= 8'h00
            reg_file[15904] <= 8'h00
            reg_file[15905] <= 8'h00
            reg_file[15906] <= 8'h00
            reg_file[15907] <= 8'h00
            reg_file[15908] <= 8'h00
            reg_file[15909] <= 8'h00
            reg_file[15910] <= 8'h00
            reg_file[15911] <= 8'h00
            reg_file[15912] <= 8'h00
            reg_file[15913] <= 8'h00
            reg_file[15914] <= 8'h00
            reg_file[15915] <= 8'h00
            reg_file[15916] <= 8'h00
            reg_file[15917] <= 8'h00
            reg_file[15918] <= 8'h00
            reg_file[15919] <= 8'h00
            reg_file[15920] <= 8'h00
            reg_file[15921] <= 8'h00
            reg_file[15922] <= 8'h00
            reg_file[15923] <= 8'h00
            reg_file[15924] <= 8'h00
            reg_file[15925] <= 8'h00
            reg_file[15926] <= 8'h00
            reg_file[15927] <= 8'h00
            reg_file[15928] <= 8'h00
            reg_file[15929] <= 8'h00
            reg_file[15930] <= 8'h00
            reg_file[15931] <= 8'h00
            reg_file[15932] <= 8'h00
            reg_file[15933] <= 8'h00
            reg_file[15934] <= 8'h00
            reg_file[15935] <= 8'h00
            reg_file[15936] <= 8'h00
            reg_file[15937] <= 8'h00
            reg_file[15938] <= 8'h00
            reg_file[15939] <= 8'h00
            reg_file[15940] <= 8'h00
            reg_file[15941] <= 8'h00
            reg_file[15942] <= 8'h00
            reg_file[15943] <= 8'h00
            reg_file[15944] <= 8'h00
            reg_file[15945] <= 8'h00
            reg_file[15946] <= 8'h00
            reg_file[15947] <= 8'h00
            reg_file[15948] <= 8'h00
            reg_file[15949] <= 8'h00
            reg_file[15950] <= 8'h00
            reg_file[15951] <= 8'h00
            reg_file[15952] <= 8'h00
            reg_file[15953] <= 8'h00
            reg_file[15954] <= 8'h00
            reg_file[15955] <= 8'h00
            reg_file[15956] <= 8'h00
            reg_file[15957] <= 8'h00
            reg_file[15958] <= 8'h00
            reg_file[15959] <= 8'h00
            reg_file[15960] <= 8'h00
            reg_file[15961] <= 8'h00
            reg_file[15962] <= 8'h00
            reg_file[15963] <= 8'h00
            reg_file[15964] <= 8'h00
            reg_file[15965] <= 8'h00
            reg_file[15966] <= 8'h00
            reg_file[15967] <= 8'h00
            reg_file[15968] <= 8'h00
            reg_file[15969] <= 8'h00
            reg_file[15970] <= 8'h00
            reg_file[15971] <= 8'h00
            reg_file[15972] <= 8'h00
            reg_file[15973] <= 8'h00
            reg_file[15974] <= 8'h00
            reg_file[15975] <= 8'h00
            reg_file[15976] <= 8'h00
            reg_file[15977] <= 8'h00
            reg_file[15978] <= 8'h00
            reg_file[15979] <= 8'h00
            reg_file[15980] <= 8'h00
            reg_file[15981] <= 8'h00
            reg_file[15982] <= 8'h00
            reg_file[15983] <= 8'h00
            reg_file[15984] <= 8'h00
            reg_file[15985] <= 8'h00
            reg_file[15986] <= 8'h00
            reg_file[15987] <= 8'h00
            reg_file[15988] <= 8'h00
            reg_file[15989] <= 8'h00
            reg_file[15990] <= 8'h00
            reg_file[15991] <= 8'h00
            reg_file[15992] <= 8'h00
            reg_file[15993] <= 8'h00
            reg_file[15994] <= 8'h00
            reg_file[15995] <= 8'h00
            reg_file[15996] <= 8'h00
            reg_file[15997] <= 8'h00
            reg_file[15998] <= 8'h00
            reg_file[15999] <= 8'h00
            reg_file[16000] <= 8'h00
            reg_file[16001] <= 8'h00
            reg_file[16002] <= 8'h00
            reg_file[16003] <= 8'h00
            reg_file[16004] <= 8'h00
            reg_file[16005] <= 8'h00
            reg_file[16006] <= 8'h00
            reg_file[16007] <= 8'h00
            reg_file[16008] <= 8'h00
            reg_file[16009] <= 8'h00
            reg_file[16010] <= 8'h00
            reg_file[16011] <= 8'h00
            reg_file[16012] <= 8'h00
            reg_file[16013] <= 8'h00
            reg_file[16014] <= 8'h00
            reg_file[16015] <= 8'h00
            reg_file[16016] <= 8'h00
            reg_file[16017] <= 8'h00
            reg_file[16018] <= 8'h00
            reg_file[16019] <= 8'h00
            reg_file[16020] <= 8'h00
            reg_file[16021] <= 8'h00
            reg_file[16022] <= 8'h00
            reg_file[16023] <= 8'h00
            reg_file[16024] <= 8'h00
            reg_file[16025] <= 8'h00
            reg_file[16026] <= 8'h00
            reg_file[16027] <= 8'h00
            reg_file[16028] <= 8'h00
            reg_file[16029] <= 8'h00
            reg_file[16030] <= 8'h00
            reg_file[16031] <= 8'h00
            reg_file[16032] <= 8'h00
            reg_file[16033] <= 8'h00
            reg_file[16034] <= 8'h00
            reg_file[16035] <= 8'h00
            reg_file[16036] <= 8'h00
            reg_file[16037] <= 8'h00
            reg_file[16038] <= 8'h00
            reg_file[16039] <= 8'h00
            reg_file[16040] <= 8'h00
            reg_file[16041] <= 8'h00
            reg_file[16042] <= 8'h00
            reg_file[16043] <= 8'h00
            reg_file[16044] <= 8'h00
            reg_file[16045] <= 8'h00
            reg_file[16046] <= 8'h00
            reg_file[16047] <= 8'h00
            reg_file[16048] <= 8'h00
            reg_file[16049] <= 8'h00
            reg_file[16050] <= 8'h00
            reg_file[16051] <= 8'h00
            reg_file[16052] <= 8'h00
            reg_file[16053] <= 8'h00
            reg_file[16054] <= 8'h00
            reg_file[16055] <= 8'h00
            reg_file[16056] <= 8'h00
            reg_file[16057] <= 8'h00
            reg_file[16058] <= 8'h00
            reg_file[16059] <= 8'h00
            reg_file[16060] <= 8'h00
            reg_file[16061] <= 8'h00
            reg_file[16062] <= 8'h00
            reg_file[16063] <= 8'h00
            reg_file[16064] <= 8'h00
            reg_file[16065] <= 8'h00
            reg_file[16066] <= 8'h00
            reg_file[16067] <= 8'h00
            reg_file[16068] <= 8'h00
            reg_file[16069] <= 8'h00
            reg_file[16070] <= 8'h00
            reg_file[16071] <= 8'h00
            reg_file[16072] <= 8'h00
            reg_file[16073] <= 8'h00
            reg_file[16074] <= 8'h00
            reg_file[16075] <= 8'h00
            reg_file[16076] <= 8'h00
            reg_file[16077] <= 8'h00
            reg_file[16078] <= 8'h00
            reg_file[16079] <= 8'h00
            reg_file[16080] <= 8'h00
            reg_file[16081] <= 8'h00
            reg_file[16082] <= 8'h00
            reg_file[16083] <= 8'h00
            reg_file[16084] <= 8'h00
            reg_file[16085] <= 8'h00
            reg_file[16086] <= 8'h00
            reg_file[16087] <= 8'h00
            reg_file[16088] <= 8'h00
            reg_file[16089] <= 8'h00
            reg_file[16090] <= 8'h00
            reg_file[16091] <= 8'h00
            reg_file[16092] <= 8'h00
            reg_file[16093] <= 8'h00
            reg_file[16094] <= 8'h00
            reg_file[16095] <= 8'h00
            reg_file[16096] <= 8'h00
            reg_file[16097] <= 8'h00
            reg_file[16098] <= 8'h00
            reg_file[16099] <= 8'h00
            reg_file[16100] <= 8'h00
            reg_file[16101] <= 8'h00
            reg_file[16102] <= 8'h00
            reg_file[16103] <= 8'h00
            reg_file[16104] <= 8'h00
            reg_file[16105] <= 8'h00
            reg_file[16106] <= 8'h00
            reg_file[16107] <= 8'h00
            reg_file[16108] <= 8'h00
            reg_file[16109] <= 8'h00
            reg_file[16110] <= 8'h00
            reg_file[16111] <= 8'h00
            reg_file[16112] <= 8'h00
            reg_file[16113] <= 8'h00
            reg_file[16114] <= 8'h00
            reg_file[16115] <= 8'h00
            reg_file[16116] <= 8'h00
            reg_file[16117] <= 8'h00
            reg_file[16118] <= 8'h00
            reg_file[16119] <= 8'h00
            reg_file[16120] <= 8'h00
            reg_file[16121] <= 8'h00
            reg_file[16122] <= 8'h00
            reg_file[16123] <= 8'h00
            reg_file[16124] <= 8'h00
            reg_file[16125] <= 8'h00
            reg_file[16126] <= 8'h00
            reg_file[16127] <= 8'h00
            reg_file[16128] <= 8'h00
            reg_file[16129] <= 8'h00
            reg_file[16130] <= 8'h00
            reg_file[16131] <= 8'h00
            reg_file[16132] <= 8'h00
            reg_file[16133] <= 8'h00
            reg_file[16134] <= 8'h00
            reg_file[16135] <= 8'h00
            reg_file[16136] <= 8'h00
            reg_file[16137] <= 8'h00
            reg_file[16138] <= 8'h00
            reg_file[16139] <= 8'h00
            reg_file[16140] <= 8'h00
            reg_file[16141] <= 8'h00
            reg_file[16142] <= 8'h00
            reg_file[16143] <= 8'h00
            reg_file[16144] <= 8'h00
            reg_file[16145] <= 8'h00
            reg_file[16146] <= 8'h00
            reg_file[16147] <= 8'h00
            reg_file[16148] <= 8'h00
            reg_file[16149] <= 8'h00
            reg_file[16150] <= 8'h00
            reg_file[16151] <= 8'h00
            reg_file[16152] <= 8'h00
            reg_file[16153] <= 8'h00
            reg_file[16154] <= 8'h00
            reg_file[16155] <= 8'h00
            reg_file[16156] <= 8'h00
            reg_file[16157] <= 8'h00
            reg_file[16158] <= 8'h00
            reg_file[16159] <= 8'h00
            reg_file[16160] <= 8'h00
            reg_file[16161] <= 8'h00
            reg_file[16162] <= 8'h00
            reg_file[16163] <= 8'h00
            reg_file[16164] <= 8'h00
            reg_file[16165] <= 8'h00
            reg_file[16166] <= 8'h00
            reg_file[16167] <= 8'h00
            reg_file[16168] <= 8'h00
            reg_file[16169] <= 8'h00
            reg_file[16170] <= 8'h00
            reg_file[16171] <= 8'h00
            reg_file[16172] <= 8'h00
            reg_file[16173] <= 8'h00
            reg_file[16174] <= 8'h00
            reg_file[16175] <= 8'h00
            reg_file[16176] <= 8'h00
            reg_file[16177] <= 8'h00
            reg_file[16178] <= 8'h00
            reg_file[16179] <= 8'h00
            reg_file[16180] <= 8'h00
            reg_file[16181] <= 8'h00
            reg_file[16182] <= 8'h00
            reg_file[16183] <= 8'h00
            reg_file[16184] <= 8'h00
            reg_file[16185] <= 8'h00
            reg_file[16186] <= 8'h00
            reg_file[16187] <= 8'h00
            reg_file[16188] <= 8'h00
            reg_file[16189] <= 8'h00
            reg_file[16190] <= 8'h00
            reg_file[16191] <= 8'h00
            reg_file[16192] <= 8'h00
            reg_file[16193] <= 8'h00
            reg_file[16194] <= 8'h00
            reg_file[16195] <= 8'h00
            reg_file[16196] <= 8'h00
            reg_file[16197] <= 8'h00
            reg_file[16198] <= 8'h00
            reg_file[16199] <= 8'h00
            reg_file[16200] <= 8'h00
            reg_file[16201] <= 8'h00
            reg_file[16202] <= 8'h00
            reg_file[16203] <= 8'h00
            reg_file[16204] <= 8'h00
            reg_file[16205] <= 8'h00
            reg_file[16206] <= 8'h00
            reg_file[16207] <= 8'h00
            reg_file[16208] <= 8'h00
            reg_file[16209] <= 8'h00
            reg_file[16210] <= 8'h00
            reg_file[16211] <= 8'h00
            reg_file[16212] <= 8'h00
            reg_file[16213] <= 8'h00
            reg_file[16214] <= 8'h00
            reg_file[16215] <= 8'h00
            reg_file[16216] <= 8'h00
            reg_file[16217] <= 8'h00
            reg_file[16218] <= 8'h00
            reg_file[16219] <= 8'h00
            reg_file[16220] <= 8'h00
            reg_file[16221] <= 8'h00
            reg_file[16222] <= 8'h00
            reg_file[16223] <= 8'h00
            reg_file[16224] <= 8'h00
            reg_file[16225] <= 8'h00
            reg_file[16226] <= 8'h00
            reg_file[16227] <= 8'h00
            reg_file[16228] <= 8'h00
            reg_file[16229] <= 8'h00
            reg_file[16230] <= 8'h00
            reg_file[16231] <= 8'h00
            reg_file[16232] <= 8'h00
            reg_file[16233] <= 8'h00
            reg_file[16234] <= 8'h00
            reg_file[16235] <= 8'h00
            reg_file[16236] <= 8'h00
            reg_file[16237] <= 8'h00
            reg_file[16238] <= 8'h00
            reg_file[16239] <= 8'h00
            reg_file[16240] <= 8'h00
            reg_file[16241] <= 8'h00
            reg_file[16242] <= 8'h00
            reg_file[16243] <= 8'h00
            reg_file[16244] <= 8'h00
            reg_file[16245] <= 8'h00
            reg_file[16246] <= 8'h00
            reg_file[16247] <= 8'h00
            reg_file[16248] <= 8'h00
            reg_file[16249] <= 8'h00
            reg_file[16250] <= 8'h00
            reg_file[16251] <= 8'h00
            reg_file[16252] <= 8'h00
            reg_file[16253] <= 8'h00
            reg_file[16254] <= 8'h00
            reg_file[16255] <= 8'h00
            reg_file[16256] <= 8'h00
            reg_file[16257] <= 8'h00
            reg_file[16258] <= 8'h00
            reg_file[16259] <= 8'h00
            reg_file[16260] <= 8'h00
            reg_file[16261] <= 8'h00
            reg_file[16262] <= 8'h00
            reg_file[16263] <= 8'h00
            reg_file[16264] <= 8'h00
            reg_file[16265] <= 8'h00
            reg_file[16266] <= 8'h00
            reg_file[16267] <= 8'h00
            reg_file[16268] <= 8'h00
            reg_file[16269] <= 8'h00
            reg_file[16270] <= 8'h00
            reg_file[16271] <= 8'h00
            reg_file[16272] <= 8'h00
            reg_file[16273] <= 8'h00
            reg_file[16274] <= 8'h00
            reg_file[16275] <= 8'h00
            reg_file[16276] <= 8'h00
            reg_file[16277] <= 8'h00
            reg_file[16278] <= 8'h00
            reg_file[16279] <= 8'h00
            reg_file[16280] <= 8'h00
            reg_file[16281] <= 8'h00
            reg_file[16282] <= 8'h00
            reg_file[16283] <= 8'h00
            reg_file[16284] <= 8'h00
            reg_file[16285] <= 8'h00
            reg_file[16286] <= 8'h00
            reg_file[16287] <= 8'h00
            reg_file[16288] <= 8'h00
            reg_file[16289] <= 8'h00
            reg_file[16290] <= 8'h00
            reg_file[16291] <= 8'h00
            reg_file[16292] <= 8'h00
            reg_file[16293] <= 8'h00
            reg_file[16294] <= 8'h00
            reg_file[16295] <= 8'h00
            reg_file[16296] <= 8'h00
            reg_file[16297] <= 8'h00
            reg_file[16298] <= 8'h00
            reg_file[16299] <= 8'h00
            reg_file[16300] <= 8'h00
            reg_file[16301] <= 8'h00
            reg_file[16302] <= 8'h00
            reg_file[16303] <= 8'h00
            reg_file[16304] <= 8'h00
            reg_file[16305] <= 8'h00
            reg_file[16306] <= 8'h00
            reg_file[16307] <= 8'h00
            reg_file[16308] <= 8'h00
            reg_file[16309] <= 8'h00
            reg_file[16310] <= 8'h00
            reg_file[16311] <= 8'h00
            reg_file[16312] <= 8'h00
            reg_file[16313] <= 8'h00
            reg_file[16314] <= 8'h00
            reg_file[16315] <= 8'h00
            reg_file[16316] <= 8'h00
            reg_file[16317] <= 8'h00
            reg_file[16318] <= 8'h00
            reg_file[16319] <= 8'h00
            reg_file[16320] <= 8'h00
            reg_file[16321] <= 8'h00
            reg_file[16322] <= 8'h00
            reg_file[16323] <= 8'h00
            reg_file[16324] <= 8'h00
            reg_file[16325] <= 8'h00
            reg_file[16326] <= 8'h00
            reg_file[16327] <= 8'h00
            reg_file[16328] <= 8'h00
            reg_file[16329] <= 8'h00
            reg_file[16330] <= 8'h00
            reg_file[16331] <= 8'h00
            reg_file[16332] <= 8'h00
            reg_file[16333] <= 8'h00
            reg_file[16334] <= 8'h00
            reg_file[16335] <= 8'h00
            reg_file[16336] <= 8'h00
            reg_file[16337] <= 8'h00
            reg_file[16338] <= 8'h00
            reg_file[16339] <= 8'h00
            reg_file[16340] <= 8'h00
            reg_file[16341] <= 8'h00
            reg_file[16342] <= 8'h00
            reg_file[16343] <= 8'h00
            reg_file[16344] <= 8'h00
            reg_file[16345] <= 8'h00
            reg_file[16346] <= 8'h00
            reg_file[16347] <= 8'h00
            reg_file[16348] <= 8'h00
            reg_file[16349] <= 8'h00
            reg_file[16350] <= 8'h00
            reg_file[16351] <= 8'h00
            reg_file[16352] <= 8'h00
            reg_file[16353] <= 8'h00
            reg_file[16354] <= 8'h00
            reg_file[16355] <= 8'h00
            reg_file[16356] <= 8'h00
            reg_file[16357] <= 8'h00
            reg_file[16358] <= 8'h00
            reg_file[16359] <= 8'h00
            reg_file[16360] <= 8'h00
            reg_file[16361] <= 8'h00
            reg_file[16362] <= 8'h00
            reg_file[16363] <= 8'h00
            reg_file[16364] <= 8'h00
            reg_file[16365] <= 8'h00
            reg_file[16366] <= 8'h00
            reg_file[16367] <= 8'h00
            reg_file[16368] <= 8'h00
            reg_file[16369] <= 8'h00
            reg_file[16370] <= 8'h00
            reg_file[16371] <= 8'h00
            reg_file[16372] <= 8'h00
            reg_file[16373] <= 8'h00
            reg_file[16374] <= 8'h00
            reg_file[16375] <= 8'h00
            reg_file[16376] <= 8'h00
            reg_file[16377] <= 8'h00
            reg_file[16378] <= 8'h00
            reg_file[16379] <= 8'h00
            reg_file[16380] <= 8'h00
            reg_file[16381] <= 8'h00
            reg_file[16382] <= 8'h00
            reg_file[16383] <= 8'h00
        end
        else
        begin
            reg_file <= next_reg_file;
        end
    end

    // other combinational logic for memory interface
    always_comb begin : OTHER_MEM_COMB_LOGIC

        // mem_req_ready = 1'b1;           // always ready for request
        mem_rsp_valid = mem_req_valid;  // read ready immediately
            // update to buffer to later clock cycle
                // along with data read value

        mem_rsp_tag = mem_req_tag;      // match req immediately
    end

    // delayed mem_req_ready signals
    parameter MEM_REQ_READY_DELAY = 0;
    logic [MEM_REQ_READY_DELAY-1:0] mem_req_ready_reg, next_mem_req_ready_reg; 

    // delayed mem_req_ready reg logic
    always_ff @ (posedge clk) begin : MEM_REQ_READY_REG_LOGIC
    
        if (reset)
        begin
            mem_req_ready_reg = '0;
        end
        else
        begin
            mem_req_ready_reg = next_mem_req_ready_reg;
        end
    end

    // delayed mem_req_ready delay next state logic
    always_comb begin : MEM_REQ_READY_DELAY_NEXT_STATE_LOGIC

        next_mem_req_ready_reg = {mem_req_ready_reg[MEM_REQ_READY_DELAY-2:0], 1'b1};    // shift 1 left
        mem_req_ready = mem_req_ready_reg[MEM_REQ_READY_DELAY-1];                       // msb of shifter
    end

    // NOTES:
    // don't know what to do with: 
        // busy

endmodule

