/*
    socet115 / zlagpaca@purdue.edu
    Zach Lagpacan

    module for faking memory with basic register file which can interface with Vortex memory interface
*/

// temporary include to have defined vals
// `include "local_mem.vh"
`include "../include/VX_define.vh"
// `include "VX_define.vh"

module local_mem #(
)(
    // seq
    input clk, reset,

    // Memory Request:
    // vortex outputs
    input logic                             mem_req_valid,
    input logic                             mem_req_rw,
    input logic [`VX_MEM_BYTEEN_WIDTH-1:0]  mem_req_byteen, // 64 (512 / 8)
    input logic [`VX_MEM_ADDR_WIDTH-1:0]    mem_req_addr,   // 26
    input logic [`VX_MEM_DATA_WIDTH-1:0]    mem_req_data,   // 512
    input logic [`VX_MEM_TAG_WIDTH-1:0]     mem_req_tag,    // 56 (55 for SM disabled)
    // vortex inputs
    output logic                            mem_req_ready,

    // Memory response:
    // vortex inputs
    output logic                            mem_rsp_valid,        
    output logic [`VX_MEM_DATA_WIDTH-1:0]   mem_rsp_data,   // 512
    output logic [`VX_MEM_TAG_WIDTH-1:0]    mem_rsp_tag,    // 56 (55 for SM disabled)
    // vortex outputs
    input logic                             mem_rsp_ready,

    // Status:
    // vortex outputs
    input logic                             busy,

    // tb:
    output logic                            tb_addr_out_of_bounds
);
    // register file instances
    
    // chunk 0
    logic wen_0_80000000;
    logic [6-1:0] wsel_0_80000000;
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_0_80000000;
    logic [6-1:0] rsel_0_80000000;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_0_80000000;
    
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_0_80000000 [64-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_0_80000000 [64-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_0_80000000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_0_80000000[0][31:0] <= 32'hFC102573;
            reg_val_0_80000000[0][63:32] <= 32'h00000597;
            reg_val_0_80000000[0][95:64] <= 32'h09C58593;
            reg_val_0_80000000[0][127:96] <= 32'h00B5106B;
            reg_val_0_80000000[0][159:128] <= 32'h090000EF;
            reg_val_0_80000000[0][191:160] <= 32'h00100513;
            reg_val_0_80000000[0][223:192] <= 32'h0005006B;
            reg_val_0_80000000[0][255:224] <= 32'hFC102573;
            reg_val_0_80000000[0][287:256] <= 32'h00000597;
            reg_val_0_80000000[0][319:288] <= 32'h12058593;
            reg_val_0_80000000[0][351:320] <= 32'h00B5106B;
            reg_val_0_80000000[0][383:352] <= 32'h114000EF;
            reg_val_0_80000000[0][415:384] <= 32'h00100513;
            reg_val_0_80000000[0][447:416] <= 32'h0005006B;
            reg_val_0_80000000[0][479:448] <= 32'h00001517;
            reg_val_0_80000000[0][511:480] <= 32'h40850513;
            reg_val_0_80000000[1][31:0] <= 32'h00001617;
            reg_val_0_80000000[1][63:32] <= 32'h48060613;
            reg_val_0_80000000[1][95:64] <= 32'h40A60633;
            reg_val_0_80000000[1][127:96] <= 32'h00000593;
            reg_val_0_80000000[1][159:128] <= 32'h29D000EF;
            reg_val_0_80000000[1][191:160] <= 32'h00000517;
            reg_val_0_80000000[1][223:192] <= 32'h1DC50513;
            reg_val_0_80000000[1][255:224] <= 32'h12D000EF;
            reg_val_0_80000000[1][287:256] <= 32'h13C000EF;
            reg_val_0_80000000[1][319:288] <= 32'h008000EF;
            reg_val_0_80000000[1][351:320] <= 32'h1350006F;
            reg_val_0_80000000[1][383:352] <= 32'hFFF00793;
            reg_val_0_80000000[1][415:384] <= 32'h0007806B;
            reg_val_0_80000000[1][447:416] <= 32'h00000513;
            reg_val_0_80000000[1][479:448] <= 32'h00008067;
            reg_val_0_80000000[1][511:480] <= 32'h00000793;
            reg_val_0_80000000[2][31:0] <= 32'h00078863;
            reg_val_0_80000000[2][63:32] <= 32'h80000537;
            reg_val_0_80000000[2][95:64] <= 32'h23050513;
            reg_val_0_80000000[2][127:96] <= 32'h0FD0006F;
            reg_val_0_80000000[2][159:128] <= 32'h00008067;
            reg_val_0_80000000[2][191:160] <= 32'h00040193;
            reg_val_0_80000000[2][223:192] <= 32'h00000513;
            reg_val_0_80000000[2][255:224] <= 32'h0005006B;
            reg_val_0_80000000[2][287:256] <= 32'hFFF00513;
            reg_val_0_80000000[2][319:288] <= 32'h0005006B;
            reg_val_0_80000000[2][351:320] <= 32'h00001197;
            reg_val_0_80000000[2][383:352] <= 32'h76018193;
            reg_val_0_80000000[2][415:384] <= 32'hFF000137;
            reg_val_0_80000000[2][447:416] <= 32'hCC102573;
            reg_val_0_80000000[2][479:448] <= 32'h00A51593;
            reg_val_0_80000000[2][511:480] <= 32'h40B10133;
            reg_val_0_80000000[3][31:0] <= 32'h00000593;
            reg_val_0_80000000[3][63:32] <= 32'h02B50533;
            reg_val_0_80000000[3][95:64] <= 32'h00001217;
            reg_val_0_80000000[3][127:96] <= 32'h43720213;
            reg_val_0_80000000[3][159:128] <= 32'h00A20233;
            reg_val_0_80000000[3][191:160] <= 32'hFC027213;
            reg_val_0_80000000[3][223:192] <= 32'hCC3026F3;
            reg_val_0_80000000[3][255:224] <= 32'h00068663;
            reg_val_0_80000000[3][287:256] <= 32'h00000513;
            reg_val_0_80000000[3][319:288] <= 32'h0005006B;
            reg_val_0_80000000[3][351:320] <= 32'h00008067;
            reg_val_0_80000000[3][383:352] <= 32'hFFF00513;
            reg_val_0_80000000[3][415:384] <= 32'h00008067;
            reg_val_0_80000000[3][447:416] <= 32'hFFF00513;
            reg_val_0_80000000[3][479:448] <= 32'h00008067;
            reg_val_0_80000000[3][511:480] <= 32'h00000513;
            reg_val_0_80000000[4][31:0] <= 32'h00008067;
            reg_val_0_80000000[4][63:32] <= 32'h00000513;
            reg_val_0_80000000[4][95:64] <= 32'h00008067;
            reg_val_0_80000000[4][127:96] <= 32'hFFF00513;
            reg_val_0_80000000[4][159:128] <= 32'h00008067;
            reg_val_0_80000000[4][191:160] <= 32'hFFF00513;
            reg_val_0_80000000[4][223:192] <= 32'h00008067;
            reg_val_0_80000000[4][255:224] <= 32'h00100073;
            reg_val_0_80000000[4][287:256] <= 32'h00000513;
            reg_val_0_80000000[4][319:288] <= 32'h00008067;
            reg_val_0_80000000[4][351:320] <= 32'h00060513;
            reg_val_0_80000000[4][383:352] <= 32'h00008067;
            reg_val_0_80000000[4][415:384] <= 32'hFFF00513;
            reg_val_0_80000000[4][447:416] <= 32'h00008067;
            reg_val_0_80000000[4][479:448] <= 32'hF1402573;
            reg_val_0_80000000[4][511:480] <= 32'h00008067;
            reg_val_0_80000000[5][31:0] <= 32'hFF010113;
            reg_val_0_80000000[5][63:32] <= 32'h00112623;
            reg_val_0_80000000[5][95:64] <= 32'h00812423;
            reg_val_0_80000000[5][127:96] <= 32'hFFF00793;
            reg_val_0_80000000[5][159:128] <= 32'h0007806B;
            reg_val_0_80000000[5][191:160] <= 32'h00000613;
            reg_val_0_80000000[5][223:192] <= 32'h00020513;
            reg_val_0_80000000[5][255:224] <= 32'h00001597;
            reg_val_0_80000000[5][287:256] <= 32'hEA458593;
            reg_val_0_80000000[5][319:288] <= 32'h00020413;
            reg_val_0_80000000[5][351:320] <= 32'h069000EF;
            reg_val_0_80000000[5][383:352] <= 32'h00000513;
            reg_val_0_80000000[5][415:384] <= 32'h00000613;
            reg_val_0_80000000[5][447:416] <= 32'h00000593;
            reg_val_0_80000000[5][479:448] <= 32'h00A40533;
            reg_val_0_80000000[5][511:480] <= 32'h171000EF;
            reg_val_0_80000000[6][31:0] <= 32'hCC3027F3;
            reg_val_0_80000000[6][63:32] <= 32'h0017B793;
            reg_val_0_80000000[6][95:64] <= 32'h0007806B;
            reg_val_0_80000000[6][127:96] <= 32'h00C12083;
            reg_val_0_80000000[6][159:128] <= 32'h00812403;
            reg_val_0_80000000[6][191:160] <= 32'h01010113;
            reg_val_0_80000000[6][223:192] <= 32'h00008067;
            reg_val_0_80000000[6][255:224] <= 32'hFF010113;
            reg_val_0_80000000[6][287:256] <= 32'h00812423;
            reg_val_0_80000000[6][319:288] <= 32'h01212023;
            reg_val_0_80000000[6][351:320] <= 32'h00001417;
            reg_val_0_80000000[6][383:352] <= 32'hE5840413;
            reg_val_0_80000000[6][415:384] <= 32'h00001917;
            reg_val_0_80000000[6][447:416] <= 32'hE5090913;
            reg_val_0_80000000[6][479:448] <= 32'h40890933;
            reg_val_0_80000000[6][511:480] <= 32'h00112623;
            reg_val_0_80000000[7][31:0] <= 32'h00912223;
            reg_val_0_80000000[7][63:32] <= 32'h40295913;
            reg_val_0_80000000[7][95:64] <= 32'h00090E63;
            reg_val_0_80000000[7][127:96] <= 32'h00000493;
            reg_val_0_80000000[7][159:128] <= 32'h00042783;
            reg_val_0_80000000[7][191:160] <= 32'h00148493;
            reg_val_0_80000000[7][223:192] <= 32'h00440413;
            reg_val_0_80000000[7][255:224] <= 32'h000780E7;
            reg_val_0_80000000[7][287:256] <= 32'hFE9918E3;
            reg_val_0_80000000[7][319:288] <= 32'h00001417;
            reg_val_0_80000000[7][351:320] <= 32'hE1C40413;
            reg_val_0_80000000[7][383:352] <= 32'h00001917;
            reg_val_0_80000000[7][415:384] <= 32'hE1890913;
            reg_val_0_80000000[7][447:416] <= 32'h40890933;
            reg_val_0_80000000[7][479:448] <= 32'h40295913;
            reg_val_0_80000000[7][511:480] <= 32'h00090E63;
            reg_val_0_80000000[8][31:0] <= 32'h00000493;
            reg_val_0_80000000[8][63:32] <= 32'h00042783;
            reg_val_0_80000000[8][95:64] <= 32'h00148493;
            reg_val_0_80000000[8][127:96] <= 32'h00440413;
            reg_val_0_80000000[8][159:128] <= 32'h000780E7;
            reg_val_0_80000000[8][191:160] <= 32'hFE9918E3;
            reg_val_0_80000000[8][223:192] <= 32'h00C12083;
            reg_val_0_80000000[8][255:224] <= 32'h00812403;
            reg_val_0_80000000[8][287:256] <= 32'h00412483;
            reg_val_0_80000000[8][319:288] <= 32'h00012903;
            reg_val_0_80000000[8][351:320] <= 32'h01010113;
            reg_val_0_80000000[8][383:352] <= 32'h00008067;
            reg_val_0_80000000[8][415:384] <= 32'hFF010113;
            reg_val_0_80000000[8][447:416] <= 32'h00812423;
            reg_val_0_80000000[8][479:448] <= 32'h00001797;
            reg_val_0_80000000[8][511:480] <= 32'hDCC78793;
            reg_val_0_80000000[9][31:0] <= 32'h00001417;
            reg_val_0_80000000[9][63:32] <= 32'hDC440413;
            reg_val_0_80000000[9][95:64] <= 32'h408787B3;
            reg_val_0_80000000[9][127:96] <= 32'h00912223;
            reg_val_0_80000000[9][159:128] <= 32'h00112623;
            reg_val_0_80000000[9][191:160] <= 32'h4027D493;
            reg_val_0_80000000[9][223:192] <= 32'h02048063;
            reg_val_0_80000000[9][255:224] <= 32'hFFC78793;
            reg_val_0_80000000[9][287:256] <= 32'h00878433;
            reg_val_0_80000000[9][319:288] <= 32'h00042783;
            reg_val_0_80000000[9][351:320] <= 32'hFFF48493;
            reg_val_0_80000000[9][383:352] <= 32'hFFC40413;
            reg_val_0_80000000[9][415:384] <= 32'h000780E7;
            reg_val_0_80000000[9][447:416] <= 32'hFE0498E3;
            reg_val_0_80000000[9][479:448] <= 32'h00C12083;
            reg_val_0_80000000[9][511:480] <= 32'h00812403;
            reg_val_0_80000000[10][31:0] <= 32'h00412483;
            reg_val_0_80000000[10][63:32] <= 32'h01010113;
            reg_val_0_80000000[10][95:64] <= 32'h00008067;
            reg_val_0_80000000[10][127:96] <= 32'hFF010113;
            reg_val_0_80000000[10][159:128] <= 32'h00112623;
            reg_val_0_80000000[10][191:160] <= 32'h00812423;
            reg_val_0_80000000[10][223:192] <= 32'h00912223;
            reg_val_0_80000000[10][255:224] <= 32'h01212023;
            reg_val_0_80000000[10][287:256] <= 32'hCC5027F3;
            reg_val_0_80000000[10][319:288] <= 32'hCC302773;
            reg_val_0_80000000[10][351:320] <= 32'hCC0026F3;
            reg_val_0_80000000[10][383:352] <= 32'hFC0025F3;
            reg_val_0_80000000[10][415:384] <= 32'h00279613;
            reg_val_0_80000000[10][447:416] <= 32'h00001797;
            reg_val_0_80000000[10][479:448] <= 32'h18C78793;
            reg_val_0_80000000[10][511:480] <= 32'h00C787B3;
            reg_val_0_80000000[11][31:0] <= 32'h0007A483;
            reg_val_0_80000000[11][63:32] <= 32'h0104A403;
            reg_val_0_80000000[11][95:64] <= 32'h00C4A603;
            reg_val_0_80000000[11][127:96] <= 32'h00872933;
            reg_val_0_80000000[11][159:128] <= 32'h00040793;
            reg_val_0_80000000[11][191:160] <= 32'h00C90933;
            reg_val_0_80000000[11][223:192] <= 32'h02E60433;
            reg_val_0_80000000[11][255:224] <= 32'h00F75463;
            reg_val_0_80000000[11][287:256] <= 32'h00070793;
            reg_val_0_80000000[11][319:288] <= 32'h00F40433;
            reg_val_0_80000000[11][351:320] <= 32'h0084A703;
            reg_val_0_80000000[11][383:352] <= 32'h02B40433;
            reg_val_0_80000000[11][415:384] <= 32'h02D907B3;
            reg_val_0_80000000[11][447:416] <= 32'h00E40433;
            reg_val_0_80000000[11][479:448] <= 32'h00F40433;
            reg_val_0_80000000[11][511:480] <= 32'h00890933;
            reg_val_0_80000000[12][31:0] <= 32'h01245E63;
            reg_val_0_80000000[12][63:32] <= 32'h0004A783;
            reg_val_0_80000000[12][95:64] <= 32'h0044A583;
            reg_val_0_80000000[12][127:96] <= 32'h00040513;
            reg_val_0_80000000[12][159:128] <= 32'h00140413;
            reg_val_0_80000000[12][191:160] <= 32'h000780E7;
            reg_val_0_80000000[12][223:192] <= 32'hFE8916E3;
            reg_val_0_80000000[12][255:224] <= 32'h0144A703;
            reg_val_0_80000000[12][287:256] <= 32'h00000793;
            reg_val_0_80000000[12][319:288] <= 32'h00E7C06B;
            reg_val_0_80000000[12][351:320] <= 32'h00C12083;
            reg_val_0_80000000[12][383:352] <= 32'h00812403;
            reg_val_0_80000000[12][415:384] <= 32'h00412483;
            reg_val_0_80000000[12][447:416] <= 32'h00012903;
            reg_val_0_80000000[12][479:448] <= 32'h01010113;
            reg_val_0_80000000[12][511:480] <= 32'h00008067;
            reg_val_0_80000000[13][31:0] <= 32'hCC5027F3;
            reg_val_0_80000000[13][63:32] <= 32'hCC202573;
            reg_val_0_80000000[13][95:64] <= 32'h00279713;
            reg_val_0_80000000[13][127:96] <= 32'h00001797;
            reg_val_0_80000000[13][159:128] <= 32'h0F478793;
            reg_val_0_80000000[13][191:160] <= 32'h00E787B3;
            reg_val_0_80000000[13][223:192] <= 32'h0007A783;
            reg_val_0_80000000[13][255:224] <= 32'h0087A703;
            reg_val_0_80000000[13][287:256] <= 32'h0007A303;
            reg_val_0_80000000[13][319:288] <= 32'h0047A583;
            reg_val_0_80000000[13][351:320] <= 32'h00E50533;
            reg_val_0_80000000[13][383:352] <= 32'h00030067;
            reg_val_0_80000000[13][415:384] <= 32'hFF010113;
            reg_val_0_80000000[13][447:416] <= 32'h00112623;
            reg_val_0_80000000[13][479:448] <= 32'hFFF00793;
            reg_val_0_80000000[13][511:480] <= 32'h0007806B;
            reg_val_0_80000000[14][31:0] <= 32'hF0DFF0EF;
            reg_val_0_80000000[14][63:32] <= 32'hCC3027F3;
            reg_val_0_80000000[14][95:64] <= 32'h0017B793;
            reg_val_0_80000000[14][127:96] <= 32'h0007806B;
            reg_val_0_80000000[14][159:128] <= 32'h00C12083;
            reg_val_0_80000000[14][191:160] <= 32'h01010113;
            reg_val_0_80000000[14][223:192] <= 32'h00008067;
            reg_val_0_80000000[14][255:224] <= 32'hFE010113;
            reg_val_0_80000000[14][287:256] <= 32'h00112E23;
            reg_val_0_80000000[14][319:288] <= 32'h00812C23;
            reg_val_0_80000000[14][351:320] <= 32'h00912A23;
            reg_val_0_80000000[14][383:352] <= 32'h01212823;
            reg_val_0_80000000[14][415:384] <= 32'h01312623;
            reg_val_0_80000000[14][447:416] <= 32'h01412423;
            reg_val_0_80000000[14][479:448] <= 32'hCC5027F3;
            reg_val_0_80000000[14][511:480] <= 32'hCC302773;
            reg_val_0_80000000[15][31:0] <= 32'hCC0026F3;
            reg_val_0_80000000[15][63:32] <= 32'hFC002573;
            reg_val_0_80000000[15][95:64] <= 32'h00279613;
            reg_val_0_80000000[15][127:96] <= 32'h00001797;
            reg_val_0_80000000[15][159:128] <= 32'h07478793;
            reg_val_0_80000000[15][191:160] <= 32'h00C787B3;
            reg_val_0_80000000[15][223:192] <= 32'h0007A403;
            reg_val_0_80000000[15][255:224] <= 32'h01442483;
            reg_val_0_80000000[15][287:256] <= 32'h01042603;
            reg_val_0_80000000[15][319:288] <= 32'h00972A33;
            reg_val_0_80000000[15][351:320] <= 32'h00048793;
            reg_val_0_80000000[15][383:352] <= 32'h00CA0A33;
            reg_val_0_80000000[15][415:384] <= 32'h02E604B3;
            reg_val_0_80000000[15][447:416] <= 32'h00F75463;
            reg_val_0_80000000[15][479:448] <= 32'h00070793;
            reg_val_0_80000000[15][511:480] <= 32'h00F484B3;
            reg_val_0_80000000[16][31:0] <= 32'h00042583;
            reg_val_0_80000000[16][63:32] <= 32'h00C42703;
            reg_val_0_80000000[16][95:64] <= 32'h0005A903;
            reg_val_0_80000000[16][127:96] <= 32'h0045A983;
            reg_val_0_80000000[16][159:128] <= 32'h02A484B3;
            reg_val_0_80000000[16][191:160] <= 32'h02DA07B3;
            reg_val_0_80000000[16][223:192] <= 32'h00E484B3;
            reg_val_0_80000000[16][255:224] <= 32'h00F484B3;
            reg_val_0_80000000[16][287:256] <= 32'h009A0A33;
            reg_val_0_80000000[16][319:288] <= 32'h033909B3;
            reg_val_0_80000000[16][351:320] <= 32'h0744C063;
            reg_val_0_80000000[16][383:352] <= 32'h0800006F;
            reg_val_0_80000000[16][415:384] <= 32'h01E44703;
            reg_val_0_80000000[16][447:416] <= 32'h01D44683;
            reg_val_0_80000000[16][479:448] <= 32'h40E4D733;
            reg_val_0_80000000[16][511:480] <= 32'h033707B3;
            reg_val_0_80000000[17][31:0] <= 32'h40F487B3;
            reg_val_0_80000000[17][63:32] <= 32'h06068063;
            reg_val_0_80000000[17][95:64] <= 32'h01F44683;
            reg_val_0_80000000[17][127:96] <= 32'h40D7D6B3;
            reg_val_0_80000000[17][159:128] <= 32'h032688B3;
            reg_val_0_80000000[17][191:160] <= 32'h0145AE03;
            reg_val_0_80000000[17][223:192] <= 32'h0105A303;
            reg_val_0_80000000[17][255:224] <= 32'h00C5A603;
            reg_val_0_80000000[17][287:256] <= 32'h00442803;
            reg_val_0_80000000[17][319:288] <= 32'h00842503;
            reg_val_0_80000000[17][351:320] <= 32'h00148493;
            reg_val_0_80000000[17][383:352] <= 32'h01C70733;
            reg_val_0_80000000[17][415:384] <= 32'h006686B3;
            reg_val_0_80000000[17][447:416] <= 32'h411787B3;
            reg_val_0_80000000[17][479:448] <= 32'h00C78633;
            reg_val_0_80000000[17][511:480] <= 32'h000800E7;
            reg_val_0_80000000[18][31:0] <= 32'h029A0663;
            reg_val_0_80000000[18][63:32] <= 32'h00042583;
            reg_val_0_80000000[18][95:64] <= 32'h01C44783;
            reg_val_0_80000000[18][127:96] <= 32'hFA0792E3;
            reg_val_0_80000000[18][159:128] <= 32'h0334C733;
            reg_val_0_80000000[18][191:160] <= 32'h01D44683;
            reg_val_0_80000000[18][223:192] <= 32'h033707B3;
            reg_val_0_80000000[18][255:224] <= 32'h40F487B3;
            reg_val_0_80000000[18][287:256] <= 32'hFA0694E3;
            reg_val_0_80000000[18][319:288] <= 32'h0327C6B3;
            reg_val_0_80000000[18][351:320] <= 32'hFA9FF06F;
            reg_val_0_80000000[18][383:352] <= 32'h01842703;
            reg_val_0_80000000[18][415:384] <= 32'h00000793;
            reg_val_0_80000000[18][447:416] <= 32'h00E7C06B;
            reg_val_0_80000000[18][479:448] <= 32'h01C12083;
            reg_val_0_80000000[18][511:480] <= 32'h01812403;
            reg_val_0_80000000[19][31:0] <= 32'h01412483;
            reg_val_0_80000000[19][63:32] <= 32'h01012903;
            reg_val_0_80000000[19][95:64] <= 32'h00C12983;
            reg_val_0_80000000[19][127:96] <= 32'h00812A03;
            reg_val_0_80000000[19][159:128] <= 32'h02010113;
            reg_val_0_80000000[19][191:160] <= 32'h00008067;
            reg_val_0_80000000[19][223:192] <= 32'hCC502773;
            reg_val_0_80000000[19][255:224] <= 32'hCC2027F3;
            reg_val_0_80000000[19][287:256] <= 32'h00271693;
            reg_val_0_80000000[19][319:288] <= 32'h00001717;
            reg_val_0_80000000[19][351:320] <= 32'hF5C70713;
            reg_val_0_80000000[19][383:352] <= 32'h00D70733;
            reg_val_0_80000000[19][415:384] <= 32'h00072503;
            reg_val_0_80000000[19][447:416] <= 32'h00052583;
            reg_val_0_80000000[19][479:448] <= 32'h00C52683;
            reg_val_0_80000000[19][511:480] <= 32'h01C54703;
            reg_val_0_80000000[20][31:0] <= 32'h0005A883;
            reg_val_0_80000000[20][63:32] <= 32'h0045A603;
            reg_val_0_80000000[20][95:64] <= 32'h00D787B3;
            reg_val_0_80000000[20][127:96] <= 32'h02C88633;
            reg_val_0_80000000[20][159:128] <= 32'h04070863;
            reg_val_0_80000000[20][191:160] <= 32'h01E54703;
            reg_val_0_80000000[20][223:192] <= 32'h01D54683;
            reg_val_0_80000000[20][255:224] <= 32'h40E7D733;
            reg_val_0_80000000[20][287:256] <= 32'h02C70633;
            reg_val_0_80000000[20][319:288] <= 32'h40C787B3;
            reg_val_0_80000000[20][351:320] <= 32'h04068663;
            reg_val_0_80000000[20][383:352] <= 32'h01F54683;
            reg_val_0_80000000[20][415:384] <= 32'h40D7D833;
            reg_val_0_80000000[20][447:416] <= 32'h0105A683;
            reg_val_0_80000000[20][479:448] <= 32'h0145AE03;
            reg_val_0_80000000[20][511:480] <= 32'h00C5A603;
            reg_val_0_80000000[21][31:0] <= 32'h00D806B3;
            reg_val_0_80000000[21][63:32] <= 32'h03180833;
            reg_val_0_80000000[21][95:64] <= 32'h00452303;
            reg_val_0_80000000[21][127:96] <= 32'h00852503;
            reg_val_0_80000000[21][159:128] <= 32'h01C70733;
            reg_val_0_80000000[21][191:160] <= 32'h410787B3;
            reg_val_0_80000000[21][223:192] <= 32'h00C78633;
            reg_val_0_80000000[21][255:224] <= 32'h00030067;
            reg_val_0_80000000[21][287:256] <= 32'h02C7C733;
            reg_val_0_80000000[21][319:288] <= 32'h01D54683;
            reg_val_0_80000000[21][351:320] <= 32'h02C70633;
            reg_val_0_80000000[21][383:352] <= 32'h40C787B3;
            reg_val_0_80000000[21][415:384] <= 32'hFA069EE3;
            reg_val_0_80000000[21][447:416] <= 32'h0317C833;
            reg_val_0_80000000[21][479:448] <= 32'hFBDFF06F;
            reg_val_0_80000000[21][511:480] <= 32'hFF010113;
            reg_val_0_80000000[22][31:0] <= 32'h00112623;
            reg_val_0_80000000[22][63:32] <= 32'hFFF00793;
            reg_val_0_80000000[22][95:64] <= 32'h0007806B;
            reg_val_0_80000000[22][127:96] <= 32'hE11FF0EF;
            reg_val_0_80000000[22][159:128] <= 32'hCC3027F3;
            reg_val_0_80000000[22][191:160] <= 32'h0017B793;
            reg_val_0_80000000[22][223:192] <= 32'h0007806B;
            reg_val_0_80000000[22][255:224] <= 32'h00C12083;
            reg_val_0_80000000[22][287:256] <= 32'h01010113;
            reg_val_0_80000000[22][319:288] <= 32'h00008067;
            reg_val_0_80000000[22][351:320] <= 32'hFD010113;
            reg_val_0_80000000[22][383:352] <= 32'h02112623;
            reg_val_0_80000000[22][415:384] <= 32'h02812423;
            reg_val_0_80000000[22][447:416] <= 32'h02912223;
            reg_val_0_80000000[22][479:448] <= 32'h03212023;
            reg_val_0_80000000[22][511:480] <= 32'hFC2026F3;
            reg_val_0_80000000[23][31:0] <= 32'hFC1028F3;
            reg_val_0_80000000[23][63:32] <= 32'hFC0024F3;
            reg_val_0_80000000[23][95:64] <= 32'hCC5027F3;
            reg_val_0_80000000[23][127:96] <= 32'h01F00713;
            reg_val_0_80000000[23][159:128] <= 32'h08F74863;
            reg_val_0_80000000[23][191:160] <= 32'h03148833;
            reg_val_0_80000000[23][223:192] <= 32'h00100713;
            reg_val_0_80000000[23][255:224] <= 32'h00A85463;
            reg_val_0_80000000[23][287:256] <= 32'h03054733;
            reg_val_0_80000000[23][319:288] <= 32'h08E6CA63;
            reg_val_0_80000000[23][351:320] <= 32'h06E7DC63;
            reg_val_0_80000000[23][383:352] <= 32'hFFF68693;
            reg_val_0_80000000[23][415:384] <= 32'h02E54333;
            reg_val_0_80000000[23][447:416] <= 32'h00030813;
            reg_val_0_80000000[23][479:448] <= 32'h00F69663;
            reg_val_0_80000000[23][511:480] <= 32'h02E56533;
            reg_val_0_80000000[24][31:0] <= 32'h00650833;
            reg_val_0_80000000[24][63:32] <= 32'h02984933;
            reg_val_0_80000000[24][95:64] <= 32'h02986433;
            reg_val_0_80000000[24][127:96] <= 32'h07194C63;
            reg_val_0_80000000[24][159:128] <= 32'h00100513;
            reg_val_0_80000000[24][191:160] <= 32'h031946B3;
            reg_val_0_80000000[24][223:192] <= 32'h00068663;
            reg_val_0_80000000[24][255:224] <= 32'h00068513;
            reg_val_0_80000000[24][287:256] <= 32'h031966B3;
            reg_val_0_80000000[24][319:288] <= 32'h00001717;
            reg_val_0_80000000[24][351:320] <= 32'hE1C70713;
            reg_val_0_80000000[24][383:352] <= 32'h00B12423;
            reg_val_0_80000000[24][415:384] <= 32'h00C12623;
            reg_val_0_80000000[24][447:416] <= 32'h00A12A23;
            reg_val_0_80000000[24][479:448] <= 32'h00D12C23;
            reg_val_0_80000000[24][511:480] <= 32'h00012E23;
            reg_val_0_80000000[25][31:0] <= 32'h02F30333;
            reg_val_0_80000000[25][63:32] <= 32'h00279793;
            reg_val_0_80000000[25][95:64] <= 32'h00F707B3;
            reg_val_0_80000000[25][127:96] <= 32'h00810713;
            reg_val_0_80000000[25][159:128] <= 32'h00E7A023;
            reg_val_0_80000000[25][191:160] <= 32'h00612823;
            reg_val_0_80000000[25][223:192] <= 32'h03204C63;
            reg_val_0_80000000[25][255:224] <= 32'h06041663;
            reg_val_0_80000000[25][287:256] <= 32'h02C12083;
            reg_val_0_80000000[25][319:288] <= 32'h02812403;
            reg_val_0_80000000[25][351:320] <= 32'h02412483;
            reg_val_0_80000000[25][383:352] <= 32'h02012903;
            reg_val_0_80000000[25][415:384] <= 32'h03010113;
            reg_val_0_80000000[25][447:416] <= 32'h00008067;
            reg_val_0_80000000[25][479:448] <= 32'h00068713;
            reg_val_0_80000000[25][511:480] <= 32'hF6E7C8E3;
            reg_val_0_80000000[26][31:0] <= 32'hFE1FF06F;
            reg_val_0_80000000[26][63:32] <= 32'h00000693;
            reg_val_0_80000000[26][95:64] <= 32'h00100513;
            reg_val_0_80000000[26][127:96] <= 32'hF99FF06F;
            reg_val_0_80000000[26][159:128] <= 32'h00090793;
            reg_val_0_80000000[26][191:160] <= 32'h0128D463;
            reg_val_0_80000000[26][223:192] <= 32'h00088793;
            reg_val_0_80000000[26][255:224] <= 32'h00F12E23;
            reg_val_0_80000000[26][287:256] <= 32'h00000717;
            reg_val_0_80000000[26][319:288] <= 32'hCD070713;
            reg_val_0_80000000[26][351:320] <= 32'h00E7906B;
            reg_val_0_80000000[26][383:352] <= 32'hFFF00793;
            reg_val_0_80000000[26][415:384] <= 32'h0007806B;
            reg_val_0_80000000[26][447:416] <= 32'hBD9FF0EF;
            reg_val_0_80000000[26][479:448] <= 32'hCC3027F3;
            reg_val_0_80000000[26][511:480] <= 32'h0017B793;
            reg_val_0_80000000[27][31:0] <= 32'h0007806B;
            reg_val_0_80000000[27][63:32] <= 32'hF8040EE3;
            reg_val_0_80000000[27][95:64] <= 32'h029904B3;
            reg_val_0_80000000[27][127:96] <= 32'h00100913;
            reg_val_0_80000000[27][159:128] <= 32'h00891833;
            reg_val_0_80000000[27][191:160] <= 32'hFFF80813;
            reg_val_0_80000000[27][223:192] <= 32'h00912823;
            reg_val_0_80000000[27][255:224] <= 32'h0008006B;
            reg_val_0_80000000[27][287:256] <= 32'hC61FF0EF;
            reg_val_0_80000000[27][319:288] <= 32'h0009006B;
            reg_val_0_80000000[27][351:320] <= 32'h02C12083;
            reg_val_0_80000000[27][383:352] <= 32'h02812403;
            reg_val_0_80000000[27][415:384] <= 32'h02412483;
            reg_val_0_80000000[27][447:416] <= 32'h02012903;
            reg_val_0_80000000[27][479:448] <= 32'h03010113;
            reg_val_0_80000000[27][511:480] <= 32'h00008067;
            reg_val_0_80000000[28][31:0] <= 32'hFD010113;
            reg_val_0_80000000[28][63:32] <= 32'h02112623;
            reg_val_0_80000000[28][95:64] <= 32'h02812423;
            reg_val_0_80000000[28][127:96] <= 32'h02912223;
            reg_val_0_80000000[28][159:128] <= 32'h03212023;
            reg_val_0_80000000[28][191:160] <= 32'hFC2028F3;
            reg_val_0_80000000[28][223:192] <= 32'hFC102373;
            reg_val_0_80000000[28][255:224] <= 32'hFC0024F3;
            reg_val_0_80000000[28][287:256] <= 32'hCC5027F3;
            reg_val_0_80000000[28][319:288] <= 32'h01F00713;
            reg_val_0_80000000[28][351:320] <= 32'h0EF74663;
            reg_val_0_80000000[28][383:352] <= 32'h00052E03;
            reg_val_0_80000000[28][415:384] <= 32'h00452683;
            reg_val_0_80000000[28][447:416] <= 32'h00852803;
            reg_val_0_80000000[28][479:448] <= 32'h02930EB3;
            reg_val_0_80000000[28][511:480] <= 32'h00100713;
            reg_val_0_80000000[29][31:0] <= 32'h02DE06B3;
            reg_val_0_80000000[29][63:32] <= 32'h03068833;
            reg_val_0_80000000[29][95:64] <= 32'h010ED463;
            reg_val_0_80000000[29][127:96] <= 32'h03D84733;
            reg_val_0_80000000[29][159:128] <= 32'h0CE8CE63;
            reg_val_0_80000000[29][191:160] <= 32'h0CE7D063;
            reg_val_0_80000000[29][223:192] <= 32'hFFF88893;
            reg_val_0_80000000[29][255:224] <= 32'h02E84F33;
            reg_val_0_80000000[29][287:256] <= 32'h000F0413;
            reg_val_0_80000000[29][319:288] <= 32'h00F89663;
            reg_val_0_80000000[29][351:320] <= 32'h02E86733;
            reg_val_0_80000000[29][383:352] <= 32'h01E70433;
            reg_val_0_80000000[29][415:384] <= 32'h02944933;
            reg_val_0_80000000[29][447:416] <= 32'h02946433;
            reg_val_0_80000000[29][479:448] <= 32'h0C694063;
            reg_val_0_80000000[29][511:480] <= 32'h00100293;
            reg_val_0_80000000[30][31:0] <= 32'h02694FB3;
            reg_val_0_80000000[30][63:32] <= 32'h000F8663;
            reg_val_0_80000000[30][95:64] <= 32'h000F8293;
            reg_val_0_80000000[30][127:96] <= 32'h02696FB3;
            reg_val_0_80000000[30][159:128] <= 32'hD006F7D3;
            reg_val_0_80000000[30][191:160] <= 32'hFFFE0893;
            reg_val_0_80000000[30][223:192] <= 32'hFFF68E93;
            reg_val_0_80000000[30][255:224] <= 32'hE0078853;
            reg_val_0_80000000[30][287:256] <= 32'hD00E77D3;
            reg_val_0_80000000[30][319:288] <= 32'h00DEF6B3;
            reg_val_0_80000000[30][351:320] <= 32'h01C8FE33;
            reg_val_0_80000000[30][383:352] <= 32'hE0078753;
            reg_val_0_80000000[30][415:384] <= 32'h41785813;
            reg_val_0_80000000[30][447:416] <= 32'h00001897;
            reg_val_0_80000000[30][479:448] <= 32'hC8C88893;
            reg_val_0_80000000[30][511:480] <= 32'h41775713;
            reg_val_0_80000000[31][31:0] <= 32'h0016B693;
            reg_val_0_80000000[31][63:32] <= 32'h001E3E13;
            reg_val_0_80000000[31][95:64] <= 32'hF8180813;
            reg_val_0_80000000[31][127:96] <= 32'hF8170713;
            reg_val_0_80000000[31][159:128] <= 32'h00A12023;
            reg_val_0_80000000[31][191:160] <= 32'h00B12223;
            reg_val_0_80000000[31][223:192] <= 32'h00C12423;
            reg_val_0_80000000[31][255:224] <= 32'h00512823;
            reg_val_0_80000000[31][287:256] <= 32'h01F12A23;
            reg_val_0_80000000[31][319:288] <= 32'h00012C23;
            reg_val_0_80000000[31][351:320] <= 32'h00D10E23;
            reg_val_0_80000000[31][383:352] <= 32'h01C10EA3;
            reg_val_0_80000000[31][415:384] <= 32'h01010F23;
            reg_val_0_80000000[31][447:416] <= 32'h00E10FA3;
            reg_val_0_80000000[31][479:448] <= 32'h02FF0F33;
            reg_val_0_80000000[31][511:480] <= 32'h00279793;
            reg_val_0_80000000[32][31:0] <= 32'h00F887B3;
            reg_val_0_80000000[32][63:32] <= 32'h0027A023;
            reg_val_0_80000000[32][95:64] <= 32'h01E12623;
            reg_val_0_80000000[32][127:96] <= 32'h03204C63;
            reg_val_0_80000000[32][159:128] <= 32'h06041663;
            reg_val_0_80000000[32][191:160] <= 32'h02C12083;
            reg_val_0_80000000[32][223:192] <= 32'h02812403;
            reg_val_0_80000000[32][255:224] <= 32'h02412483;
            reg_val_0_80000000[32][287:256] <= 32'h02012903;
            reg_val_0_80000000[32][319:288] <= 32'h03010113;
            reg_val_0_80000000[32][351:320] <= 32'h00008067;
            reg_val_0_80000000[32][383:352] <= 32'h00088713;
            reg_val_0_80000000[32][415:384] <= 32'hF2E7C4E3;
            reg_val_0_80000000[32][447:416] <= 32'hFE1FF06F;
            reg_val_0_80000000[32][479:448] <= 32'h00000F93;
            reg_val_0_80000000[32][511:480] <= 32'h00100293;
            reg_val_0_80000000[33][31:0] <= 32'hF51FF06F;
            reg_val_0_80000000[33][63:32] <= 32'h00090793;
            reg_val_0_80000000[33][95:64] <= 32'h01235463;
            reg_val_0_80000000[33][127:96] <= 32'h00030793;
            reg_val_0_80000000[33][159:128] <= 32'h00F12C23;
            reg_val_0_80000000[33][191:160] <= 32'h00000717;
            reg_val_0_80000000[33][223:192] <= 32'hD2870713;
            reg_val_0_80000000[33][255:224] <= 32'h00E7906B;
            reg_val_0_80000000[33][287:256] <= 32'hFFF00793;
            reg_val_0_80000000[33][319:288] <= 32'h0007806B;
            reg_val_0_80000000[33][351:320] <= 32'hB35FF0EF;
            reg_val_0_80000000[33][383:352] <= 32'hCC3027F3;
            reg_val_0_80000000[33][415:384] <= 32'h0017B793;
            reg_val_0_80000000[33][447:416] <= 32'h0007806B;
            reg_val_0_80000000[33][479:448] <= 32'hF8040EE3;
            reg_val_0_80000000[33][511:480] <= 32'h029904B3;
            reg_val_0_80000000[34][31:0] <= 32'h00100913;
            reg_val_0_80000000[34][63:32] <= 32'h00891433;
            reg_val_0_80000000[34][95:64] <= 32'hFFF40413;
            reg_val_0_80000000[34][127:96] <= 32'h00912623;
            reg_val_0_80000000[34][159:128] <= 32'h0004006B;
            reg_val_0_80000000[34][191:160] <= 32'hC45FF0EF;
            reg_val_0_80000000[34][223:192] <= 32'h0009006B;
            reg_val_0_80000000[34][255:224] <= 32'h02C12083;
            reg_val_0_80000000[34][287:256] <= 32'h02812403;
            reg_val_0_80000000[34][319:288] <= 32'h02412483;
            reg_val_0_80000000[34][351:320] <= 32'h02012903;
            reg_val_0_80000000[34][383:352] <= 32'h03010113;
            reg_val_0_80000000[34][415:384] <= 32'h00008067;
            reg_val_0_80000000[34][447:416] <= 32'hFE810113;
            reg_val_0_80000000[34][479:448] <= 32'h00112A23;
            reg_val_0_80000000[34][511:480] <= 32'h01412823;
            reg_val_0_80000000[35][31:0] <= 32'h01312623;
            reg_val_0_80000000[35][63:32] <= 32'h01212423;
            reg_val_0_80000000[35][95:64] <= 32'h00912223;
            reg_val_0_80000000[35][127:96] <= 32'h00812023;
            reg_val_0_80000000[35][159:128] <= 32'h00050A13;
            reg_val_0_80000000[35][191:160] <= 32'h00058993;
            reg_val_0_80000000[35][223:192] <= 32'hFC002973;
            reg_val_0_80000000[35][255:224] <= 32'hCC0024F3;
            reg_val_0_80000000[35][287:256] <= 32'h00000413;
            reg_val_0_80000000[35][319:288] <= 32'h409402B3;
            reg_val_0_80000000[35][351:320] <= 32'h0012B313;
            reg_val_0_80000000[35][383:352] <= 32'h0003206B;
            reg_val_0_80000000[35][415:384] <= 32'h00029663;
            reg_val_0_80000000[35][447:416] <= 32'h00098513;
            reg_val_0_80000000[35][479:448] <= 32'h000A00E7;
            reg_val_0_80000000[35][511:480] <= 32'h0000306B;
            reg_val_0_80000000[36][31:0] <= 32'h00140413;
            reg_val_0_80000000[36][63:32] <= 32'hFF2440E3;
            reg_val_0_80000000[36][95:64] <= 32'h01412083;
            reg_val_0_80000000[36][127:96] <= 32'h01012A03;
            reg_val_0_80000000[36][159:128] <= 32'h00C12983;
            reg_val_0_80000000[36][191:160] <= 32'h00812903;
            reg_val_0_80000000[36][223:192] <= 32'h00412483;
            reg_val_0_80000000[36][255:224] <= 32'h00012403;
            reg_val_0_80000000[36][287:256] <= 32'h01810113;
            reg_val_0_80000000[36][319:288] <= 32'h00008067;
            reg_val_0_80000000[36][351:320] <= 32'hFFF00513;
            reg_val_0_80000000[36][383:352] <= 32'h00008067;
            reg_val_0_80000000[36][415:384] <= 32'hFFF00513;
            reg_val_0_80000000[36][447:416] <= 32'h00008067;
            reg_val_0_80000000[36][479:448] <= 32'hFFF00513;
            reg_val_0_80000000[36][511:480] <= 32'h00008067;
            reg_val_0_80000000[37][31:0] <= 32'hFFF00513;
            reg_val_0_80000000[37][63:32] <= 32'h00008067;
            reg_val_0_80000000[37][95:64] <= 32'hFFF00513;
            reg_val_0_80000000[37][127:96] <= 32'h00008067;
            reg_val_0_80000000[37][159:128] <= 32'hFFF00513;
            reg_val_0_80000000[37][191:160] <= 32'h00008067;
            reg_val_0_80000000[37][223:192] <= 32'h00000513;
            reg_val_0_80000000[37][255:224] <= 32'h00008067;
            reg_val_0_80000000[37][287:256] <= 32'hFFF00513;
            reg_val_0_80000000[37][319:288] <= 32'h00008067;
            reg_val_0_80000000[37][351:320] <= 32'hFFF00513;
            reg_val_0_80000000[37][383:352] <= 32'h00008067;
            reg_val_0_80000000[37][415:384] <= 32'hFFF00513;
            reg_val_0_80000000[37][447:416] <= 32'h00008067;
            reg_val_0_80000000[37][479:448] <= 32'hFFF00513;
            reg_val_0_80000000[37][511:480] <= 32'h00008067;
            reg_val_0_80000000[38][31:0] <= 32'hFFF00513;
            reg_val_0_80000000[38][63:32] <= 32'h00008067;
            reg_val_0_80000000[38][95:64] <= 32'h00050593;
            reg_val_0_80000000[38][127:96] <= 32'h00000693;
            reg_val_0_80000000[38][159:128] <= 32'h00000613;
            reg_val_0_80000000[38][191:160] <= 32'h00000513;
            reg_val_0_80000000[38][223:192] <= 32'h2300006F;
            reg_val_0_80000000[38][255:224] <= 32'hFF010113;
            reg_val_0_80000000[38][287:256] <= 32'h00000593;
            reg_val_0_80000000[38][319:288] <= 32'h00812423;
            reg_val_0_80000000[38][351:320] <= 32'h00112623;
            reg_val_0_80000000[38][383:352] <= 32'h00050413;
            reg_val_0_80000000[38][415:384] <= 32'h2B4000EF;
            reg_val_0_80000000[38][447:416] <= 32'h800017B7;
            reg_val_0_80000000[38][479:448] <= 32'h4387A503;
            reg_val_0_80000000[38][511:480] <= 32'h03C52783;
            reg_val_0_80000000[39][31:0] <= 32'h00078463;
            reg_val_0_80000000[39][63:32] <= 32'h000780E7;
            reg_val_0_80000000[39][95:64] <= 32'h00040513;
            reg_val_0_80000000[39][127:96] <= 32'hEC8FF0EF;
            reg_val_0_80000000[39][159:128] <= 32'h00A5C7B3;
            reg_val_0_80000000[39][191:160] <= 32'h0037F793;
            reg_val_0_80000000[39][223:192] <= 32'h00C508B3;
            reg_val_0_80000000[39][255:224] <= 32'h06079263;
            reg_val_0_80000000[39][287:256] <= 32'h00300793;
            reg_val_0_80000000[39][319:288] <= 32'h04C7FE63;
            reg_val_0_80000000[39][351:320] <= 32'h00357793;
            reg_val_0_80000000[39][383:352] <= 32'h00050713;
            reg_val_0_80000000[39][415:384] <= 32'h06079863;
            reg_val_0_80000000[39][447:416] <= 32'hFFC8F613;
            reg_val_0_80000000[39][479:448] <= 32'hFE060793;
            reg_val_0_80000000[39][511:480] <= 32'h08F76C63;
            reg_val_0_80000000[40][31:0] <= 32'h02C77C63;
            reg_val_0_80000000[40][63:32] <= 32'h00058693;
            reg_val_0_80000000[40][95:64] <= 32'h00070793;
            reg_val_0_80000000[40][127:96] <= 32'h0006A803;
            reg_val_0_80000000[40][159:128] <= 32'h00478793;
            reg_val_0_80000000[40][191:160] <= 32'h00468693;
            reg_val_0_80000000[40][223:192] <= 32'hFF07AE23;
            reg_val_0_80000000[40][255:224] <= 32'hFEC7E8E3;
            reg_val_0_80000000[40][287:256] <= 32'hFFF60793;
            reg_val_0_80000000[40][319:288] <= 32'h40E787B3;
            reg_val_0_80000000[40][351:320] <= 32'hFFC7F793;
            reg_val_0_80000000[40][383:352] <= 32'h00478793;
            reg_val_0_80000000[40][415:384] <= 32'h00F70733;
            reg_val_0_80000000[40][447:416] <= 32'h00F585B3;
            reg_val_0_80000000[40][479:448] <= 32'h01176863;
            reg_val_0_80000000[40][511:480] <= 32'h00008067;
            reg_val_0_80000000[41][31:0] <= 32'h00050713;
            reg_val_0_80000000[41][63:32] <= 32'hFF157CE3;
            reg_val_0_80000000[41][95:64] <= 32'h0005C783;
            reg_val_0_80000000[41][127:96] <= 32'h00170713;
            reg_val_0_80000000[41][159:128] <= 32'h00158593;
            reg_val_0_80000000[41][191:160] <= 32'hFEF70FA3;
            reg_val_0_80000000[41][223:192] <= 32'hFF1768E3;
            reg_val_0_80000000[41][255:224] <= 32'h00008067;
            reg_val_0_80000000[41][287:256] <= 32'h0005C683;
            reg_val_0_80000000[41][319:288] <= 32'h00170713;
            reg_val_0_80000000[41][351:320] <= 32'h00377793;
            reg_val_0_80000000[41][383:352] <= 32'hFED70FA3;
            reg_val_0_80000000[41][415:384] <= 32'h00158593;
            reg_val_0_80000000[41][447:416] <= 32'hF80780E3;
            reg_val_0_80000000[41][479:448] <= 32'h0005C683;
            reg_val_0_80000000[41][511:480] <= 32'h00170713;
            reg_val_0_80000000[42][31:0] <= 32'h00377793;
            reg_val_0_80000000[42][63:32] <= 32'hFED70FA3;
            reg_val_0_80000000[42][95:64] <= 32'h00158593;
            reg_val_0_80000000[42][127:96] <= 32'hFC079AE3;
            reg_val_0_80000000[42][159:128] <= 32'hF65FF06F;
            reg_val_0_80000000[42][191:160] <= 32'h0045A683;
            reg_val_0_80000000[42][223:192] <= 32'h0005A283;
            reg_val_0_80000000[42][255:224] <= 32'h0085AF83;
            reg_val_0_80000000[42][287:256] <= 32'h00C5AF03;
            reg_val_0_80000000[42][319:288] <= 32'h0105AE83;
            reg_val_0_80000000[42][351:320] <= 32'h0145AE03;
            reg_val_0_80000000[42][383:352] <= 32'h0185A303;
            reg_val_0_80000000[42][415:384] <= 32'h01C5A803;
            reg_val_0_80000000[42][447:416] <= 32'h00D72223;
            reg_val_0_80000000[42][479:448] <= 32'h0205A683;
            reg_val_0_80000000[42][511:480] <= 32'h00572023;
            reg_val_0_80000000[43][31:0] <= 32'h01F72423;
            reg_val_0_80000000[43][63:32] <= 32'h01E72623;
            reg_val_0_80000000[43][95:64] <= 32'h01D72823;
            reg_val_0_80000000[43][127:96] <= 32'h01C72A23;
            reg_val_0_80000000[43][159:128] <= 32'h00672C23;
            reg_val_0_80000000[43][191:160] <= 32'h01072E23;
            reg_val_0_80000000[43][223:192] <= 32'h02D72023;
            reg_val_0_80000000[43][255:224] <= 32'h02470713;
            reg_val_0_80000000[43][287:256] <= 32'h02458593;
            reg_val_0_80000000[43][319:288] <= 32'hFAF768E3;
            reg_val_0_80000000[43][351:320] <= 32'hF19FF06F;
            reg_val_0_80000000[43][383:352] <= 32'h00F00313;
            reg_val_0_80000000[43][415:384] <= 32'h00050713;
            reg_val_0_80000000[43][447:416] <= 32'h02C37E63;
            reg_val_0_80000000[43][479:448] <= 32'h00F77793;
            reg_val_0_80000000[43][511:480] <= 32'h0A079063;
            reg_val_0_80000000[44][31:0] <= 32'h08059263;
            reg_val_0_80000000[44][63:32] <= 32'hFF067693;
            reg_val_0_80000000[44][95:64] <= 32'h00F67613;
            reg_val_0_80000000[44][127:96] <= 32'h00E686B3;
            reg_val_0_80000000[44][159:128] <= 32'h00B72023;
            reg_val_0_80000000[44][191:160] <= 32'h00B72223;
            reg_val_0_80000000[44][223:192] <= 32'h00B72423;
            reg_val_0_80000000[44][255:224] <= 32'h00B72623;
            reg_val_0_80000000[44][287:256] <= 32'h01070713;
            reg_val_0_80000000[44][319:288] <= 32'hFED766E3;
            reg_val_0_80000000[44][351:320] <= 32'h00061463;
            reg_val_0_80000000[44][383:352] <= 32'h00008067;
            reg_val_0_80000000[44][415:384] <= 32'h40C306B3;
            reg_val_0_80000000[44][447:416] <= 32'h00269693;
            reg_val_0_80000000[44][479:448] <= 32'h00000297;
            reg_val_0_80000000[44][511:480] <= 32'h005686B3;
            reg_val_0_80000000[45][31:0] <= 32'h00C68067;
            reg_val_0_80000000[45][63:32] <= 32'h00B70723;
            reg_val_0_80000000[45][95:64] <= 32'h00B706A3;
            reg_val_0_80000000[45][127:96] <= 32'h00B70623;
            reg_val_0_80000000[45][159:128] <= 32'h00B705A3;
            reg_val_0_80000000[45][191:160] <= 32'h00B70523;
            reg_val_0_80000000[45][223:192] <= 32'h00B704A3;
            reg_val_0_80000000[45][255:224] <= 32'h00B70423;
            reg_val_0_80000000[45][287:256] <= 32'h00B703A3;
            reg_val_0_80000000[45][319:288] <= 32'h00B70323;
            reg_val_0_80000000[45][351:320] <= 32'h00B702A3;
            reg_val_0_80000000[45][383:352] <= 32'h00B70223;
            reg_val_0_80000000[45][415:384] <= 32'h00B701A3;
            reg_val_0_80000000[45][447:416] <= 32'h00B70123;
            reg_val_0_80000000[45][479:448] <= 32'h00B700A3;
            reg_val_0_80000000[45][511:480] <= 32'h00B70023;
            reg_val_0_80000000[46][31:0] <= 32'h00008067;
            reg_val_0_80000000[46][63:32] <= 32'h0FF5F593;
            reg_val_0_80000000[46][95:64] <= 32'h00859693;
            reg_val_0_80000000[46][127:96] <= 32'h00D5E5B3;
            reg_val_0_80000000[46][159:128] <= 32'h01059693;
            reg_val_0_80000000[46][191:160] <= 32'h00D5E5B3;
            reg_val_0_80000000[46][223:192] <= 32'hF6DFF06F;
            reg_val_0_80000000[46][255:224] <= 32'h00279693;
            reg_val_0_80000000[46][287:256] <= 32'h00000297;
            reg_val_0_80000000[46][319:288] <= 32'h005686B3;
            reg_val_0_80000000[46][351:320] <= 32'h00008293;
            reg_val_0_80000000[46][383:352] <= 32'hFA0680E7;
            reg_val_0_80000000[46][415:384] <= 32'h00028093;
            reg_val_0_80000000[46][447:416] <= 32'hFF078793;
            reg_val_0_80000000[46][479:448] <= 32'h40F70733;
            reg_val_0_80000000[46][511:480] <= 32'h00F60633;
            reg_val_0_80000000[47][31:0] <= 32'hF6C378E3;
            reg_val_0_80000000[47][63:32] <= 32'hF3DFF06F;
            reg_val_0_80000000[47][95:64] <= 32'h800017B7;
            reg_val_0_80000000[47][127:96] <= 32'h4387A703;
            reg_val_0_80000000[47][159:128] <= 32'h14872783;
            reg_val_0_80000000[47][191:160] <= 32'h04078C63;
            reg_val_0_80000000[47][223:192] <= 32'h0047A703;
            reg_val_0_80000000[47][255:224] <= 32'h01F00813;
            reg_val_0_80000000[47][287:256] <= 32'h06E84E63;
            reg_val_0_80000000[47][319:288] <= 32'h00271813;
            reg_val_0_80000000[47][351:320] <= 32'h02050663;
            reg_val_0_80000000[47][383:352] <= 32'h01078333;
            reg_val_0_80000000[47][415:384] <= 32'h08C32423;
            reg_val_0_80000000[47][447:416] <= 32'h1887A883;
            reg_val_0_80000000[47][479:448] <= 32'h00100613;
            reg_val_0_80000000[47][511:480] <= 32'h00E61633;
            reg_val_0_80000000[48][31:0] <= 32'h00C8E8B3;
            reg_val_0_80000000[48][63:32] <= 32'h1917A423;
            reg_val_0_80000000[48][95:64] <= 32'h10D32423;
            reg_val_0_80000000[48][127:96] <= 32'h00200693;
            reg_val_0_80000000[48][159:128] <= 32'h02D50463;
            reg_val_0_80000000[48][191:160] <= 32'h00170713;
            reg_val_0_80000000[48][223:192] <= 32'h00E7A223;
            reg_val_0_80000000[48][255:224] <= 32'h010787B3;
            reg_val_0_80000000[48][287:256] <= 32'h00B7A423;
            reg_val_0_80000000[48][319:288] <= 32'h00000513;
            reg_val_0_80000000[48][351:320] <= 32'h00008067;
            reg_val_0_80000000[48][383:352] <= 32'h14C70793;
            reg_val_0_80000000[48][415:384] <= 32'h14F72423;
            reg_val_0_80000000[48][447:416] <= 32'hFA5FF06F;
            reg_val_0_80000000[48][479:448] <= 32'h18C7A683;
            reg_val_0_80000000[48][511:480] <= 32'h00170713;
            reg_val_0_80000000[49][31:0] <= 32'h00E7A223;
            reg_val_0_80000000[49][63:32] <= 32'h00C6E633;
            reg_val_0_80000000[49][95:64] <= 32'h18C7A623;
            reg_val_0_80000000[49][127:96] <= 32'h010787B3;
            reg_val_0_80000000[49][159:128] <= 32'h00B7A423;
            reg_val_0_80000000[49][191:160] <= 32'h00000513;
            reg_val_0_80000000[49][223:192] <= 32'h00008067;
            reg_val_0_80000000[49][255:224] <= 32'hFFF00513;
            reg_val_0_80000000[49][287:256] <= 32'h00008067;
            reg_val_0_80000000[49][319:288] <= 32'hFD010113;
            reg_val_0_80000000[49][351:320] <= 32'h800017B7;
            reg_val_0_80000000[49][383:352] <= 32'h01412C23;
            reg_val_0_80000000[49][415:384] <= 32'h4387AA03;
            reg_val_0_80000000[49][447:416] <= 32'h03212023;
            reg_val_0_80000000[49][479:448] <= 32'h02112623;
            reg_val_0_80000000[49][511:480] <= 32'h148A2903;
            reg_val_0_80000000[50][31:0] <= 32'h02812423;
            reg_val_0_80000000[50][63:32] <= 32'h02912223;
            reg_val_0_80000000[50][95:64] <= 32'h01312E23;
            reg_val_0_80000000[50][127:96] <= 32'h01512A23;
            reg_val_0_80000000[50][159:128] <= 32'h01612823;
            reg_val_0_80000000[50][191:160] <= 32'h01712623;
            reg_val_0_80000000[50][223:192] <= 32'h01812423;
            reg_val_0_80000000[50][255:224] <= 32'h04090063;
            reg_val_0_80000000[50][287:256] <= 32'h00050B13;
            reg_val_0_80000000[50][319:288] <= 32'h00058B93;
            reg_val_0_80000000[50][351:320] <= 32'h00100A93;
            reg_val_0_80000000[50][383:352] <= 32'hFFF00993;
            reg_val_0_80000000[50][415:384] <= 32'h00492483;
            reg_val_0_80000000[50][447:416] <= 32'hFFF48413;
            reg_val_0_80000000[50][479:448] <= 32'h02044263;
            reg_val_0_80000000[50][511:480] <= 32'h00249493;
            reg_val_0_80000000[51][31:0] <= 32'h009904B3;
            reg_val_0_80000000[51][63:32] <= 32'h040B8463;
            reg_val_0_80000000[51][95:64] <= 32'h1044A783;
            reg_val_0_80000000[51][127:96] <= 32'h05778063;
            reg_val_0_80000000[51][159:128] <= 32'hFFF40413;
            reg_val_0_80000000[51][191:160] <= 32'hFFC48493;
            reg_val_0_80000000[51][223:192] <= 32'hFF3416E3;
            reg_val_0_80000000[51][255:224] <= 32'h02C12083;
            reg_val_0_80000000[51][287:256] <= 32'h02812403;
            reg_val_0_80000000[51][319:288] <= 32'h02412483;
            reg_val_0_80000000[51][351:320] <= 32'h02012903;
            reg_val_0_80000000[51][383:352] <= 32'h01C12983;
            reg_val_0_80000000[51][415:384] <= 32'h01812A03;
            reg_val_0_80000000[51][447:416] <= 32'h01412A83;
            reg_val_0_80000000[51][479:448] <= 32'h01012B03;
            reg_val_0_80000000[51][511:480] <= 32'h00C12B83;
            reg_val_0_80000000[52][31:0] <= 32'h00812C03;
            reg_val_0_80000000[52][63:32] <= 32'h03010113;
            reg_val_0_80000000[52][95:64] <= 32'h00008067;
            reg_val_0_80000000[52][127:96] <= 32'h00492783;
            reg_val_0_80000000[52][159:128] <= 32'h0044A683;
            reg_val_0_80000000[52][191:160] <= 32'hFFF78793;
            reg_val_0_80000000[52][223:192] <= 32'h04878E63;
            reg_val_0_80000000[52][255:224] <= 32'h0004A223;
            reg_val_0_80000000[52][287:256] <= 32'hFA0688E3;
            reg_val_0_80000000[52][319:288] <= 32'h18892783;
            reg_val_0_80000000[52][351:320] <= 32'h008A9733;
            reg_val_0_80000000[52][383:352] <= 32'h00492C03;
            reg_val_0_80000000[52][415:384] <= 32'h00F777B3;
            reg_val_0_80000000[52][447:416] <= 32'h02079263;
            reg_val_0_80000000[52][479:448] <= 32'h000680E7;
            reg_val_0_80000000[52][511:480] <= 32'h00492703;
            reg_val_0_80000000[53][31:0] <= 32'h148A2783;
            reg_val_0_80000000[53][63:32] <= 32'h01871463;
            reg_val_0_80000000[53][95:64] <= 32'hF8F904E3;
            reg_val_0_80000000[53][127:96] <= 32'hF80788E3;
            reg_val_0_80000000[53][159:128] <= 32'h00078913;
            reg_val_0_80000000[53][191:160] <= 32'hF5DFF06F;
            reg_val_0_80000000[53][223:192] <= 32'h18C92783;
            reg_val_0_80000000[53][255:224] <= 32'h0844A583;
            reg_val_0_80000000[53][287:256] <= 32'h00F77733;
            reg_val_0_80000000[53][319:288] <= 32'h00071C63;
            reg_val_0_80000000[53][351:320] <= 32'h000B0513;
            reg_val_0_80000000[53][383:352] <= 32'h000680E7;
            reg_val_0_80000000[53][415:384] <= 32'hFCDFF06F;
            reg_val_0_80000000[53][447:416] <= 32'h00892223;
            reg_val_0_80000000[53][479:448] <= 32'hFA9FF06F;
            reg_val_0_80000000[53][511:480] <= 32'h00058513;
            reg_val_0_80000000[54][31:0] <= 32'h000680E7;
            reg_val_0_80000000[54][63:32] <= 32'hFB9FF06F;
            reg_val_0_80000000[54][95:64] <= 32'h00000010;
            reg_val_0_80000000[54][127:96] <= 32'h00000000;
            reg_val_0_80000000[54][159:128] <= 32'h00527A03;
            reg_val_0_80000000[54][191:160] <= 32'h01017C01;
            reg_val_0_80000000[54][223:192] <= 32'h00020D1B;
            reg_val_0_80000000[54][255:224] <= 32'h00000010;
            reg_val_0_80000000[54][287:256] <= 32'h00000018;
            reg_val_0_80000000[54][319:288] <= 32'hFFFFFB84;
            reg_val_0_80000000[54][351:320] <= 32'h00000008;
            reg_val_0_80000000[54][383:352] <= 32'h00000000;
            reg_val_0_80000000[54][415:384] <= 32'h00000010;
            reg_val_0_80000000[54][447:416] <= 32'h0000002C;
            reg_val_0_80000000[54][479:448] <= 32'hFFFFFB78;
            reg_val_0_80000000[54][511:480] <= 32'h00000008;
            reg_val_0_80000000[55][31:0] <= 32'h00000000;
            reg_val_0_80000000[55][63:32] <= 32'h00000010;
            reg_val_0_80000000[55][95:64] <= 32'h00000040;
            reg_val_0_80000000[55][127:96] <= 32'hFFFFFB6C;
            reg_val_0_80000000[55][159:128] <= 32'h00000008;
            reg_val_0_80000000[55][191:160] <= 32'h00000000;
            reg_val_0_80000000[55][223:192] <= 32'h00000010;
            reg_val_0_80000000[55][255:224] <= 32'h00000054;
            reg_val_0_80000000[55][287:256] <= 32'hFFFFFB60;
            reg_val_0_80000000[55][319:288] <= 32'h00000008;
            reg_val_0_80000000[55][351:320] <= 32'h00000000;
            reg_val_0_80000000[55][383:352] <= 32'h00000010;
            reg_val_0_80000000[55][415:384] <= 32'h00000068;
            reg_val_0_80000000[55][447:416] <= 32'hFFFFFB54;
            reg_val_0_80000000[55][479:448] <= 32'h00000008;
            reg_val_0_80000000[55][511:480] <= 32'h00000000;
            reg_val_0_80000000[56][31:0] <= 32'h00000010;
            reg_val_0_80000000[56][63:32] <= 32'h0000007C;
            reg_val_0_80000000[56][95:64] <= 32'hFFFFFB48;
            reg_val_0_80000000[56][127:96] <= 32'h00000008;
            reg_val_0_80000000[56][159:128] <= 32'h00000000;
            reg_val_0_80000000[56][191:160] <= 32'h00000010;
            reg_val_0_80000000[56][223:192] <= 32'h00000090;
            reg_val_0_80000000[56][255:224] <= 32'hFFFFFB3C;
            reg_val_0_80000000[56][287:256] <= 32'h00000008;
            reg_val_0_80000000[56][319:288] <= 32'h00000000;
            reg_val_0_80000000[56][351:320] <= 32'h00000010;
            reg_val_0_80000000[56][383:352] <= 32'h000000A4;
            reg_val_0_80000000[56][415:384] <= 32'hFFFFFB30;
            reg_val_0_80000000[56][447:416] <= 32'h00000008;
            reg_val_0_80000000[56][479:448] <= 32'h00000000;
            reg_val_0_80000000[56][511:480] <= 32'h00000010;
            reg_val_0_80000000[57][31:0] <= 32'h000000B8;
            reg_val_0_80000000[57][63:32] <= 32'hFFFFFB24;
            reg_val_0_80000000[57][95:64] <= 32'h00000008;
            reg_val_0_80000000[57][127:96] <= 32'h00000000;
            reg_val_0_80000000[57][159:128] <= 32'h00000010;
            reg_val_0_80000000[57][191:160] <= 32'h000000CC;
            reg_val_0_80000000[57][223:192] <= 32'hFFFFFB18;
            reg_val_0_80000000[57][255:224] <= 32'h00000008;
            reg_val_0_80000000[57][287:256] <= 32'h00000000;
            reg_val_0_80000000[57][319:288] <= 32'h00000010;
            reg_val_0_80000000[57][351:320] <= 32'h000000E0;
            reg_val_0_80000000[57][383:352] <= 32'hFFFFFB0C;
            reg_val_0_80000000[57][415:384] <= 32'h00000008;
            reg_val_0_80000000[57][447:416] <= 32'h00000000;
            reg_val_0_80000000[57][479:448] <= 32'h00000010;
            reg_val_0_80000000[57][511:480] <= 32'h000000F4;
            reg_val_0_80000000[58][31:0] <= 32'hFFFFFB00;
            reg_val_0_80000000[58][63:32] <= 32'h00000008;
            reg_val_0_80000000[58][95:64] <= 32'h00000000;
            // fill-in reset values:
            reg_val_0_80000000[58][127:96] <= 32'h00000000;
            reg_val_0_80000000[58][159:128] <= 32'h00000000;
            reg_val_0_80000000[58][191:160] <= 32'h00000000;
            reg_val_0_80000000[58][223:192] <= 32'h00000000;
            reg_val_0_80000000[58][255:224] <= 32'h00000000;
            reg_val_0_80000000[58][287:256] <= 32'h00000000;
            reg_val_0_80000000[58][319:288] <= 32'h00000000;
            reg_val_0_80000000[58][351:320] <= 32'h00000000;
            reg_val_0_80000000[58][383:352] <= 32'h00000000;
            reg_val_0_80000000[58][415:384] <= 32'h00000000;
            reg_val_0_80000000[58][447:416] <= 32'h00000000;
            reg_val_0_80000000[58][479:448] <= 32'h00000000;
            reg_val_0_80000000[58][511:480] <= 32'h00000000;
            reg_val_0_80000000[59][31:0] <= 32'h00000000;
            reg_val_0_80000000[59][63:32] <= 32'h00000000;
            reg_val_0_80000000[59][95:64] <= 32'h00000000;
            reg_val_0_80000000[59][127:96] <= 32'h00000000;
            reg_val_0_80000000[59][159:128] <= 32'h00000000;
            reg_val_0_80000000[59][191:160] <= 32'h00000000;
            reg_val_0_80000000[59][223:192] <= 32'h00000000;
            reg_val_0_80000000[59][255:224] <= 32'h00000000;
            reg_val_0_80000000[59][287:256] <= 32'h00000000;
            reg_val_0_80000000[59][319:288] <= 32'h00000000;
            reg_val_0_80000000[59][351:320] <= 32'h00000000;
            reg_val_0_80000000[59][383:352] <= 32'h00000000;
            reg_val_0_80000000[59][415:384] <= 32'h00000000;
            reg_val_0_80000000[59][447:416] <= 32'h00000000;
            reg_val_0_80000000[59][479:448] <= 32'h00000000;
            reg_val_0_80000000[59][511:480] <= 32'h00000000;
            reg_val_0_80000000[60][31:0] <= 32'h00000000;
            reg_val_0_80000000[60][63:32] <= 32'h00000000;
            reg_val_0_80000000[60][95:64] <= 32'h00000000;
            reg_val_0_80000000[60][127:96] <= 32'h00000000;
            reg_val_0_80000000[60][159:128] <= 32'h00000000;
            reg_val_0_80000000[60][191:160] <= 32'h00000000;
            reg_val_0_80000000[60][223:192] <= 32'h00000000;
            reg_val_0_80000000[60][255:224] <= 32'h00000000;
            reg_val_0_80000000[60][287:256] <= 32'h00000000;
            reg_val_0_80000000[60][319:288] <= 32'h00000000;
            reg_val_0_80000000[60][351:320] <= 32'h00000000;
            reg_val_0_80000000[60][383:352] <= 32'h00000000;
            reg_val_0_80000000[60][415:384] <= 32'h00000000;
            reg_val_0_80000000[60][447:416] <= 32'h00000000;
            reg_val_0_80000000[60][479:448] <= 32'h00000000;
            reg_val_0_80000000[60][511:480] <= 32'h00000000;
            reg_val_0_80000000[61][31:0] <= 32'h00000000;
            reg_val_0_80000000[61][63:32] <= 32'h00000000;
            reg_val_0_80000000[61][95:64] <= 32'h00000000;
            reg_val_0_80000000[61][127:96] <= 32'h00000000;
            reg_val_0_80000000[61][159:128] <= 32'h00000000;
            reg_val_0_80000000[61][191:160] <= 32'h00000000;
            reg_val_0_80000000[61][223:192] <= 32'h00000000;
            reg_val_0_80000000[61][255:224] <= 32'h00000000;
            reg_val_0_80000000[61][287:256] <= 32'h00000000;
            reg_val_0_80000000[61][319:288] <= 32'h00000000;
            reg_val_0_80000000[61][351:320] <= 32'h00000000;
            reg_val_0_80000000[61][383:352] <= 32'h00000000;
            reg_val_0_80000000[61][415:384] <= 32'h00000000;
            reg_val_0_80000000[61][447:416] <= 32'h00000000;
            reg_val_0_80000000[61][479:448] <= 32'h00000000;
            reg_val_0_80000000[61][511:480] <= 32'h00000000;
            reg_val_0_80000000[62][31:0] <= 32'h00000000;
            reg_val_0_80000000[62][63:32] <= 32'h00000000;
            reg_val_0_80000000[62][95:64] <= 32'h00000000;
            reg_val_0_80000000[62][127:96] <= 32'h00000000;
            reg_val_0_80000000[62][159:128] <= 32'h00000000;
            reg_val_0_80000000[62][191:160] <= 32'h00000000;
            reg_val_0_80000000[62][223:192] <= 32'h00000000;
            reg_val_0_80000000[62][255:224] <= 32'h00000000;
            reg_val_0_80000000[62][287:256] <= 32'h00000000;
            reg_val_0_80000000[62][319:288] <= 32'h00000000;
            reg_val_0_80000000[62][351:320] <= 32'h00000000;
            reg_val_0_80000000[62][383:352] <= 32'h00000000;
            reg_val_0_80000000[62][415:384] <= 32'h00000000;
            reg_val_0_80000000[62][447:416] <= 32'h00000000;
            reg_val_0_80000000[62][479:448] <= 32'h00000000;
            reg_val_0_80000000[62][511:480] <= 32'h00000000;
            reg_val_0_80000000[63][31:0] <= 32'h00000000;
            reg_val_0_80000000[63][63:32] <= 32'h00000000;
            reg_val_0_80000000[63][95:64] <= 32'h00000000;
            reg_val_0_80000000[63][127:96] <= 32'h00000000;
            reg_val_0_80000000[63][159:128] <= 32'h00000000;
            reg_val_0_80000000[63][191:160] <= 32'h00000000;
            reg_val_0_80000000[63][223:192] <= 32'h00000000;
            reg_val_0_80000000[63][255:224] <= 32'h00000000;
            reg_val_0_80000000[63][287:256] <= 32'h00000000;
            reg_val_0_80000000[63][319:288] <= 32'h00000000;
            reg_val_0_80000000[63][351:320] <= 32'h00000000;
            reg_val_0_80000000[63][383:352] <= 32'h00000000;
            reg_val_0_80000000[63][415:384] <= 32'h00000000;
            reg_val_0_80000000[63][447:416] <= 32'h00000000;
            reg_val_0_80000000[63][479:448] <= 32'h00000000;
            reg_val_0_80000000[63][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_0_80000000 = next_reg_val_0_80000000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_0_80000000
        // hold reg val by default
        for (int i = 0; i < 64; i++)
        begin
            next_reg_val_0_80000000[i] = reg_val_0_80000000[i];
        end
        // update reg val if wen
        if (wen_0_80000000)
        begin
            next_reg_val_0_80000000[wsel_0_80000000] = wdata_0_80000000;
        end
    end
    
    always_comb begin : READ_LOGIC_0_80000000
        // read val at rsel
        rdata_0_80000000 = reg_val_0_80000000[rsel_0_80000000];
    end
    
    // chunk 1
    logic wen_1_80001000;
    logic [1-1:0] wsel_1_80001000;
    // logic wsel_1_80001000;
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_1_80001000;
    logic [1-1:0] rsel_1_80001000;
    // logic rsel_1_80001000;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_1_80001000;
    
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_1_80001000 [2-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_1_80001000 [2-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_1_80001000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_1_80001000[0][31:0] <= 32'h8000007C;
            // fill-in reset values:
            reg_val_1_80001000[0][63:32] <= 32'h00000000;
            reg_val_1_80001000[0][95:64] <= 32'h00000000;
            reg_val_1_80001000[0][127:96] <= 32'h00000000;
            reg_val_1_80001000[0][159:128] <= 32'h00000000;
            reg_val_1_80001000[0][191:160] <= 32'h00000000;
            reg_val_1_80001000[0][223:192] <= 32'h00000000;
            reg_val_1_80001000[0][255:224] <= 32'h00000000;
            reg_val_1_80001000[0][287:256] <= 32'h00000000;
            reg_val_1_80001000[0][319:288] <= 32'h00000000;
            reg_val_1_80001000[0][351:320] <= 32'h00000000;
            reg_val_1_80001000[0][383:352] <= 32'h00000000;
            reg_val_1_80001000[0][415:384] <= 32'h00000000;
            reg_val_1_80001000[0][447:416] <= 32'h00000000;
            reg_val_1_80001000[0][479:448] <= 32'h00000000;
            reg_val_1_80001000[0][511:480] <= 32'h00000000;
            reg_val_1_80001000[1][63:32] <= 32'h00000000;
            reg_val_1_80001000[1][95:64] <= 32'h00000000;
            reg_val_1_80001000[1][127:96] <= 32'h00000000;
            reg_val_1_80001000[1][159:128] <= 32'h00000000;
            reg_val_1_80001000[1][191:160] <= 32'h00000000;
            reg_val_1_80001000[1][223:192] <= 32'h00000000;
            reg_val_1_80001000[1][255:224] <= 32'h00000000;
            reg_val_1_80001000[1][287:256] <= 32'h00000000;
            reg_val_1_80001000[1][319:288] <= 32'h00000000;
            reg_val_1_80001000[1][351:320] <= 32'h00000000;
            reg_val_1_80001000[1][383:352] <= 32'h00000000;
            reg_val_1_80001000[1][415:384] <= 32'h00000000;
            reg_val_1_80001000[1][447:416] <= 32'h00000000;
            reg_val_1_80001000[1][479:448] <= 32'h00000000;
            reg_val_1_80001000[1][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_1_80001000 = next_reg_val_1_80001000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_1_80001000
        // hold reg val by default
        for (int i = 0; i < 1; i++)
        begin
            next_reg_val_1_80001000[i] = reg_val_1_80001000[i];
        end
        // update reg val if wen
        if (wen_1_80001000)
        begin
            next_reg_val_1_80001000[wsel_1_80001000] = wdata_1_80001000;
        end
    end
    
    always_comb begin : READ_LOGIC_1_80001000
        // read val at rsel
        rdata_1_80001000 = reg_val_1_80001000[rsel_1_80001000];
    end
    
    // chunk 2
    logic wen_2_80001008;
    logic [5-1:0] wsel_2_80001008;
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_2_80001008;
    logic [5-1:0] rsel_2_80001008;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_2_80001008;
    
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_2_80001008 [32-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_2_80001008 [32-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_2_80001008
        if (reset)
        begin
            // enumerated reset values:
            reg_val_2_80001008[0][31:0] <= 32'h00000000;
            reg_val_2_80001008[0][63:32] <= 32'h00000000;
            reg_val_2_80001008[0][95:64] <= 32'h00000000;
            reg_val_2_80001008[0][127:96] <= 32'h800012FC;
            reg_val_2_80001008[0][159:128] <= 32'h80001364;
            reg_val_2_80001008[0][191:160] <= 32'h800013CC;
            reg_val_2_80001008[0][223:192] <= 32'h00000000;
            reg_val_2_80001008[0][255:224] <= 32'h00000000;
            reg_val_2_80001008[0][287:256] <= 32'h00000000;
            reg_val_2_80001008[0][319:288] <= 32'h00000000;
            reg_val_2_80001008[0][351:320] <= 32'h00000000;
            reg_val_2_80001008[0][383:352] <= 32'h00000000;
            reg_val_2_80001008[0][415:384] <= 32'h00000000;
            reg_val_2_80001008[0][447:416] <= 32'h00000000;
            reg_val_2_80001008[0][479:448] <= 32'h00000000;
            reg_val_2_80001008[0][511:480] <= 32'h00000000;
            reg_val_2_80001008[1][31:0] <= 32'h00000000;
            reg_val_2_80001008[1][63:32] <= 32'h00000000;
            reg_val_2_80001008[1][95:64] <= 32'h00000000;
            reg_val_2_80001008[1][127:96] <= 32'h00000000;
            reg_val_2_80001008[1][159:128] <= 32'h00000000;
            reg_val_2_80001008[1][191:160] <= 32'h00000000;
            reg_val_2_80001008[1][223:192] <= 32'h00000000;
            reg_val_2_80001008[1][255:224] <= 32'h00000000;
            reg_val_2_80001008[1][287:256] <= 32'h00000000;
            reg_val_2_80001008[1][319:288] <= 32'h00000000;
            reg_val_2_80001008[1][351:320] <= 32'h00000000;
            reg_val_2_80001008[1][383:352] <= 32'h00000000;
            reg_val_2_80001008[1][415:384] <= 32'h00000000;
            reg_val_2_80001008[1][447:416] <= 32'h00000000;
            reg_val_2_80001008[1][479:448] <= 32'h00000000;
            reg_val_2_80001008[1][511:480] <= 32'h00000000;
            reg_val_2_80001008[2][31:0] <= 32'h00000000;
            reg_val_2_80001008[2][63:32] <= 32'h00000000;
            reg_val_2_80001008[2][95:64] <= 32'h00000000;
            reg_val_2_80001008[2][127:96] <= 32'h00000000;
            reg_val_2_80001008[2][159:128] <= 32'h00000000;
            reg_val_2_80001008[2][191:160] <= 32'h00000000;
            reg_val_2_80001008[2][223:192] <= 32'h00000000;
            reg_val_2_80001008[2][255:224] <= 32'h00000000;
            reg_val_2_80001008[2][287:256] <= 32'h00000000;
            reg_val_2_80001008[2][319:288] <= 32'h00000000;
            reg_val_2_80001008[2][351:320] <= 32'h00000000;
            reg_val_2_80001008[2][383:352] <= 32'h00000000;
            reg_val_2_80001008[2][415:384] <= 32'h00000001;
            reg_val_2_80001008[2][447:416] <= 32'h00000000;
            reg_val_2_80001008[2][479:448] <= 32'hABCD330E;
            reg_val_2_80001008[2][511:480] <= 32'hE66D1234;
            reg_val_2_80001008[3][31:0] <= 32'h0005DEEC;
            reg_val_2_80001008[3][63:32] <= 32'h0000000B;
            reg_val_2_80001008[3][95:64] <= 32'h00000000;
            reg_val_2_80001008[3][127:96] <= 32'h00000000;
            reg_val_2_80001008[3][159:128] <= 32'h00000000;
            reg_val_2_80001008[3][191:160] <= 32'h00000000;
            reg_val_2_80001008[3][223:192] <= 32'h00000000;
            reg_val_2_80001008[3][255:224] <= 32'h00000000;
            reg_val_2_80001008[3][287:256] <= 32'h00000000;
            reg_val_2_80001008[3][319:288] <= 32'h00000000;
            reg_val_2_80001008[3][351:320] <= 32'h00000000;
            reg_val_2_80001008[3][383:352] <= 32'h00000000;
            reg_val_2_80001008[3][415:384] <= 32'h00000000;
            reg_val_2_80001008[3][447:416] <= 32'h00000000;
            reg_val_2_80001008[3][479:448] <= 32'h00000000;
            reg_val_2_80001008[3][511:480] <= 32'h00000000;
            reg_val_2_80001008[4][31:0] <= 32'h00000000;
            reg_val_2_80001008[4][63:32] <= 32'h00000000;
            reg_val_2_80001008[4][95:64] <= 32'h00000000;
            reg_val_2_80001008[4][127:96] <= 32'h00000000;
            reg_val_2_80001008[4][159:128] <= 32'h00000000;
            reg_val_2_80001008[4][191:160] <= 32'h00000000;
            reg_val_2_80001008[4][223:192] <= 32'h00000000;
            reg_val_2_80001008[4][255:224] <= 32'h00000000;
            reg_val_2_80001008[4][287:256] <= 32'h00000000;
            reg_val_2_80001008[4][319:288] <= 32'h00000000;
            reg_val_2_80001008[4][351:320] <= 32'h00000000;
            reg_val_2_80001008[4][383:352] <= 32'h00000000;
            reg_val_2_80001008[4][415:384] <= 32'h00000000;
            reg_val_2_80001008[4][447:416] <= 32'h00000000;
            reg_val_2_80001008[4][479:448] <= 32'h00000000;
            reg_val_2_80001008[4][511:480] <= 32'h00000000;
            reg_val_2_80001008[5][31:0] <= 32'h00000000;
            reg_val_2_80001008[5][63:32] <= 32'h00000000;
            reg_val_2_80001008[5][95:64] <= 32'h00000000;
            reg_val_2_80001008[5][127:96] <= 32'h00000000;
            reg_val_2_80001008[5][159:128] <= 32'h00000000;
            reg_val_2_80001008[5][191:160] <= 32'h00000000;
            reg_val_2_80001008[5][223:192] <= 32'h00000000;
            reg_val_2_80001008[5][255:224] <= 32'h00000000;
            reg_val_2_80001008[5][287:256] <= 32'h00000000;
            reg_val_2_80001008[5][319:288] <= 32'h00000000;
            reg_val_2_80001008[5][351:320] <= 32'h00000000;
            reg_val_2_80001008[5][383:352] <= 32'h00000000;
            reg_val_2_80001008[5][415:384] <= 32'h00000000;
            reg_val_2_80001008[5][447:416] <= 32'h00000000;
            reg_val_2_80001008[5][479:448] <= 32'h00000000;
            reg_val_2_80001008[5][511:480] <= 32'h00000000;
            reg_val_2_80001008[6][31:0] <= 32'h00000000;
            reg_val_2_80001008[6][63:32] <= 32'h00000000;
            reg_val_2_80001008[6][95:64] <= 32'h00000000;
            reg_val_2_80001008[6][127:96] <= 32'h00000000;
            reg_val_2_80001008[6][159:128] <= 32'h00000000;
            reg_val_2_80001008[6][191:160] <= 32'h00000000;
            reg_val_2_80001008[6][223:192] <= 32'h00000000;
            reg_val_2_80001008[6][255:224] <= 32'h00000000;
            reg_val_2_80001008[6][287:256] <= 32'h00000000;
            reg_val_2_80001008[6][319:288] <= 32'h00000000;
            reg_val_2_80001008[6][351:320] <= 32'h00000000;
            reg_val_2_80001008[6][383:352] <= 32'h00000000;
            reg_val_2_80001008[6][415:384] <= 32'h00000000;
            reg_val_2_80001008[6][447:416] <= 32'h00000000;
            reg_val_2_80001008[6][479:448] <= 32'h00000000;
            reg_val_2_80001008[6][511:480] <= 32'h00000000;
            reg_val_2_80001008[7][31:0] <= 32'h00000000;
            reg_val_2_80001008[7][63:32] <= 32'h00000000;
            reg_val_2_80001008[7][95:64] <= 32'h00000000;
            reg_val_2_80001008[7][127:96] <= 32'h00000000;
            reg_val_2_80001008[7][159:128] <= 32'h00000000;
            reg_val_2_80001008[7][191:160] <= 32'h00000000;
            reg_val_2_80001008[7][223:192] <= 32'h00000000;
            reg_val_2_80001008[7][255:224] <= 32'h00000000;
            reg_val_2_80001008[7][287:256] <= 32'h00000000;
            reg_val_2_80001008[7][319:288] <= 32'h00000000;
            reg_val_2_80001008[7][351:320] <= 32'h00000000;
            reg_val_2_80001008[7][383:352] <= 32'h00000000;
            reg_val_2_80001008[7][415:384] <= 32'h00000000;
            reg_val_2_80001008[7][447:416] <= 32'h00000000;
            reg_val_2_80001008[7][479:448] <= 32'h00000000;
            reg_val_2_80001008[7][511:480] <= 32'h00000000;
            reg_val_2_80001008[8][31:0] <= 32'h00000000;
            reg_val_2_80001008[8][63:32] <= 32'h00000000;
            reg_val_2_80001008[8][95:64] <= 32'h00000000;
            reg_val_2_80001008[8][127:96] <= 32'h00000000;
            reg_val_2_80001008[8][159:128] <= 32'h00000000;
            reg_val_2_80001008[8][191:160] <= 32'h00000000;
            reg_val_2_80001008[8][223:192] <= 32'h00000000;
            reg_val_2_80001008[8][255:224] <= 32'h00000000;
            reg_val_2_80001008[8][287:256] <= 32'h00000000;
            reg_val_2_80001008[8][319:288] <= 32'h00000000;
            reg_val_2_80001008[8][351:320] <= 32'h00000000;
            reg_val_2_80001008[8][383:352] <= 32'h00000000;
            reg_val_2_80001008[8][415:384] <= 32'h00000000;
            reg_val_2_80001008[8][447:416] <= 32'h00000000;
            reg_val_2_80001008[8][479:448] <= 32'h00000000;
            reg_val_2_80001008[8][511:480] <= 32'h00000000;
            reg_val_2_80001008[9][31:0] <= 32'h00000000;
            reg_val_2_80001008[9][63:32] <= 32'h00000000;
            reg_val_2_80001008[9][95:64] <= 32'h00000000;
            reg_val_2_80001008[9][127:96] <= 32'h00000000;
            reg_val_2_80001008[9][159:128] <= 32'h00000000;
            reg_val_2_80001008[9][191:160] <= 32'h00000000;
            reg_val_2_80001008[9][223:192] <= 32'h00000000;
            reg_val_2_80001008[9][255:224] <= 32'h00000000;
            reg_val_2_80001008[9][287:256] <= 32'h00000000;
            reg_val_2_80001008[9][319:288] <= 32'h00000000;
            reg_val_2_80001008[9][351:320] <= 32'h00000000;
            reg_val_2_80001008[9][383:352] <= 32'h00000000;
            reg_val_2_80001008[9][415:384] <= 32'h00000000;
            reg_val_2_80001008[9][447:416] <= 32'h00000000;
            reg_val_2_80001008[9][479:448] <= 32'h00000000;
            reg_val_2_80001008[9][511:480] <= 32'h00000000;
            reg_val_2_80001008[10][31:0] <= 32'h00000000;
            reg_val_2_80001008[10][63:32] <= 32'h00000000;
            reg_val_2_80001008[10][95:64] <= 32'h00000000;
            reg_val_2_80001008[10][127:96] <= 32'h00000000;
            reg_val_2_80001008[10][159:128] <= 32'h00000000;
            reg_val_2_80001008[10][191:160] <= 32'h00000000;
            reg_val_2_80001008[10][223:192] <= 32'h00000000;
            reg_val_2_80001008[10][255:224] <= 32'h00000000;
            reg_val_2_80001008[10][287:256] <= 32'h00000000;
            reg_val_2_80001008[10][319:288] <= 32'h00000000;
            reg_val_2_80001008[10][351:320] <= 32'h00000000;
            reg_val_2_80001008[10][383:352] <= 32'h00000000;
            reg_val_2_80001008[10][415:384] <= 32'h00000000;
            reg_val_2_80001008[10][447:416] <= 32'h00000000;
            reg_val_2_80001008[10][479:448] <= 32'h00000000;
            reg_val_2_80001008[10][511:480] <= 32'h00000000;
            reg_val_2_80001008[11][31:0] <= 32'h00000000;
            reg_val_2_80001008[11][63:32] <= 32'h00000000;
            reg_val_2_80001008[11][95:64] <= 32'h00000000;
            reg_val_2_80001008[11][127:96] <= 32'h00000000;
            reg_val_2_80001008[11][159:128] <= 32'h00000000;
            reg_val_2_80001008[11][191:160] <= 32'h00000000;
            reg_val_2_80001008[11][223:192] <= 32'h00000000;
            reg_val_2_80001008[11][255:224] <= 32'h00000000;
            reg_val_2_80001008[11][287:256] <= 32'h00000000;
            reg_val_2_80001008[11][319:288] <= 32'h00000000;
            reg_val_2_80001008[11][351:320] <= 32'h00000000;
            reg_val_2_80001008[11][383:352] <= 32'h00000000;
            reg_val_2_80001008[11][415:384] <= 32'h00000000;
            reg_val_2_80001008[11][447:416] <= 32'h00000000;
            reg_val_2_80001008[11][479:448] <= 32'h00000000;
            reg_val_2_80001008[11][511:480] <= 32'h00000000;
            reg_val_2_80001008[12][31:0] <= 32'h00000000;
            reg_val_2_80001008[12][63:32] <= 32'h00000000;
            reg_val_2_80001008[12][95:64] <= 32'h00000000;
            reg_val_2_80001008[12][127:96] <= 32'h00000000;
            reg_val_2_80001008[12][159:128] <= 32'h00000000;
            reg_val_2_80001008[12][191:160] <= 32'h00000000;
            reg_val_2_80001008[12][223:192] <= 32'h00000000;
            reg_val_2_80001008[12][255:224] <= 32'h00000000;
            reg_val_2_80001008[12][287:256] <= 32'h00000000;
            reg_val_2_80001008[12][319:288] <= 32'h00000000;
            reg_val_2_80001008[12][351:320] <= 32'h00000000;
            reg_val_2_80001008[12][383:352] <= 32'h00000000;
            reg_val_2_80001008[12][415:384] <= 32'h00000000;
            reg_val_2_80001008[12][447:416] <= 32'h00000000;
            reg_val_2_80001008[12][479:448] <= 32'h00000000;
            reg_val_2_80001008[12][511:480] <= 32'h00000000;
            reg_val_2_80001008[13][31:0] <= 32'h00000000;
            reg_val_2_80001008[13][63:32] <= 32'h00000000;
            reg_val_2_80001008[13][95:64] <= 32'h00000000;
            reg_val_2_80001008[13][127:96] <= 32'h00000000;
            reg_val_2_80001008[13][159:128] <= 32'h00000000;
            reg_val_2_80001008[13][191:160] <= 32'h00000000;
            reg_val_2_80001008[13][223:192] <= 32'h00000000;
            reg_val_2_80001008[13][255:224] <= 32'h00000000;
            reg_val_2_80001008[13][287:256] <= 32'h00000000;
            reg_val_2_80001008[13][319:288] <= 32'h00000000;
            reg_val_2_80001008[13][351:320] <= 32'h00000000;
            reg_val_2_80001008[13][383:352] <= 32'h00000000;
            reg_val_2_80001008[13][415:384] <= 32'h00000000;
            reg_val_2_80001008[13][447:416] <= 32'h00000000;
            reg_val_2_80001008[13][479:448] <= 32'h00000000;
            reg_val_2_80001008[13][511:480] <= 32'h00000000;
            reg_val_2_80001008[14][31:0] <= 32'h00000000;
            reg_val_2_80001008[14][63:32] <= 32'h00000000;
            reg_val_2_80001008[14][95:64] <= 32'h00000000;
            reg_val_2_80001008[14][127:96] <= 32'h00000000;
            reg_val_2_80001008[14][159:128] <= 32'h00000000;
            reg_val_2_80001008[14][191:160] <= 32'h00000000;
            reg_val_2_80001008[14][223:192] <= 32'h00000000;
            reg_val_2_80001008[14][255:224] <= 32'h00000000;
            reg_val_2_80001008[14][287:256] <= 32'h00000000;
            reg_val_2_80001008[14][319:288] <= 32'h00000000;
            reg_val_2_80001008[14][351:320] <= 32'h00000000;
            reg_val_2_80001008[14][383:352] <= 32'h00000000;
            reg_val_2_80001008[14][415:384] <= 32'h00000000;
            reg_val_2_80001008[14][447:416] <= 32'h00000000;
            reg_val_2_80001008[14][479:448] <= 32'h00000000;
            reg_val_2_80001008[14][511:480] <= 32'h00000000;
            reg_val_2_80001008[15][31:0] <= 32'h00000000;
            reg_val_2_80001008[15][63:32] <= 32'h00000000;
            reg_val_2_80001008[15][95:64] <= 32'h00000000;
            reg_val_2_80001008[15][127:96] <= 32'h00000000;
            reg_val_2_80001008[15][159:128] <= 32'h00000000;
            reg_val_2_80001008[15][191:160] <= 32'h00000000;
            reg_val_2_80001008[15][223:192] <= 32'h00000000;
            reg_val_2_80001008[15][255:224] <= 32'h00000000;
            reg_val_2_80001008[15][287:256] <= 32'h00000000;
            reg_val_2_80001008[15][319:288] <= 32'h00000000;
            reg_val_2_80001008[15][351:320] <= 32'h00000000;
            reg_val_2_80001008[15][383:352] <= 32'h00000000;
            reg_val_2_80001008[15][415:384] <= 32'h00000000;
            reg_val_2_80001008[15][447:416] <= 32'h00000000;
            reg_val_2_80001008[15][479:448] <= 32'h00000000;
            reg_val_2_80001008[15][511:480] <= 32'h00000000;
            reg_val_2_80001008[16][31:0] <= 32'h00000000;
            reg_val_2_80001008[16][63:32] <= 32'h00000000;
            reg_val_2_80001008[16][95:64] <= 32'h00000000;
            reg_val_2_80001008[16][127:96] <= 32'h00000000;
            reg_val_2_80001008[16][159:128] <= 32'h00000000;
            reg_val_2_80001008[16][191:160] <= 32'h00000000;
            reg_val_2_80001008[16][223:192] <= 32'h00000000;
            reg_val_2_80001008[16][255:224] <= 32'h00000000;
            reg_val_2_80001008[16][287:256] <= 32'h00000000;
            reg_val_2_80001008[16][319:288] <= 32'h00000000;
            reg_val_2_80001008[16][351:320] <= 32'h00000000;
            reg_val_2_80001008[16][383:352] <= 32'h00000000;
            reg_val_2_80001008[16][415:384] <= 32'h80001010;
            reg_val_2_80001008[16][447:416] <= 32'h80001010;
            // fill-in reset values:
            reg_val_2_80001008[16][479:448] <= 32'h00000000;
            reg_val_2_80001008[16][511:480] <= 32'h00000000;
            reg_val_2_80001008[17][31:0] <= 32'h00000000;
            reg_val_2_80001008[17][63:32] <= 32'h00000000;
            reg_val_2_80001008[17][95:64] <= 32'h00000000;
            reg_val_2_80001008[17][127:96] <= 32'h00000000;
            reg_val_2_80001008[17][159:128] <= 32'h00000000;
            reg_val_2_80001008[17][191:160] <= 32'h00000000;
            reg_val_2_80001008[17][223:192] <= 32'h00000000;
            reg_val_2_80001008[17][255:224] <= 32'h00000000;
            reg_val_2_80001008[17][287:256] <= 32'h00000000;
            reg_val_2_80001008[17][319:288] <= 32'h00000000;
            reg_val_2_80001008[17][351:320] <= 32'h00000000;
            reg_val_2_80001008[17][383:352] <= 32'h00000000;
            reg_val_2_80001008[17][415:384] <= 32'h00000000;
            reg_val_2_80001008[17][447:416] <= 32'h00000000;
            reg_val_2_80001008[17][479:448] <= 32'h00000000;
            reg_val_2_80001008[17][511:480] <= 32'h00000000;
            reg_val_2_80001008[18][31:0] <= 32'h00000000;
            reg_val_2_80001008[18][63:32] <= 32'h00000000;
            reg_val_2_80001008[18][95:64] <= 32'h00000000;
            reg_val_2_80001008[18][127:96] <= 32'h00000000;
            reg_val_2_80001008[18][159:128] <= 32'h00000000;
            reg_val_2_80001008[18][191:160] <= 32'h00000000;
            reg_val_2_80001008[18][223:192] <= 32'h00000000;
            reg_val_2_80001008[18][255:224] <= 32'h00000000;
            reg_val_2_80001008[18][287:256] <= 32'h00000000;
            reg_val_2_80001008[18][319:288] <= 32'h00000000;
            reg_val_2_80001008[18][351:320] <= 32'h00000000;
            reg_val_2_80001008[18][383:352] <= 32'h00000000;
            reg_val_2_80001008[18][415:384] <= 32'h00000000;
            reg_val_2_80001008[18][447:416] <= 32'h00000000;
            reg_val_2_80001008[18][479:448] <= 32'h00000000;
            reg_val_2_80001008[18][511:480] <= 32'h00000000;
            reg_val_2_80001008[19][31:0] <= 32'h00000000;
            reg_val_2_80001008[19][63:32] <= 32'h00000000;
            reg_val_2_80001008[19][95:64] <= 32'h00000000;
            reg_val_2_80001008[19][127:96] <= 32'h00000000;
            reg_val_2_80001008[19][159:128] <= 32'h00000000;
            reg_val_2_80001008[19][191:160] <= 32'h00000000;
            reg_val_2_80001008[19][223:192] <= 32'h00000000;
            reg_val_2_80001008[19][255:224] <= 32'h00000000;
            reg_val_2_80001008[19][287:256] <= 32'h00000000;
            reg_val_2_80001008[19][319:288] <= 32'h00000000;
            reg_val_2_80001008[19][351:320] <= 32'h00000000;
            reg_val_2_80001008[19][383:352] <= 32'h00000000;
            reg_val_2_80001008[19][415:384] <= 32'h00000000;
            reg_val_2_80001008[19][447:416] <= 32'h00000000;
            reg_val_2_80001008[19][479:448] <= 32'h00000000;
            reg_val_2_80001008[19][511:480] <= 32'h00000000;
            reg_val_2_80001008[20][31:0] <= 32'h00000000;
            reg_val_2_80001008[20][63:32] <= 32'h00000000;
            reg_val_2_80001008[20][95:64] <= 32'h00000000;
            reg_val_2_80001008[20][127:96] <= 32'h00000000;
            reg_val_2_80001008[20][159:128] <= 32'h00000000;
            reg_val_2_80001008[20][191:160] <= 32'h00000000;
            reg_val_2_80001008[20][223:192] <= 32'h00000000;
            reg_val_2_80001008[20][255:224] <= 32'h00000000;
            reg_val_2_80001008[20][287:256] <= 32'h00000000;
            reg_val_2_80001008[20][319:288] <= 32'h00000000;
            reg_val_2_80001008[20][351:320] <= 32'h00000000;
            reg_val_2_80001008[20][383:352] <= 32'h00000000;
            reg_val_2_80001008[20][415:384] <= 32'h00000000;
            reg_val_2_80001008[20][447:416] <= 32'h00000000;
            reg_val_2_80001008[20][479:448] <= 32'h00000000;
            reg_val_2_80001008[20][511:480] <= 32'h00000000;
            reg_val_2_80001008[21][31:0] <= 32'h00000000;
            reg_val_2_80001008[21][63:32] <= 32'h00000000;
            reg_val_2_80001008[21][95:64] <= 32'h00000000;
            reg_val_2_80001008[21][127:96] <= 32'h00000000;
            reg_val_2_80001008[21][159:128] <= 32'h00000000;
            reg_val_2_80001008[21][191:160] <= 32'h00000000;
            reg_val_2_80001008[21][223:192] <= 32'h00000000;
            reg_val_2_80001008[21][255:224] <= 32'h00000000;
            reg_val_2_80001008[21][287:256] <= 32'h00000000;
            reg_val_2_80001008[21][319:288] <= 32'h00000000;
            reg_val_2_80001008[21][351:320] <= 32'h00000000;
            reg_val_2_80001008[21][383:352] <= 32'h00000000;
            reg_val_2_80001008[21][415:384] <= 32'h00000000;
            reg_val_2_80001008[21][447:416] <= 32'h00000000;
            reg_val_2_80001008[21][479:448] <= 32'h00000000;
            reg_val_2_80001008[21][511:480] <= 32'h00000000;
            reg_val_2_80001008[22][31:0] <= 32'h00000000;
            reg_val_2_80001008[22][63:32] <= 32'h00000000;
            reg_val_2_80001008[22][95:64] <= 32'h00000000;
            reg_val_2_80001008[22][127:96] <= 32'h00000000;
            reg_val_2_80001008[22][159:128] <= 32'h00000000;
            reg_val_2_80001008[22][191:160] <= 32'h00000000;
            reg_val_2_80001008[22][223:192] <= 32'h00000000;
            reg_val_2_80001008[22][255:224] <= 32'h00000000;
            reg_val_2_80001008[22][287:256] <= 32'h00000000;
            reg_val_2_80001008[22][319:288] <= 32'h00000000;
            reg_val_2_80001008[22][351:320] <= 32'h00000000;
            reg_val_2_80001008[22][383:352] <= 32'h00000000;
            reg_val_2_80001008[22][415:384] <= 32'h00000000;
            reg_val_2_80001008[22][447:416] <= 32'h00000000;
            reg_val_2_80001008[22][479:448] <= 32'h00000000;
            reg_val_2_80001008[22][511:480] <= 32'h00000000;
            reg_val_2_80001008[23][31:0] <= 32'h00000000;
            reg_val_2_80001008[23][63:32] <= 32'h00000000;
            reg_val_2_80001008[23][95:64] <= 32'h00000000;
            reg_val_2_80001008[23][127:96] <= 32'h00000000;
            reg_val_2_80001008[23][159:128] <= 32'h00000000;
            reg_val_2_80001008[23][191:160] <= 32'h00000000;
            reg_val_2_80001008[23][223:192] <= 32'h00000000;
            reg_val_2_80001008[23][255:224] <= 32'h00000000;
            reg_val_2_80001008[23][287:256] <= 32'h00000000;
            reg_val_2_80001008[23][319:288] <= 32'h00000000;
            reg_val_2_80001008[23][351:320] <= 32'h00000000;
            reg_val_2_80001008[23][383:352] <= 32'h00000000;
            reg_val_2_80001008[23][415:384] <= 32'h00000000;
            reg_val_2_80001008[23][447:416] <= 32'h00000000;
            reg_val_2_80001008[23][479:448] <= 32'h00000000;
            reg_val_2_80001008[23][511:480] <= 32'h00000000;
            reg_val_2_80001008[24][31:0] <= 32'h00000000;
            reg_val_2_80001008[24][63:32] <= 32'h00000000;
            reg_val_2_80001008[24][95:64] <= 32'h00000000;
            reg_val_2_80001008[24][127:96] <= 32'h00000000;
            reg_val_2_80001008[24][159:128] <= 32'h00000000;
            reg_val_2_80001008[24][191:160] <= 32'h00000000;
            reg_val_2_80001008[24][223:192] <= 32'h00000000;
            reg_val_2_80001008[24][255:224] <= 32'h00000000;
            reg_val_2_80001008[24][287:256] <= 32'h00000000;
            reg_val_2_80001008[24][319:288] <= 32'h00000000;
            reg_val_2_80001008[24][351:320] <= 32'h00000000;
            reg_val_2_80001008[24][383:352] <= 32'h00000000;
            reg_val_2_80001008[24][415:384] <= 32'h00000000;
            reg_val_2_80001008[24][447:416] <= 32'h00000000;
            reg_val_2_80001008[24][479:448] <= 32'h00000000;
            reg_val_2_80001008[24][511:480] <= 32'h00000000;
            reg_val_2_80001008[25][31:0] <= 32'h00000000;
            reg_val_2_80001008[25][63:32] <= 32'h00000000;
            reg_val_2_80001008[25][95:64] <= 32'h00000000;
            reg_val_2_80001008[25][127:96] <= 32'h00000000;
            reg_val_2_80001008[25][159:128] <= 32'h00000000;
            reg_val_2_80001008[25][191:160] <= 32'h00000000;
            reg_val_2_80001008[25][223:192] <= 32'h00000000;
            reg_val_2_80001008[25][255:224] <= 32'h00000000;
            reg_val_2_80001008[25][287:256] <= 32'h00000000;
            reg_val_2_80001008[25][319:288] <= 32'h00000000;
            reg_val_2_80001008[25][351:320] <= 32'h00000000;
            reg_val_2_80001008[25][383:352] <= 32'h00000000;
            reg_val_2_80001008[25][415:384] <= 32'h00000000;
            reg_val_2_80001008[25][447:416] <= 32'h00000000;
            reg_val_2_80001008[25][479:448] <= 32'h00000000;
            reg_val_2_80001008[25][511:480] <= 32'h00000000;
            reg_val_2_80001008[26][31:0] <= 32'h00000000;
            reg_val_2_80001008[26][63:32] <= 32'h00000000;
            reg_val_2_80001008[26][95:64] <= 32'h00000000;
            reg_val_2_80001008[26][127:96] <= 32'h00000000;
            reg_val_2_80001008[26][159:128] <= 32'h00000000;
            reg_val_2_80001008[26][191:160] <= 32'h00000000;
            reg_val_2_80001008[26][223:192] <= 32'h00000000;
            reg_val_2_80001008[26][255:224] <= 32'h00000000;
            reg_val_2_80001008[26][287:256] <= 32'h00000000;
            reg_val_2_80001008[26][319:288] <= 32'h00000000;
            reg_val_2_80001008[26][351:320] <= 32'h00000000;
            reg_val_2_80001008[26][383:352] <= 32'h00000000;
            reg_val_2_80001008[26][415:384] <= 32'h00000000;
            reg_val_2_80001008[26][447:416] <= 32'h00000000;
            reg_val_2_80001008[26][479:448] <= 32'h00000000;
            reg_val_2_80001008[26][511:480] <= 32'h00000000;
            reg_val_2_80001008[27][31:0] <= 32'h00000000;
            reg_val_2_80001008[27][63:32] <= 32'h00000000;
            reg_val_2_80001008[27][95:64] <= 32'h00000000;
            reg_val_2_80001008[27][127:96] <= 32'h00000000;
            reg_val_2_80001008[27][159:128] <= 32'h00000000;
            reg_val_2_80001008[27][191:160] <= 32'h00000000;
            reg_val_2_80001008[27][223:192] <= 32'h00000000;
            reg_val_2_80001008[27][255:224] <= 32'h00000000;
            reg_val_2_80001008[27][287:256] <= 32'h00000000;
            reg_val_2_80001008[27][319:288] <= 32'h00000000;
            reg_val_2_80001008[27][351:320] <= 32'h00000000;
            reg_val_2_80001008[27][383:352] <= 32'h00000000;
            reg_val_2_80001008[27][415:384] <= 32'h00000000;
            reg_val_2_80001008[27][447:416] <= 32'h00000000;
            reg_val_2_80001008[27][479:448] <= 32'h00000000;
            reg_val_2_80001008[27][511:480] <= 32'h00000000;
            reg_val_2_80001008[28][31:0] <= 32'h00000000;
            reg_val_2_80001008[28][63:32] <= 32'h00000000;
            reg_val_2_80001008[28][95:64] <= 32'h00000000;
            reg_val_2_80001008[28][127:96] <= 32'h00000000;
            reg_val_2_80001008[28][159:128] <= 32'h00000000;
            reg_val_2_80001008[28][191:160] <= 32'h00000000;
            reg_val_2_80001008[28][223:192] <= 32'h00000000;
            reg_val_2_80001008[28][255:224] <= 32'h00000000;
            reg_val_2_80001008[28][287:256] <= 32'h00000000;
            reg_val_2_80001008[28][319:288] <= 32'h00000000;
            reg_val_2_80001008[28][351:320] <= 32'h00000000;
            reg_val_2_80001008[28][383:352] <= 32'h00000000;
            reg_val_2_80001008[28][415:384] <= 32'h00000000;
            reg_val_2_80001008[28][447:416] <= 32'h00000000;
            reg_val_2_80001008[28][479:448] <= 32'h00000000;
            reg_val_2_80001008[28][511:480] <= 32'h00000000;
            reg_val_2_80001008[29][31:0] <= 32'h00000000;
            reg_val_2_80001008[29][63:32] <= 32'h00000000;
            reg_val_2_80001008[29][95:64] <= 32'h00000000;
            reg_val_2_80001008[29][127:96] <= 32'h00000000;
            reg_val_2_80001008[29][159:128] <= 32'h00000000;
            reg_val_2_80001008[29][191:160] <= 32'h00000000;
            reg_val_2_80001008[29][223:192] <= 32'h00000000;
            reg_val_2_80001008[29][255:224] <= 32'h00000000;
            reg_val_2_80001008[29][287:256] <= 32'h00000000;
            reg_val_2_80001008[29][319:288] <= 32'h00000000;
            reg_val_2_80001008[29][351:320] <= 32'h00000000;
            reg_val_2_80001008[29][383:352] <= 32'h00000000;
            reg_val_2_80001008[29][415:384] <= 32'h00000000;
            reg_val_2_80001008[29][447:416] <= 32'h00000000;
            reg_val_2_80001008[29][479:448] <= 32'h00000000;
            reg_val_2_80001008[29][511:480] <= 32'h00000000;
            reg_val_2_80001008[30][31:0] <= 32'h00000000;
            reg_val_2_80001008[30][63:32] <= 32'h00000000;
            reg_val_2_80001008[30][95:64] <= 32'h00000000;
            reg_val_2_80001008[30][127:96] <= 32'h00000000;
            reg_val_2_80001008[30][159:128] <= 32'h00000000;
            reg_val_2_80001008[30][191:160] <= 32'h00000000;
            reg_val_2_80001008[30][223:192] <= 32'h00000000;
            reg_val_2_80001008[30][255:224] <= 32'h00000000;
            reg_val_2_80001008[30][287:256] <= 32'h00000000;
            reg_val_2_80001008[30][319:288] <= 32'h00000000;
            reg_val_2_80001008[30][351:320] <= 32'h00000000;
            reg_val_2_80001008[30][383:352] <= 32'h00000000;
            reg_val_2_80001008[30][415:384] <= 32'h00000000;
            reg_val_2_80001008[30][447:416] <= 32'h00000000;
            reg_val_2_80001008[30][479:448] <= 32'h00000000;
            reg_val_2_80001008[30][511:480] <= 32'h00000000;
            reg_val_2_80001008[31][31:0] <= 32'h00000000;
            reg_val_2_80001008[31][63:32] <= 32'h00000000;
            reg_val_2_80001008[31][95:64] <= 32'h00000000;
            reg_val_2_80001008[31][127:96] <= 32'h00000000;
            reg_val_2_80001008[31][159:128] <= 32'h00000000;
            reg_val_2_80001008[31][191:160] <= 32'h00000000;
            reg_val_2_80001008[31][223:192] <= 32'h00000000;
            reg_val_2_80001008[31][255:224] <= 32'h00000000;
            reg_val_2_80001008[31][287:256] <= 32'h00000000;
            reg_val_2_80001008[31][319:288] <= 32'h00000000;
            reg_val_2_80001008[31][351:320] <= 32'h00000000;
            reg_val_2_80001008[31][383:352] <= 32'h00000000;
            reg_val_2_80001008[31][415:384] <= 32'h00000000;
            reg_val_2_80001008[31][447:416] <= 32'h00000000;
            reg_val_2_80001008[31][479:448] <= 32'h00000000;
            reg_val_2_80001008[31][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_2_80001008 = next_reg_val_2_80001008;
        end
    end
    
    always_comb begin : WRITE_LOGIC_2_80001008
        // hold reg val by default
        for (int i = 0; i < 32; i++)
        begin
            next_reg_val_2_80001008[i] = reg_val_2_80001008[i];
        end
        // update reg val if wen
        if (wen_2_80001008)
        begin
            next_reg_val_2_80001008[wsel_2_80001008] = wdata_2_80001008;
        end
    end
    
    always_comb begin : READ_LOGIC_2_80001008
        // read val at rsel
        rdata_2_80001008 = reg_val_2_80001008[rsel_2_80001008];
    end
    
    // need reg file/chunk selection signal
    logic [2-1:0] chunk_sel;

    // addr hashing logic
    always_comb begin : ADDR_HASHING_LOGIC
        // default as address not out of bounds
        tb_addr_out_of_bounds = 1'b0;
        
        // bad address assertion:
        assert (
            (26'b10000000000000000000000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000000000000 + 64) ||
            (26'b10000000000000000001000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000001000000 + 1) ||
            (26'b10000000000000000001000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000001000000 + 32)
        ) else begin
            $display("mem request at address 0x%h = 0b%b not available in chunks", mem_req_addr, mem_req_addr);
            tb_addr_out_of_bounds = 1'b1;
        end
        
        // bit = 1 branch
        if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 20] == 1'b1)
        begin
            if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 26] == 1'b0)
            begin
                // select chunk @ 0x80001000
                chunk_sel = 1;
            end
            else if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 26] == 1'b0)
            begin
                // select chunk @ 0x80001008
                chunk_sel = 2;
            end
        end
        // bit = 0 branch
        else if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 20] == 1'b0)
        begin
            // select chunk @ 0x80000000
            chunk_sel = 0;
        end
        else
        begin
            $display("error: got to else in high-level branch");
            tb_addr_out_of_bounds = 1'b1;
        end
        
        // hardwired outputs:
        // hardwiring for chunk 0
        wsel_0_80000000 = mem_req_addr[6-1 : 0];
        wdata_0_80000000 = mem_req_data;
        rsel_0_80000000 = mem_req_addr[6-1 : 0];
        // hardwiring for chunk 1
        wsel_1_80001000 = mem_req_addr[1-1 : 0];
        wdata_1_80001000 = mem_req_data;
        rsel_1_80001000 = mem_req_addr[1-1 : 0];
        // hardwiring for chunk 2
        wsel_2_80001008 = mem_req_addr[5-1 : 0];
        wdata_2_80001008 = mem_req_data;
        rsel_2_80001008 = mem_req_addr[5-1 : 0];
        
        // default outputs:
        mem_rsp_data = {16{32'hdeadbeef}};
        // chunk wen's:
        wen_0_80000000 = 1'b0;
        wen_1_80001000 = 1'b0;
        wen_2_80001008 = 1'b0;
        
        // case for routing to diff reg file chunks
        casez (chunk_sel)
        
            // select chunk 0 @ 0x80000000
            0:
            begin
                // write routing
                wen_0_80000000 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_0_80000000;
            end
        
            // select chunk 1 @ 0x80001000
            1:
            begin
                // write routing
                wen_1_80001000 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_1_80001000;
            end
        
            // select chunk 2 @ 0x80001008
            2:
            begin
                // write routing
                wen_2_80001008 = mem_req_rw;
                // read routing
                mem_rsp_data = rdata_2_80001008;
            end
        
            // shouldn't get here
            default:
            begin
                $display("error: got to default in chunk_sel case");
                mem_rsp_data = {16{32'hdeadbeef}};
                tb_addr_out_of_bounds = 1'b1;
            end
        endcase
    end

    // other combinational logic for memory interface
    always_comb begin : OTHER_MEM_COMB_LOGIC

        // mem_req_ready = 1'b1;           // always ready for request
        mem_rsp_valid = mem_req_valid;  // read ready immediately
            // update to buffer to later clock cycle
                // along with data read value

        mem_rsp_tag = mem_req_tag;      // match req immediately
    end

    // delayed mem_req_ready signals
    parameter MEM_REQ_READY_DELAY = 15;
    logic [MEM_REQ_READY_DELAY-1:0] mem_req_ready_reg, next_mem_req_ready_reg; 

    // delayed mem_req_ready reg logic
    always_ff @ (posedge clk) begin : MEM_REQ_READY_REG_LOGIC
    
        if (reset)
        begin
            mem_req_ready_reg = '0;
        end
        else
        begin
            mem_req_ready_reg = next_mem_req_ready_reg;
        end
    end

    // delayed mem_req_ready delay next state logic
    always_comb begin : MEM_REQ_READY_DELAY_NEXT_STATE_LOGIC

        next_mem_req_ready_reg = {mem_req_ready_reg[MEM_REQ_READY_DELAY-2:0], 1'b1};    // shift 1 left
        mem_req_ready = mem_req_ready_reg[MEM_REQ_READY_DELAY-1];                       // msb of shifter
    end

    // NOTES:
    // don't know what to do with: 
        // mem_req_byteen
        // busy

endmodule

