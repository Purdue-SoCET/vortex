// `ifndef LOCAL_MEM_DEFINE
// `define LOCAL_MEM_DEFINE

// // temporary hardcoded values 
// `define VX_MEM_BYTEEN_WIDTH     1
// `define VX_MEM_ADDR_WIDTH       32
// `define VX_MEM_DATA_WIDTH       32
// `define VX_MEM_TAG_WIDTH        4     

// `endif
