/*
    socet115 / zlagpaca@purdue.edu
    Zach Lagpacan

    module for faking memory with basic register file which can interface with Vortex memory interface
*/

// temporary include to have defined vals
// `include "local_mem.vh"
`include "../include/VX_define.vh"
// `include "VX_define.vh"

module local_mem #(
)(
    // seq
    input clk, reset,

    // Memory Request:
    // vortex outputs
    input logic                             mem_req_valid,
    input logic                             mem_req_rw,
    input logic [`VX_MEM_BYTEEN_WIDTH-1:0]  mem_req_byteen, // 64 (512 / 8)
    input logic [`VX_MEM_ADDR_WIDTH-1:0]    mem_req_addr,   // 26
    input logic [`VX_MEM_DATA_WIDTH-1:0]    mem_req_data,   // 512
    input logic [`VX_MEM_TAG_WIDTH-1:0]     mem_req_tag,    // 56 (55 for SM disabled)
    // vortex inputs
    output logic                            mem_req_ready,

    // Memory response:
    // vortex inputs
    output logic                            mem_rsp_valid,        
    output logic [`VX_MEM_DATA_WIDTH-1:0]   mem_rsp_data,   // 512
    output logic [`VX_MEM_TAG_WIDTH-1:0]    mem_rsp_tag,    // 56 (55 for SM disabled)
    // vortex outputs
    input logic                             mem_rsp_ready,

    // Status:
    // vortex outputs
    input logic                             busy,

    // tb:
    output logic                            tb_addr_out_of_bounds
);
    // register file instances
    
    // chunk 0
    logic wen_0_80000000;
    
    // block selection within reg file
    logic [5-1:0] wsel_0_80000000;
    logic [5-1:0] rsel_0_80000000;
    
    // lock-sized reg file write input and read output
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_0_80000000;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_0_80000000;
    
    // 2D register file
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_0_80000000 [32-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_0_80000000 [32-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_0_80000000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_0_80000000[0][31:0] <= 32'h0480006F;
            reg_val_0_80000000[0][63:32] <= 32'h34202F73;
            reg_val_0_80000000[0][95:64] <= 32'h00800F93;
            reg_val_0_80000000[0][127:96] <= 32'h03FF0863;
            reg_val_0_80000000[0][159:128] <= 32'h00900F93;
            reg_val_0_80000000[0][191:160] <= 32'h03FF0463;
            reg_val_0_80000000[0][223:192] <= 32'h00B00F93;
            reg_val_0_80000000[0][255:224] <= 32'h03FF0063;
            reg_val_0_80000000[0][287:256] <= 32'h00000F13;
            reg_val_0_80000000[0][319:288] <= 32'h000F0463;
            reg_val_0_80000000[0][351:320] <= 32'h000F0067;
            reg_val_0_80000000[0][383:352] <= 32'h34202F73;
            reg_val_0_80000000[0][415:384] <= 32'h000F5463;
            reg_val_0_80000000[0][447:416] <= 32'h0040006F;
            reg_val_0_80000000[0][479:448] <= 32'h5391E193;
            reg_val_0_80000000[0][511:480] <= 32'h00001F17;
            reg_val_0_80000000[1][31:0] <= 32'hFC3F2223;
            reg_val_0_80000000[1][63:32] <= 32'hFF9FF06F;
            reg_val_0_80000000[1][95:64] <= 32'h00000093;
            reg_val_0_80000000[1][127:96] <= 32'h00000113;
            reg_val_0_80000000[1][159:128] <= 32'h00000193;
            reg_val_0_80000000[1][191:160] <= 32'h00000213;
            reg_val_0_80000000[1][223:192] <= 32'h00000293;
            reg_val_0_80000000[1][255:224] <= 32'h00000313;
            reg_val_0_80000000[1][287:256] <= 32'h00000393;
            reg_val_0_80000000[1][319:288] <= 32'h00000413;
            reg_val_0_80000000[1][351:320] <= 32'h00000493;
            reg_val_0_80000000[1][383:352] <= 32'h00000513;
            reg_val_0_80000000[1][415:384] <= 32'h00000593;
            reg_val_0_80000000[1][447:416] <= 32'h00000613;
            reg_val_0_80000000[1][479:448] <= 32'h00000693;
            reg_val_0_80000000[1][511:480] <= 32'h00000713;
            reg_val_0_80000000[2][31:0] <= 32'h00000793;
            reg_val_0_80000000[2][63:32] <= 32'h00000813;
            reg_val_0_80000000[2][95:64] <= 32'h00000893;
            reg_val_0_80000000[2][127:96] <= 32'h00000913;
            reg_val_0_80000000[2][159:128] <= 32'h00000993;
            reg_val_0_80000000[2][191:160] <= 32'h00000A13;
            reg_val_0_80000000[2][223:192] <= 32'h00000A93;
            reg_val_0_80000000[2][255:224] <= 32'h00000B13;
            reg_val_0_80000000[2][287:256] <= 32'h00000B93;
            reg_val_0_80000000[2][319:288] <= 32'h00000C13;
            reg_val_0_80000000[2][351:320] <= 32'h00000C93;
            reg_val_0_80000000[2][383:352] <= 32'h00000D13;
            reg_val_0_80000000[2][415:384] <= 32'h00000D93;
            reg_val_0_80000000[2][447:416] <= 32'h00000E13;
            reg_val_0_80000000[2][479:448] <= 32'h00000E93;
            reg_val_0_80000000[2][511:480] <= 32'h00000F13;
            reg_val_0_80000000[3][31:0] <= 32'h00000F93;
            reg_val_0_80000000[3][63:32] <= 32'hF1402573;
            reg_val_0_80000000[3][95:64] <= 32'h00051063;
            reg_val_0_80000000[3][127:96] <= 32'h00000297;
            reg_val_0_80000000[3][159:128] <= 32'h01028293;
            reg_val_0_80000000[3][191:160] <= 32'h30529073;
            reg_val_0_80000000[3][223:192] <= 32'h18005073;
            reg_val_0_80000000[3][255:224] <= 32'h00000297;
            reg_val_0_80000000[3][287:256] <= 32'h02028293;
            reg_val_0_80000000[3][319:288] <= 32'h30529073;
            reg_val_0_80000000[3][351:320] <= 32'h800002B7;
            reg_val_0_80000000[3][383:352] <= 32'hFFF28293;
            reg_val_0_80000000[3][415:384] <= 32'h3B029073;
            reg_val_0_80000000[3][447:416] <= 32'h01F00293;
            reg_val_0_80000000[3][479:448] <= 32'h3A029073;
            reg_val_0_80000000[3][511:480] <= 32'h30405073;
            reg_val_0_80000000[4][31:0] <= 32'h00000297;
            reg_val_0_80000000[4][63:32] <= 32'h01428293;
            reg_val_0_80000000[4][95:64] <= 32'h30529073;
            reg_val_0_80000000[4][127:96] <= 32'h30205073;
            reg_val_0_80000000[4][159:128] <= 32'h30305073;
            reg_val_0_80000000[4][191:160] <= 32'h00000193;
            reg_val_0_80000000[4][223:192] <= 32'h00000297;
            reg_val_0_80000000[4][255:224] <= 32'hEEC28293;
            reg_val_0_80000000[4][287:256] <= 32'h30529073;
            reg_val_0_80000000[4][319:288] <= 32'h00100513;
            reg_val_0_80000000[4][351:320] <= 32'h01F51513;
            reg_val_0_80000000[4][383:352] <= 32'h00054C63;
            reg_val_0_80000000[4][415:384] <= 32'h0FF0000F;
            reg_val_0_80000000[4][447:416] <= 32'h00100193;
            reg_val_0_80000000[4][479:448] <= 32'h05D00893;
            reg_val_0_80000000[4][511:480] <= 32'h00000513;
            reg_val_0_80000000[5][31:0] <= 32'h00000073;
            reg_val_0_80000000[5][63:32] <= 32'h00000293;
            reg_val_0_80000000[5][95:64] <= 32'h00028A63;
            reg_val_0_80000000[5][127:96] <= 32'h10529073;
            reg_val_0_80000000[5][159:128] <= 32'h0000B2B7;
            reg_val_0_80000000[5][191:160] <= 32'h10928293;
            reg_val_0_80000000[5][223:192] <= 32'h30229073;
            reg_val_0_80000000[5][255:224] <= 32'h30005073;
            reg_val_0_80000000[5][287:256] <= 32'h00002537;
            reg_val_0_80000000[5][319:288] <= 32'h30052073;
            reg_val_0_80000000[5][351:320] <= 32'h00305073;
            reg_val_0_80000000[5][383:352] <= 32'h00000297;
            reg_val_0_80000000[5][415:384] <= 32'h01428293;
            reg_val_0_80000000[5][447:416] <= 32'h34129073;
            reg_val_0_80000000[5][479:448] <= 32'hF1402573;
            reg_val_0_80000000[5][511:480] <= 32'h30200073;
            reg_val_0_80000000[6][31:0] <= 32'h00200193;
            reg_val_0_80000000[6][63:32] <= 32'h00002517;
            reg_val_0_80000000[6][95:64] <= 32'hE7C50513;
            reg_val_0_80000000[6][127:96] <= 32'h00053007;
            reg_val_0_80000000[6][159:128] <= 32'h00853087;
            reg_val_0_80000000[6][191:160] <= 32'h01053107;
            reg_val_0_80000000[6][223:192] <= 32'h01852683;
            reg_val_0_80000000[6][255:224] <= 32'h01C52303;
            reg_val_0_80000000[6][287:256] <= 32'h021071D3;
            reg_val_0_80000000[6][319:288] <= 32'h00353027;
            reg_val_0_80000000[6][351:320] <= 32'h00452383;
            reg_val_0_80000000[6][383:352] <= 32'h00052503;
            reg_val_0_80000000[6][415:384] <= 32'h001015F3;
            reg_val_0_80000000[6][447:416] <= 32'h00000613;
            reg_val_0_80000000[6][479:448] <= 32'h26D51A63;
            reg_val_0_80000000[6][511:480] <= 32'h26731863;
            reg_val_0_80000000[7][31:0] <= 32'h26C59663;
            reg_val_0_80000000[7][63:32] <= 32'h00300193;
            reg_val_0_80000000[7][95:64] <= 32'h00002517;
            reg_val_0_80000000[7][127:96] <= 32'hE5850513;
            reg_val_0_80000000[7][159:128] <= 32'h00053007;
            reg_val_0_80000000[7][191:160] <= 32'h00853087;
            reg_val_0_80000000[7][223:192] <= 32'h01053107;
            reg_val_0_80000000[7][255:224] <= 32'h01852683;
            reg_val_0_80000000[7][287:256] <= 32'h01C52303;
            reg_val_0_80000000[7][319:288] <= 32'h021071D3;
            reg_val_0_80000000[7][351:320] <= 32'h00353027;
            reg_val_0_80000000[7][383:352] <= 32'h00452383;
            reg_val_0_80000000[7][415:384] <= 32'h00052503;
            reg_val_0_80000000[7][447:416] <= 32'h001015F3;
            reg_val_0_80000000[7][479:448] <= 32'h00100613;
            reg_val_0_80000000[7][511:480] <= 32'h22D51863;
            reg_val_0_80000000[8][31:0] <= 32'h22731663;
            reg_val_0_80000000[8][63:32] <= 32'h22C59463;
            reg_val_0_80000000[8][95:64] <= 32'h00400193;
            reg_val_0_80000000[8][127:96] <= 32'h00002517;
            reg_val_0_80000000[8][159:128] <= 32'hE3450513;
            reg_val_0_80000000[8][191:160] <= 32'h00053007;
            reg_val_0_80000000[8][223:192] <= 32'h00853087;
            reg_val_0_80000000[8][255:224] <= 32'h01053107;
            reg_val_0_80000000[8][287:256] <= 32'h01852683;
            reg_val_0_80000000[8][319:288] <= 32'h01C52303;
            reg_val_0_80000000[8][351:320] <= 32'h021071D3;
            reg_val_0_80000000[8][383:352] <= 32'h00353027;
            reg_val_0_80000000[8][415:384] <= 32'h00452383;
            reg_val_0_80000000[8][447:416] <= 32'h00052503;
            reg_val_0_80000000[8][479:448] <= 32'h001015F3;
            reg_val_0_80000000[8][511:480] <= 32'h00100613;
            reg_val_0_80000000[9][31:0] <= 32'h1ED51663;
            reg_val_0_80000000[9][63:32] <= 32'h1E731463;
            reg_val_0_80000000[9][95:64] <= 32'h1EC59263;
            reg_val_0_80000000[9][127:96] <= 32'h00500193;
            reg_val_0_80000000[9][159:128] <= 32'h00002517;
            reg_val_0_80000000[9][191:160] <= 32'hE1050513;
            reg_val_0_80000000[9][223:192] <= 32'h00053007;
            reg_val_0_80000000[9][255:224] <= 32'h00853087;
            reg_val_0_80000000[9][287:256] <= 32'h01053107;
            reg_val_0_80000000[9][319:288] <= 32'h01852683;
            reg_val_0_80000000[9][351:320] <= 32'h01C52303;
            reg_val_0_80000000[9][383:352] <= 32'h0A1071D3;
            reg_val_0_80000000[9][415:384] <= 32'h00353027;
            reg_val_0_80000000[9][447:416] <= 32'h00452383;
            reg_val_0_80000000[9][479:448] <= 32'h00052503;
            reg_val_0_80000000[9][511:480] <= 32'h001015F3;
            reg_val_0_80000000[10][31:0] <= 32'h00000613;
            reg_val_0_80000000[10][63:32] <= 32'h1AD51463;
            reg_val_0_80000000[10][95:64] <= 32'h1A731263;
            reg_val_0_80000000[10][127:96] <= 32'h1AC59063;
            reg_val_0_80000000[10][159:128] <= 32'h00600193;
            reg_val_0_80000000[10][191:160] <= 32'h00002517;
            reg_val_0_80000000[10][223:192] <= 32'hDEC50513;
            reg_val_0_80000000[10][255:224] <= 32'h00053007;
            reg_val_0_80000000[10][287:256] <= 32'h00853087;
            reg_val_0_80000000[10][319:288] <= 32'h01053107;
            reg_val_0_80000000[10][351:320] <= 32'h01852683;
            reg_val_0_80000000[10][383:352] <= 32'h01C52303;
            reg_val_0_80000000[10][415:384] <= 32'h0A1071D3;
            reg_val_0_80000000[10][447:416] <= 32'h00353027;
            reg_val_0_80000000[10][479:448] <= 32'h00452383;
            reg_val_0_80000000[10][511:480] <= 32'h00052503;
            reg_val_0_80000000[11][31:0] <= 32'h001015F3;
            reg_val_0_80000000[11][63:32] <= 32'h00100613;
            reg_val_0_80000000[11][95:64] <= 32'h16D51263;
            reg_val_0_80000000[11][127:96] <= 32'h16731063;
            reg_val_0_80000000[11][159:128] <= 32'h14C59E63;
            reg_val_0_80000000[11][191:160] <= 32'h00700193;
            reg_val_0_80000000[11][223:192] <= 32'h00002517;
            reg_val_0_80000000[11][255:224] <= 32'hDC850513;
            reg_val_0_80000000[11][287:256] <= 32'h00053007;
            reg_val_0_80000000[11][319:288] <= 32'h00853087;
            reg_val_0_80000000[11][351:320] <= 32'h01053107;
            reg_val_0_80000000[11][383:352] <= 32'h01852683;
            reg_val_0_80000000[11][415:384] <= 32'h01C52303;
            reg_val_0_80000000[11][447:416] <= 32'h0A1071D3;
            reg_val_0_80000000[11][479:448] <= 32'h00353027;
            reg_val_0_80000000[11][511:480] <= 32'h00452383;
            reg_val_0_80000000[12][31:0] <= 32'h00052503;
            reg_val_0_80000000[12][63:32] <= 32'h001015F3;
            reg_val_0_80000000[12][95:64] <= 32'h00100613;
            reg_val_0_80000000[12][127:96] <= 32'h12D51063;
            reg_val_0_80000000[12][159:128] <= 32'h10731E63;
            reg_val_0_80000000[12][191:160] <= 32'h10C59C63;
            reg_val_0_80000000[12][223:192] <= 32'h00800193;
            reg_val_0_80000000[12][255:224] <= 32'h00002517;
            reg_val_0_80000000[12][287:256] <= 32'hDA450513;
            reg_val_0_80000000[12][319:288] <= 32'h00053007;
            reg_val_0_80000000[12][351:320] <= 32'h00853087;
            reg_val_0_80000000[12][383:352] <= 32'h01053107;
            reg_val_0_80000000[12][415:384] <= 32'h01852683;
            reg_val_0_80000000[12][447:416] <= 32'h01C52303;
            reg_val_0_80000000[12][479:448] <= 32'h121071D3;
            reg_val_0_80000000[12][511:480] <= 32'h00353027;
            reg_val_0_80000000[13][31:0] <= 32'h00452383;
            reg_val_0_80000000[13][63:32] <= 32'h00052503;
            reg_val_0_80000000[13][95:64] <= 32'h001015F3;
            reg_val_0_80000000[13][127:96] <= 32'h00000613;
            reg_val_0_80000000[13][159:128] <= 32'h0CD51E63;
            reg_val_0_80000000[13][191:160] <= 32'h0C731C63;
            reg_val_0_80000000[13][223:192] <= 32'h0CC59A63;
            reg_val_0_80000000[13][255:224] <= 32'h00900193;
            reg_val_0_80000000[13][287:256] <= 32'h00002517;
            reg_val_0_80000000[13][319:288] <= 32'hD8050513;
            reg_val_0_80000000[13][351:320] <= 32'h00053007;
            reg_val_0_80000000[13][383:352] <= 32'h00853087;
            reg_val_0_80000000[13][415:384] <= 32'h01053107;
            reg_val_0_80000000[13][447:416] <= 32'h01852683;
            reg_val_0_80000000[13][479:448] <= 32'h01C52303;
            reg_val_0_80000000[13][511:480] <= 32'h121071D3;
            reg_val_0_80000000[14][31:0] <= 32'h00353027;
            reg_val_0_80000000[14][63:32] <= 32'h00452383;
            reg_val_0_80000000[14][95:64] <= 32'h00052503;
            reg_val_0_80000000[14][127:96] <= 32'h001015F3;
            reg_val_0_80000000[14][159:128] <= 32'h00100613;
            reg_val_0_80000000[14][191:160] <= 32'h08D51C63;
            reg_val_0_80000000[14][223:192] <= 32'h08731A63;
            reg_val_0_80000000[14][255:224] <= 32'h08C59863;
            reg_val_0_80000000[14][287:256] <= 32'h00A00193;
            reg_val_0_80000000[14][319:288] <= 32'h00002517;
            reg_val_0_80000000[14][351:320] <= 32'hD5C50513;
            reg_val_0_80000000[14][383:352] <= 32'h00053007;
            reg_val_0_80000000[14][415:384] <= 32'h00853087;
            reg_val_0_80000000[14][447:416] <= 32'h01053107;
            reg_val_0_80000000[14][479:448] <= 32'h01852683;
            reg_val_0_80000000[14][511:480] <= 32'h01C52303;
            reg_val_0_80000000[15][31:0] <= 32'h121071D3;
            reg_val_0_80000000[15][63:32] <= 32'h00353027;
            reg_val_0_80000000[15][95:64] <= 32'h00452383;
            reg_val_0_80000000[15][127:96] <= 32'h00052503;
            reg_val_0_80000000[15][159:128] <= 32'h001015F3;
            reg_val_0_80000000[15][191:160] <= 32'h00100613;
            reg_val_0_80000000[15][223:192] <= 32'h04D51A63;
            reg_val_0_80000000[15][255:224] <= 32'h04731863;
            reg_val_0_80000000[15][287:256] <= 32'h04C59663;
            reg_val_0_80000000[15][319:288] <= 32'h00B00193;
            reg_val_0_80000000[15][351:320] <= 32'h00002517;
            reg_val_0_80000000[15][383:352] <= 32'hD3850513;
            reg_val_0_80000000[15][415:384] <= 32'h00053007;
            reg_val_0_80000000[15][447:416] <= 32'h00853087;
            reg_val_0_80000000[15][479:448] <= 32'h01053107;
            reg_val_0_80000000[15][511:480] <= 32'h01852683;
            reg_val_0_80000000[16][31:0] <= 32'h01C52303;
            reg_val_0_80000000[16][63:32] <= 32'h0A1071D3;
            reg_val_0_80000000[16][95:64] <= 32'h00353027;
            reg_val_0_80000000[16][127:96] <= 32'h00452383;
            reg_val_0_80000000[16][159:128] <= 32'h00052503;
            reg_val_0_80000000[16][191:160] <= 32'h001015F3;
            reg_val_0_80000000[16][223:192] <= 32'h01000613;
            reg_val_0_80000000[16][255:224] <= 32'h00D51863;
            reg_val_0_80000000[16][287:256] <= 32'h00731663;
            reg_val_0_80000000[16][319:288] <= 32'h00C59463;
            reg_val_0_80000000[16][351:320] <= 32'h02301063;
            reg_val_0_80000000[16][383:352] <= 32'h0FF0000F;
            reg_val_0_80000000[16][415:384] <= 32'h00018063;
            reg_val_0_80000000[16][447:416] <= 32'h00119193;
            reg_val_0_80000000[16][479:448] <= 32'h0011E193;
            reg_val_0_80000000[16][511:480] <= 32'h05D00893;
            reg_val_0_80000000[17][31:0] <= 32'h00018513;
            reg_val_0_80000000[17][63:32] <= 32'h00000073;
            reg_val_0_80000000[17][95:64] <= 32'h0FF0000F;
            reg_val_0_80000000[17][127:96] <= 32'h00100193;
            reg_val_0_80000000[17][159:128] <= 32'h05D00893;
            reg_val_0_80000000[17][191:160] <= 32'h00000513;
            reg_val_0_80000000[17][223:192] <= 32'h00000073;
            reg_val_0_80000000[17][255:224] <= 32'hC0001073;
            reg_val_0_80000000[17][287:256] <= 32'h00000000;
            reg_val_0_80000000[17][319:288] <= 32'h00000000;
            reg_val_0_80000000[17][351:320] <= 32'h00000000;
            reg_val_0_80000000[17][383:352] <= 32'h00000000;
            reg_val_0_80000000[17][415:384] <= 32'h00000000;
            reg_val_0_80000000[17][447:416] <= 32'h00000000;
            reg_val_0_80000000[17][479:448] <= 32'h00000000;
            // fill-in reset values:
            reg_val_0_80000000[17][511:480] <= 32'h00000000;
            reg_val_0_80000000[18][31:0] <= 32'h00000000;
            reg_val_0_80000000[18][63:32] <= 32'h00000000;
            reg_val_0_80000000[18][95:64] <= 32'h00000000;
            reg_val_0_80000000[18][127:96] <= 32'h00000000;
            reg_val_0_80000000[18][159:128] <= 32'h00000000;
            reg_val_0_80000000[18][191:160] <= 32'h00000000;
            reg_val_0_80000000[18][223:192] <= 32'h00000000;
            reg_val_0_80000000[18][255:224] <= 32'h00000000;
            reg_val_0_80000000[18][287:256] <= 32'h00000000;
            reg_val_0_80000000[18][319:288] <= 32'h00000000;
            reg_val_0_80000000[18][351:320] <= 32'h00000000;
            reg_val_0_80000000[18][383:352] <= 32'h00000000;
            reg_val_0_80000000[18][415:384] <= 32'h00000000;
            reg_val_0_80000000[18][447:416] <= 32'h00000000;
            reg_val_0_80000000[18][479:448] <= 32'h00000000;
            reg_val_0_80000000[18][511:480] <= 32'h00000000;
            reg_val_0_80000000[19][31:0] <= 32'h00000000;
            reg_val_0_80000000[19][63:32] <= 32'h00000000;
            reg_val_0_80000000[19][95:64] <= 32'h00000000;
            reg_val_0_80000000[19][127:96] <= 32'h00000000;
            reg_val_0_80000000[19][159:128] <= 32'h00000000;
            reg_val_0_80000000[19][191:160] <= 32'h00000000;
            reg_val_0_80000000[19][223:192] <= 32'h00000000;
            reg_val_0_80000000[19][255:224] <= 32'h00000000;
            reg_val_0_80000000[19][287:256] <= 32'h00000000;
            reg_val_0_80000000[19][319:288] <= 32'h00000000;
            reg_val_0_80000000[19][351:320] <= 32'h00000000;
            reg_val_0_80000000[19][383:352] <= 32'h00000000;
            reg_val_0_80000000[19][415:384] <= 32'h00000000;
            reg_val_0_80000000[19][447:416] <= 32'h00000000;
            reg_val_0_80000000[19][479:448] <= 32'h00000000;
            reg_val_0_80000000[19][511:480] <= 32'h00000000;
            reg_val_0_80000000[20][31:0] <= 32'h00000000;
            reg_val_0_80000000[20][63:32] <= 32'h00000000;
            reg_val_0_80000000[20][95:64] <= 32'h00000000;
            reg_val_0_80000000[20][127:96] <= 32'h00000000;
            reg_val_0_80000000[20][159:128] <= 32'h00000000;
            reg_val_0_80000000[20][191:160] <= 32'h00000000;
            reg_val_0_80000000[20][223:192] <= 32'h00000000;
            reg_val_0_80000000[20][255:224] <= 32'h00000000;
            reg_val_0_80000000[20][287:256] <= 32'h00000000;
            reg_val_0_80000000[20][319:288] <= 32'h00000000;
            reg_val_0_80000000[20][351:320] <= 32'h00000000;
            reg_val_0_80000000[20][383:352] <= 32'h00000000;
            reg_val_0_80000000[20][415:384] <= 32'h00000000;
            reg_val_0_80000000[20][447:416] <= 32'h00000000;
            reg_val_0_80000000[20][479:448] <= 32'h00000000;
            reg_val_0_80000000[20][511:480] <= 32'h00000000;
            reg_val_0_80000000[21][31:0] <= 32'h00000000;
            reg_val_0_80000000[21][63:32] <= 32'h00000000;
            reg_val_0_80000000[21][95:64] <= 32'h00000000;
            reg_val_0_80000000[21][127:96] <= 32'h00000000;
            reg_val_0_80000000[21][159:128] <= 32'h00000000;
            reg_val_0_80000000[21][191:160] <= 32'h00000000;
            reg_val_0_80000000[21][223:192] <= 32'h00000000;
            reg_val_0_80000000[21][255:224] <= 32'h00000000;
            reg_val_0_80000000[21][287:256] <= 32'h00000000;
            reg_val_0_80000000[21][319:288] <= 32'h00000000;
            reg_val_0_80000000[21][351:320] <= 32'h00000000;
            reg_val_0_80000000[21][383:352] <= 32'h00000000;
            reg_val_0_80000000[21][415:384] <= 32'h00000000;
            reg_val_0_80000000[21][447:416] <= 32'h00000000;
            reg_val_0_80000000[21][479:448] <= 32'h00000000;
            reg_val_0_80000000[21][511:480] <= 32'h00000000;
            reg_val_0_80000000[22][31:0] <= 32'h00000000;
            reg_val_0_80000000[22][63:32] <= 32'h00000000;
            reg_val_0_80000000[22][95:64] <= 32'h00000000;
            reg_val_0_80000000[22][127:96] <= 32'h00000000;
            reg_val_0_80000000[22][159:128] <= 32'h00000000;
            reg_val_0_80000000[22][191:160] <= 32'h00000000;
            reg_val_0_80000000[22][223:192] <= 32'h00000000;
            reg_val_0_80000000[22][255:224] <= 32'h00000000;
            reg_val_0_80000000[22][287:256] <= 32'h00000000;
            reg_val_0_80000000[22][319:288] <= 32'h00000000;
            reg_val_0_80000000[22][351:320] <= 32'h00000000;
            reg_val_0_80000000[22][383:352] <= 32'h00000000;
            reg_val_0_80000000[22][415:384] <= 32'h00000000;
            reg_val_0_80000000[22][447:416] <= 32'h00000000;
            reg_val_0_80000000[22][479:448] <= 32'h00000000;
            reg_val_0_80000000[22][511:480] <= 32'h00000000;
            reg_val_0_80000000[23][31:0] <= 32'h00000000;
            reg_val_0_80000000[23][63:32] <= 32'h00000000;
            reg_val_0_80000000[23][95:64] <= 32'h00000000;
            reg_val_0_80000000[23][127:96] <= 32'h00000000;
            reg_val_0_80000000[23][159:128] <= 32'h00000000;
            reg_val_0_80000000[23][191:160] <= 32'h00000000;
            reg_val_0_80000000[23][223:192] <= 32'h00000000;
            reg_val_0_80000000[23][255:224] <= 32'h00000000;
            reg_val_0_80000000[23][287:256] <= 32'h00000000;
            reg_val_0_80000000[23][319:288] <= 32'h00000000;
            reg_val_0_80000000[23][351:320] <= 32'h00000000;
            reg_val_0_80000000[23][383:352] <= 32'h00000000;
            reg_val_0_80000000[23][415:384] <= 32'h00000000;
            reg_val_0_80000000[23][447:416] <= 32'h00000000;
            reg_val_0_80000000[23][479:448] <= 32'h00000000;
            reg_val_0_80000000[23][511:480] <= 32'h00000000;
            reg_val_0_80000000[24][31:0] <= 32'h00000000;
            reg_val_0_80000000[24][63:32] <= 32'h00000000;
            reg_val_0_80000000[24][95:64] <= 32'h00000000;
            reg_val_0_80000000[24][127:96] <= 32'h00000000;
            reg_val_0_80000000[24][159:128] <= 32'h00000000;
            reg_val_0_80000000[24][191:160] <= 32'h00000000;
            reg_val_0_80000000[24][223:192] <= 32'h00000000;
            reg_val_0_80000000[24][255:224] <= 32'h00000000;
            reg_val_0_80000000[24][287:256] <= 32'h00000000;
            reg_val_0_80000000[24][319:288] <= 32'h00000000;
            reg_val_0_80000000[24][351:320] <= 32'h00000000;
            reg_val_0_80000000[24][383:352] <= 32'h00000000;
            reg_val_0_80000000[24][415:384] <= 32'h00000000;
            reg_val_0_80000000[24][447:416] <= 32'h00000000;
            reg_val_0_80000000[24][479:448] <= 32'h00000000;
            reg_val_0_80000000[24][511:480] <= 32'h00000000;
            reg_val_0_80000000[25][31:0] <= 32'h00000000;
            reg_val_0_80000000[25][63:32] <= 32'h00000000;
            reg_val_0_80000000[25][95:64] <= 32'h00000000;
            reg_val_0_80000000[25][127:96] <= 32'h00000000;
            reg_val_0_80000000[25][159:128] <= 32'h00000000;
            reg_val_0_80000000[25][191:160] <= 32'h00000000;
            reg_val_0_80000000[25][223:192] <= 32'h00000000;
            reg_val_0_80000000[25][255:224] <= 32'h00000000;
            reg_val_0_80000000[25][287:256] <= 32'h00000000;
            reg_val_0_80000000[25][319:288] <= 32'h00000000;
            reg_val_0_80000000[25][351:320] <= 32'h00000000;
            reg_val_0_80000000[25][383:352] <= 32'h00000000;
            reg_val_0_80000000[25][415:384] <= 32'h00000000;
            reg_val_0_80000000[25][447:416] <= 32'h00000000;
            reg_val_0_80000000[25][479:448] <= 32'h00000000;
            reg_val_0_80000000[25][511:480] <= 32'h00000000;
            reg_val_0_80000000[26][31:0] <= 32'h00000000;
            reg_val_0_80000000[26][63:32] <= 32'h00000000;
            reg_val_0_80000000[26][95:64] <= 32'h00000000;
            reg_val_0_80000000[26][127:96] <= 32'h00000000;
            reg_val_0_80000000[26][159:128] <= 32'h00000000;
            reg_val_0_80000000[26][191:160] <= 32'h00000000;
            reg_val_0_80000000[26][223:192] <= 32'h00000000;
            reg_val_0_80000000[26][255:224] <= 32'h00000000;
            reg_val_0_80000000[26][287:256] <= 32'h00000000;
            reg_val_0_80000000[26][319:288] <= 32'h00000000;
            reg_val_0_80000000[26][351:320] <= 32'h00000000;
            reg_val_0_80000000[26][383:352] <= 32'h00000000;
            reg_val_0_80000000[26][415:384] <= 32'h00000000;
            reg_val_0_80000000[26][447:416] <= 32'h00000000;
            reg_val_0_80000000[26][479:448] <= 32'h00000000;
            reg_val_0_80000000[26][511:480] <= 32'h00000000;
            reg_val_0_80000000[27][31:0] <= 32'h00000000;
            reg_val_0_80000000[27][63:32] <= 32'h00000000;
            reg_val_0_80000000[27][95:64] <= 32'h00000000;
            reg_val_0_80000000[27][127:96] <= 32'h00000000;
            reg_val_0_80000000[27][159:128] <= 32'h00000000;
            reg_val_0_80000000[27][191:160] <= 32'h00000000;
            reg_val_0_80000000[27][223:192] <= 32'h00000000;
            reg_val_0_80000000[27][255:224] <= 32'h00000000;
            reg_val_0_80000000[27][287:256] <= 32'h00000000;
            reg_val_0_80000000[27][319:288] <= 32'h00000000;
            reg_val_0_80000000[27][351:320] <= 32'h00000000;
            reg_val_0_80000000[27][383:352] <= 32'h00000000;
            reg_val_0_80000000[27][415:384] <= 32'h00000000;
            reg_val_0_80000000[27][447:416] <= 32'h00000000;
            reg_val_0_80000000[27][479:448] <= 32'h00000000;
            reg_val_0_80000000[27][511:480] <= 32'h00000000;
            reg_val_0_80000000[28][31:0] <= 32'h00000000;
            reg_val_0_80000000[28][63:32] <= 32'h00000000;
            reg_val_0_80000000[28][95:64] <= 32'h00000000;
            reg_val_0_80000000[28][127:96] <= 32'h00000000;
            reg_val_0_80000000[28][159:128] <= 32'h00000000;
            reg_val_0_80000000[28][191:160] <= 32'h00000000;
            reg_val_0_80000000[28][223:192] <= 32'h00000000;
            reg_val_0_80000000[28][255:224] <= 32'h00000000;
            reg_val_0_80000000[28][287:256] <= 32'h00000000;
            reg_val_0_80000000[28][319:288] <= 32'h00000000;
            reg_val_0_80000000[28][351:320] <= 32'h00000000;
            reg_val_0_80000000[28][383:352] <= 32'h00000000;
            reg_val_0_80000000[28][415:384] <= 32'h00000000;
            reg_val_0_80000000[28][447:416] <= 32'h00000000;
            reg_val_0_80000000[28][479:448] <= 32'h00000000;
            reg_val_0_80000000[28][511:480] <= 32'h00000000;
            reg_val_0_80000000[29][31:0] <= 32'h00000000;
            reg_val_0_80000000[29][63:32] <= 32'h00000000;
            reg_val_0_80000000[29][95:64] <= 32'h00000000;
            reg_val_0_80000000[29][127:96] <= 32'h00000000;
            reg_val_0_80000000[29][159:128] <= 32'h00000000;
            reg_val_0_80000000[29][191:160] <= 32'h00000000;
            reg_val_0_80000000[29][223:192] <= 32'h00000000;
            reg_val_0_80000000[29][255:224] <= 32'h00000000;
            reg_val_0_80000000[29][287:256] <= 32'h00000000;
            reg_val_0_80000000[29][319:288] <= 32'h00000000;
            reg_val_0_80000000[29][351:320] <= 32'h00000000;
            reg_val_0_80000000[29][383:352] <= 32'h00000000;
            reg_val_0_80000000[29][415:384] <= 32'h00000000;
            reg_val_0_80000000[29][447:416] <= 32'h00000000;
            reg_val_0_80000000[29][479:448] <= 32'h00000000;
            reg_val_0_80000000[29][511:480] <= 32'h00000000;
            reg_val_0_80000000[30][31:0] <= 32'h00000000;
            reg_val_0_80000000[30][63:32] <= 32'h00000000;
            reg_val_0_80000000[30][95:64] <= 32'h00000000;
            reg_val_0_80000000[30][127:96] <= 32'h00000000;
            reg_val_0_80000000[30][159:128] <= 32'h00000000;
            reg_val_0_80000000[30][191:160] <= 32'h00000000;
            reg_val_0_80000000[30][223:192] <= 32'h00000000;
            reg_val_0_80000000[30][255:224] <= 32'h00000000;
            reg_val_0_80000000[30][287:256] <= 32'h00000000;
            reg_val_0_80000000[30][319:288] <= 32'h00000000;
            reg_val_0_80000000[30][351:320] <= 32'h00000000;
            reg_val_0_80000000[30][383:352] <= 32'h00000000;
            reg_val_0_80000000[30][415:384] <= 32'h00000000;
            reg_val_0_80000000[30][447:416] <= 32'h00000000;
            reg_val_0_80000000[30][479:448] <= 32'h00000000;
            reg_val_0_80000000[30][511:480] <= 32'h00000000;
            reg_val_0_80000000[31][31:0] <= 32'h00000000;
            reg_val_0_80000000[31][63:32] <= 32'h00000000;
            reg_val_0_80000000[31][95:64] <= 32'h00000000;
            reg_val_0_80000000[31][127:96] <= 32'h00000000;
            reg_val_0_80000000[31][159:128] <= 32'h00000000;
            reg_val_0_80000000[31][191:160] <= 32'h00000000;
            reg_val_0_80000000[31][223:192] <= 32'h00000000;
            reg_val_0_80000000[31][255:224] <= 32'h00000000;
            reg_val_0_80000000[31][287:256] <= 32'h00000000;
            reg_val_0_80000000[31][319:288] <= 32'h00000000;
            reg_val_0_80000000[31][351:320] <= 32'h00000000;
            reg_val_0_80000000[31][383:352] <= 32'h00000000;
            reg_val_0_80000000[31][415:384] <= 32'h00000000;
            reg_val_0_80000000[31][447:416] <= 32'h00000000;
            reg_val_0_80000000[31][479:448] <= 32'h00000000;
            reg_val_0_80000000[31][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_0_80000000 <= next_reg_val_0_80000000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_0_80000000
        // hold reg val by default
        for (int i = 0; i < 32; i++)
        begin
            next_reg_val_0_80000000[i] = reg_val_0_80000000[i];
        end
        // update reg val if wen
        if (wen_0_80000000)
        begin
            // check for this byte enabled
            if (mem_req_byteen[0])  next_reg_val_0_80000000[wsel_0_80000000][7:0] = wdata_0_80000000[7:0];
            if (mem_req_byteen[1])  next_reg_val_0_80000000[wsel_0_80000000][15:8] = wdata_0_80000000[15:8];
            if (mem_req_byteen[2])  next_reg_val_0_80000000[wsel_0_80000000][23:16] = wdata_0_80000000[23:16];
            if (mem_req_byteen[3])  next_reg_val_0_80000000[wsel_0_80000000][31:24] = wdata_0_80000000[31:24];
            if (mem_req_byteen[4])  next_reg_val_0_80000000[wsel_0_80000000][39:32] = wdata_0_80000000[39:32];
            if (mem_req_byteen[5])  next_reg_val_0_80000000[wsel_0_80000000][47:40] = wdata_0_80000000[47:40];
            if (mem_req_byteen[6])  next_reg_val_0_80000000[wsel_0_80000000][55:48] = wdata_0_80000000[55:48];
            if (mem_req_byteen[7])  next_reg_val_0_80000000[wsel_0_80000000][63:56] = wdata_0_80000000[63:56];
            if (mem_req_byteen[8])  next_reg_val_0_80000000[wsel_0_80000000][71:64] = wdata_0_80000000[71:64];
            if (mem_req_byteen[9])  next_reg_val_0_80000000[wsel_0_80000000][79:72] = wdata_0_80000000[79:72];
            if (mem_req_byteen[10])  next_reg_val_0_80000000[wsel_0_80000000][87:80] = wdata_0_80000000[87:80];
            if (mem_req_byteen[11])  next_reg_val_0_80000000[wsel_0_80000000][95:88] = wdata_0_80000000[95:88];
            if (mem_req_byteen[12])  next_reg_val_0_80000000[wsel_0_80000000][103:96] = wdata_0_80000000[103:96];
            if (mem_req_byteen[13])  next_reg_val_0_80000000[wsel_0_80000000][111:104] = wdata_0_80000000[111:104];
            if (mem_req_byteen[14])  next_reg_val_0_80000000[wsel_0_80000000][119:112] = wdata_0_80000000[119:112];
            if (mem_req_byteen[15])  next_reg_val_0_80000000[wsel_0_80000000][127:120] = wdata_0_80000000[127:120];
            if (mem_req_byteen[16])  next_reg_val_0_80000000[wsel_0_80000000][135:128] = wdata_0_80000000[135:128];
            if (mem_req_byteen[17])  next_reg_val_0_80000000[wsel_0_80000000][143:136] = wdata_0_80000000[143:136];
            if (mem_req_byteen[18])  next_reg_val_0_80000000[wsel_0_80000000][151:144] = wdata_0_80000000[151:144];
            if (mem_req_byteen[19])  next_reg_val_0_80000000[wsel_0_80000000][159:152] = wdata_0_80000000[159:152];
            if (mem_req_byteen[20])  next_reg_val_0_80000000[wsel_0_80000000][167:160] = wdata_0_80000000[167:160];
            if (mem_req_byteen[21])  next_reg_val_0_80000000[wsel_0_80000000][175:168] = wdata_0_80000000[175:168];
            if (mem_req_byteen[22])  next_reg_val_0_80000000[wsel_0_80000000][183:176] = wdata_0_80000000[183:176];
            if (mem_req_byteen[23])  next_reg_val_0_80000000[wsel_0_80000000][191:184] = wdata_0_80000000[191:184];
            if (mem_req_byteen[24])  next_reg_val_0_80000000[wsel_0_80000000][199:192] = wdata_0_80000000[199:192];
            if (mem_req_byteen[25])  next_reg_val_0_80000000[wsel_0_80000000][207:200] = wdata_0_80000000[207:200];
            if (mem_req_byteen[26])  next_reg_val_0_80000000[wsel_0_80000000][215:208] = wdata_0_80000000[215:208];
            if (mem_req_byteen[27])  next_reg_val_0_80000000[wsel_0_80000000][223:216] = wdata_0_80000000[223:216];
            if (mem_req_byteen[28])  next_reg_val_0_80000000[wsel_0_80000000][231:224] = wdata_0_80000000[231:224];
            if (mem_req_byteen[29])  next_reg_val_0_80000000[wsel_0_80000000][239:232] = wdata_0_80000000[239:232];
            if (mem_req_byteen[30])  next_reg_val_0_80000000[wsel_0_80000000][247:240] = wdata_0_80000000[247:240];
            if (mem_req_byteen[31])  next_reg_val_0_80000000[wsel_0_80000000][255:248] = wdata_0_80000000[255:248];
            if (mem_req_byteen[32])  next_reg_val_0_80000000[wsel_0_80000000][263:256] = wdata_0_80000000[263:256];
            if (mem_req_byteen[33])  next_reg_val_0_80000000[wsel_0_80000000][271:264] = wdata_0_80000000[271:264];
            if (mem_req_byteen[34])  next_reg_val_0_80000000[wsel_0_80000000][279:272] = wdata_0_80000000[279:272];
            if (mem_req_byteen[35])  next_reg_val_0_80000000[wsel_0_80000000][287:280] = wdata_0_80000000[287:280];
            if (mem_req_byteen[36])  next_reg_val_0_80000000[wsel_0_80000000][295:288] = wdata_0_80000000[295:288];
            if (mem_req_byteen[37])  next_reg_val_0_80000000[wsel_0_80000000][303:296] = wdata_0_80000000[303:296];
            if (mem_req_byteen[38])  next_reg_val_0_80000000[wsel_0_80000000][311:304] = wdata_0_80000000[311:304];
            if (mem_req_byteen[39])  next_reg_val_0_80000000[wsel_0_80000000][319:312] = wdata_0_80000000[319:312];
            if (mem_req_byteen[40])  next_reg_val_0_80000000[wsel_0_80000000][327:320] = wdata_0_80000000[327:320];
            if (mem_req_byteen[41])  next_reg_val_0_80000000[wsel_0_80000000][335:328] = wdata_0_80000000[335:328];
            if (mem_req_byteen[42])  next_reg_val_0_80000000[wsel_0_80000000][343:336] = wdata_0_80000000[343:336];
            if (mem_req_byteen[43])  next_reg_val_0_80000000[wsel_0_80000000][351:344] = wdata_0_80000000[351:344];
            if (mem_req_byteen[44])  next_reg_val_0_80000000[wsel_0_80000000][359:352] = wdata_0_80000000[359:352];
            if (mem_req_byteen[45])  next_reg_val_0_80000000[wsel_0_80000000][367:360] = wdata_0_80000000[367:360];
            if (mem_req_byteen[46])  next_reg_val_0_80000000[wsel_0_80000000][375:368] = wdata_0_80000000[375:368];
            if (mem_req_byteen[47])  next_reg_val_0_80000000[wsel_0_80000000][383:376] = wdata_0_80000000[383:376];
            if (mem_req_byteen[48])  next_reg_val_0_80000000[wsel_0_80000000][391:384] = wdata_0_80000000[391:384];
            if (mem_req_byteen[49])  next_reg_val_0_80000000[wsel_0_80000000][399:392] = wdata_0_80000000[399:392];
            if (mem_req_byteen[50])  next_reg_val_0_80000000[wsel_0_80000000][407:400] = wdata_0_80000000[407:400];
            if (mem_req_byteen[51])  next_reg_val_0_80000000[wsel_0_80000000][415:408] = wdata_0_80000000[415:408];
            if (mem_req_byteen[52])  next_reg_val_0_80000000[wsel_0_80000000][423:416] = wdata_0_80000000[423:416];
            if (mem_req_byteen[53])  next_reg_val_0_80000000[wsel_0_80000000][431:424] = wdata_0_80000000[431:424];
            if (mem_req_byteen[54])  next_reg_val_0_80000000[wsel_0_80000000][439:432] = wdata_0_80000000[439:432];
            if (mem_req_byteen[55])  next_reg_val_0_80000000[wsel_0_80000000][447:440] = wdata_0_80000000[447:440];
            if (mem_req_byteen[56])  next_reg_val_0_80000000[wsel_0_80000000][455:448] = wdata_0_80000000[455:448];
            if (mem_req_byteen[57])  next_reg_val_0_80000000[wsel_0_80000000][463:456] = wdata_0_80000000[463:456];
            if (mem_req_byteen[58])  next_reg_val_0_80000000[wsel_0_80000000][471:464] = wdata_0_80000000[471:464];
            if (mem_req_byteen[59])  next_reg_val_0_80000000[wsel_0_80000000][479:472] = wdata_0_80000000[479:472];
            if (mem_req_byteen[60])  next_reg_val_0_80000000[wsel_0_80000000][487:480] = wdata_0_80000000[487:480];
            if (mem_req_byteen[61])  next_reg_val_0_80000000[wsel_0_80000000][495:488] = wdata_0_80000000[495:488];
            if (mem_req_byteen[62])  next_reg_val_0_80000000[wsel_0_80000000][503:496] = wdata_0_80000000[503:496];
            if (mem_req_byteen[63])  next_reg_val_0_80000000[wsel_0_80000000][511:504] = wdata_0_80000000[511:504];
        end
    end
    
    always_comb begin : READ_LOGIC_0_80000000
        // read val at rsel
        // multi block version (need select line)
        rdata_0_80000000 = reg_val_0_80000000[rsel_0_80000000];
    end
    
    // chunk 1
    logic wen_1_80001000;
    
    // block selection within reg file
    logic [1-1:0] wsel_1_80001000;
    logic [1-1:0] rsel_1_80001000;
    
    // lock-sized reg file write input and read output
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_1_80001000;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_1_80001000;
    
    // 2D register file
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_1_80001000 [2-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_1_80001000 [2-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_1_80001000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_1_80001000[0][31:0] <= 32'h00000000;
            reg_val_1_80001000[0][63:32] <= 32'h00000000;
            reg_val_1_80001000[0][95:64] <= 32'h00000000;
            reg_val_1_80001000[0][127:96] <= 32'h00000000;
            reg_val_1_80001000[0][159:128] <= 32'h00000000;
            reg_val_1_80001000[0][191:160] <= 32'h00000000;
            reg_val_1_80001000[0][223:192] <= 32'h00000000;
            reg_val_1_80001000[0][255:224] <= 32'h00000000;
            reg_val_1_80001000[0][287:256] <= 32'h00000000;
            reg_val_1_80001000[0][319:288] <= 32'h00000000;
            reg_val_1_80001000[0][351:320] <= 32'h00000000;
            reg_val_1_80001000[0][383:352] <= 32'h00000000;
            reg_val_1_80001000[0][415:384] <= 32'h00000000;
            reg_val_1_80001000[0][447:416] <= 32'h00000000;
            reg_val_1_80001000[0][479:448] <= 32'h00000000;
            reg_val_1_80001000[0][511:480] <= 32'h00000000;
            reg_val_1_80001000[1][31:0] <= 32'h00000000;
            reg_val_1_80001000[1][63:32] <= 32'h00000000;
            // fill-in reset values:
            reg_val_1_80001000[1][95:64] <= 32'h00000000;
            reg_val_1_80001000[1][127:96] <= 32'h00000000;
            reg_val_1_80001000[1][159:128] <= 32'h00000000;
            reg_val_1_80001000[1][191:160] <= 32'h00000000;
            reg_val_1_80001000[1][223:192] <= 32'h00000000;
            reg_val_1_80001000[1][255:224] <= 32'h00000000;
            reg_val_1_80001000[1][287:256] <= 32'h00000000;
            reg_val_1_80001000[1][319:288] <= 32'h00000000;
            reg_val_1_80001000[1][351:320] <= 32'h00000000;
            reg_val_1_80001000[1][383:352] <= 32'h00000000;
            reg_val_1_80001000[1][415:384] <= 32'h00000000;
            reg_val_1_80001000[1][447:416] <= 32'h00000000;
            reg_val_1_80001000[1][479:448] <= 32'h00000000;
            reg_val_1_80001000[1][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_1_80001000 <= next_reg_val_1_80001000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_1_80001000
        // hold reg val by default
        for (int i = 0; i < 2; i++)
        begin
            next_reg_val_1_80001000[i] = reg_val_1_80001000[i];
        end
        // update reg val if wen
        if (wen_1_80001000)
        begin
            // check for this byte enabled
            if (mem_req_byteen[0])  next_reg_val_1_80001000[wsel_1_80001000][7:0] = wdata_1_80001000[7:0];
            if (mem_req_byteen[1])  next_reg_val_1_80001000[wsel_1_80001000][15:8] = wdata_1_80001000[15:8];
            if (mem_req_byteen[2])  next_reg_val_1_80001000[wsel_1_80001000][23:16] = wdata_1_80001000[23:16];
            if (mem_req_byteen[3])  next_reg_val_1_80001000[wsel_1_80001000][31:24] = wdata_1_80001000[31:24];
            if (mem_req_byteen[4])  next_reg_val_1_80001000[wsel_1_80001000][39:32] = wdata_1_80001000[39:32];
            if (mem_req_byteen[5])  next_reg_val_1_80001000[wsel_1_80001000][47:40] = wdata_1_80001000[47:40];
            if (mem_req_byteen[6])  next_reg_val_1_80001000[wsel_1_80001000][55:48] = wdata_1_80001000[55:48];
            if (mem_req_byteen[7])  next_reg_val_1_80001000[wsel_1_80001000][63:56] = wdata_1_80001000[63:56];
            if (mem_req_byteen[8])  next_reg_val_1_80001000[wsel_1_80001000][71:64] = wdata_1_80001000[71:64];
            if (mem_req_byteen[9])  next_reg_val_1_80001000[wsel_1_80001000][79:72] = wdata_1_80001000[79:72];
            if (mem_req_byteen[10])  next_reg_val_1_80001000[wsel_1_80001000][87:80] = wdata_1_80001000[87:80];
            if (mem_req_byteen[11])  next_reg_val_1_80001000[wsel_1_80001000][95:88] = wdata_1_80001000[95:88];
            if (mem_req_byteen[12])  next_reg_val_1_80001000[wsel_1_80001000][103:96] = wdata_1_80001000[103:96];
            if (mem_req_byteen[13])  next_reg_val_1_80001000[wsel_1_80001000][111:104] = wdata_1_80001000[111:104];
            if (mem_req_byteen[14])  next_reg_val_1_80001000[wsel_1_80001000][119:112] = wdata_1_80001000[119:112];
            if (mem_req_byteen[15])  next_reg_val_1_80001000[wsel_1_80001000][127:120] = wdata_1_80001000[127:120];
            if (mem_req_byteen[16])  next_reg_val_1_80001000[wsel_1_80001000][135:128] = wdata_1_80001000[135:128];
            if (mem_req_byteen[17])  next_reg_val_1_80001000[wsel_1_80001000][143:136] = wdata_1_80001000[143:136];
            if (mem_req_byteen[18])  next_reg_val_1_80001000[wsel_1_80001000][151:144] = wdata_1_80001000[151:144];
            if (mem_req_byteen[19])  next_reg_val_1_80001000[wsel_1_80001000][159:152] = wdata_1_80001000[159:152];
            if (mem_req_byteen[20])  next_reg_val_1_80001000[wsel_1_80001000][167:160] = wdata_1_80001000[167:160];
            if (mem_req_byteen[21])  next_reg_val_1_80001000[wsel_1_80001000][175:168] = wdata_1_80001000[175:168];
            if (mem_req_byteen[22])  next_reg_val_1_80001000[wsel_1_80001000][183:176] = wdata_1_80001000[183:176];
            if (mem_req_byteen[23])  next_reg_val_1_80001000[wsel_1_80001000][191:184] = wdata_1_80001000[191:184];
            if (mem_req_byteen[24])  next_reg_val_1_80001000[wsel_1_80001000][199:192] = wdata_1_80001000[199:192];
            if (mem_req_byteen[25])  next_reg_val_1_80001000[wsel_1_80001000][207:200] = wdata_1_80001000[207:200];
            if (mem_req_byteen[26])  next_reg_val_1_80001000[wsel_1_80001000][215:208] = wdata_1_80001000[215:208];
            if (mem_req_byteen[27])  next_reg_val_1_80001000[wsel_1_80001000][223:216] = wdata_1_80001000[223:216];
            if (mem_req_byteen[28])  next_reg_val_1_80001000[wsel_1_80001000][231:224] = wdata_1_80001000[231:224];
            if (mem_req_byteen[29])  next_reg_val_1_80001000[wsel_1_80001000][239:232] = wdata_1_80001000[239:232];
            if (mem_req_byteen[30])  next_reg_val_1_80001000[wsel_1_80001000][247:240] = wdata_1_80001000[247:240];
            if (mem_req_byteen[31])  next_reg_val_1_80001000[wsel_1_80001000][255:248] = wdata_1_80001000[255:248];
            if (mem_req_byteen[32])  next_reg_val_1_80001000[wsel_1_80001000][263:256] = wdata_1_80001000[263:256];
            if (mem_req_byteen[33])  next_reg_val_1_80001000[wsel_1_80001000][271:264] = wdata_1_80001000[271:264];
            if (mem_req_byteen[34])  next_reg_val_1_80001000[wsel_1_80001000][279:272] = wdata_1_80001000[279:272];
            if (mem_req_byteen[35])  next_reg_val_1_80001000[wsel_1_80001000][287:280] = wdata_1_80001000[287:280];
            if (mem_req_byteen[36])  next_reg_val_1_80001000[wsel_1_80001000][295:288] = wdata_1_80001000[295:288];
            if (mem_req_byteen[37])  next_reg_val_1_80001000[wsel_1_80001000][303:296] = wdata_1_80001000[303:296];
            if (mem_req_byteen[38])  next_reg_val_1_80001000[wsel_1_80001000][311:304] = wdata_1_80001000[311:304];
            if (mem_req_byteen[39])  next_reg_val_1_80001000[wsel_1_80001000][319:312] = wdata_1_80001000[319:312];
            if (mem_req_byteen[40])  next_reg_val_1_80001000[wsel_1_80001000][327:320] = wdata_1_80001000[327:320];
            if (mem_req_byteen[41])  next_reg_val_1_80001000[wsel_1_80001000][335:328] = wdata_1_80001000[335:328];
            if (mem_req_byteen[42])  next_reg_val_1_80001000[wsel_1_80001000][343:336] = wdata_1_80001000[343:336];
            if (mem_req_byteen[43])  next_reg_val_1_80001000[wsel_1_80001000][351:344] = wdata_1_80001000[351:344];
            if (mem_req_byteen[44])  next_reg_val_1_80001000[wsel_1_80001000][359:352] = wdata_1_80001000[359:352];
            if (mem_req_byteen[45])  next_reg_val_1_80001000[wsel_1_80001000][367:360] = wdata_1_80001000[367:360];
            if (mem_req_byteen[46])  next_reg_val_1_80001000[wsel_1_80001000][375:368] = wdata_1_80001000[375:368];
            if (mem_req_byteen[47])  next_reg_val_1_80001000[wsel_1_80001000][383:376] = wdata_1_80001000[383:376];
            if (mem_req_byteen[48])  next_reg_val_1_80001000[wsel_1_80001000][391:384] = wdata_1_80001000[391:384];
            if (mem_req_byteen[49])  next_reg_val_1_80001000[wsel_1_80001000][399:392] = wdata_1_80001000[399:392];
            if (mem_req_byteen[50])  next_reg_val_1_80001000[wsel_1_80001000][407:400] = wdata_1_80001000[407:400];
            if (mem_req_byteen[51])  next_reg_val_1_80001000[wsel_1_80001000][415:408] = wdata_1_80001000[415:408];
            if (mem_req_byteen[52])  next_reg_val_1_80001000[wsel_1_80001000][423:416] = wdata_1_80001000[423:416];
            if (mem_req_byteen[53])  next_reg_val_1_80001000[wsel_1_80001000][431:424] = wdata_1_80001000[431:424];
            if (mem_req_byteen[54])  next_reg_val_1_80001000[wsel_1_80001000][439:432] = wdata_1_80001000[439:432];
            if (mem_req_byteen[55])  next_reg_val_1_80001000[wsel_1_80001000][447:440] = wdata_1_80001000[447:440];
            if (mem_req_byteen[56])  next_reg_val_1_80001000[wsel_1_80001000][455:448] = wdata_1_80001000[455:448];
            if (mem_req_byteen[57])  next_reg_val_1_80001000[wsel_1_80001000][463:456] = wdata_1_80001000[463:456];
            if (mem_req_byteen[58])  next_reg_val_1_80001000[wsel_1_80001000][471:464] = wdata_1_80001000[471:464];
            if (mem_req_byteen[59])  next_reg_val_1_80001000[wsel_1_80001000][479:472] = wdata_1_80001000[479:472];
            if (mem_req_byteen[60])  next_reg_val_1_80001000[wsel_1_80001000][487:480] = wdata_1_80001000[487:480];
            if (mem_req_byteen[61])  next_reg_val_1_80001000[wsel_1_80001000][495:488] = wdata_1_80001000[495:488];
            if (mem_req_byteen[62])  next_reg_val_1_80001000[wsel_1_80001000][503:496] = wdata_1_80001000[503:496];
            if (mem_req_byteen[63])  next_reg_val_1_80001000[wsel_1_80001000][511:504] = wdata_1_80001000[511:504];
        end
    end
    
    always_comb begin : READ_LOGIC_1_80001000
        // read val at rsel
        // multi block version (need select line)
        rdata_1_80001000 = reg_val_1_80001000[rsel_1_80001000];
    end
    
    // chunk 2
    logic wen_2_80002000;
    
    // block selection within reg file
    logic [3-1:0] wsel_2_80002000;
    logic [3-1:0] rsel_2_80002000;
    
    // lock-sized reg file write input and read output
    logic [`VX_MEM_DATA_WIDTH-1:0] wdata_2_80002000;
    logic [`VX_MEM_DATA_WIDTH-1:0] rdata_2_80002000;
    
    // 2D register file
    logic [`VX_MEM_DATA_WIDTH-1:0] reg_val_2_80002000 [8-1:0];
    logic [`VX_MEM_DATA_WIDTH-1:0] next_reg_val_2_80002000 [8-1:0];
    
    always_ff @ (posedge clk) begin : REGISTER_LOGIC_2_80002000
        if (reset)
        begin
            // enumerated reset values:
            reg_val_2_80002000[0][31:0] <= 32'h00000000;
            reg_val_2_80002000[0][63:32] <= 32'h40040000;
            reg_val_2_80002000[0][95:64] <= 32'h00000000;
            reg_val_2_80002000[0][127:96] <= 32'h3FF00000;
            reg_val_2_80002000[0][159:128] <= 32'h00000000;
            reg_val_2_80002000[0][191:160] <= 32'h00000000;
            reg_val_2_80002000[0][223:192] <= 32'h00000000;
            reg_val_2_80002000[0][255:224] <= 32'h400C0000;
            reg_val_2_80002000[0][287:256] <= 32'h66666666;
            reg_val_2_80002000[0][319:288] <= 32'hC0934C66;
            reg_val_2_80002000[0][351:320] <= 32'h9999999A;
            reg_val_2_80002000[0][383:352] <= 32'h3FF19999;
            reg_val_2_80002000[0][415:384] <= 32'h00000000;
            reg_val_2_80002000[0][447:416] <= 32'h00000000;
            reg_val_2_80002000[0][479:448] <= 32'h00000000;
            reg_val_2_80002000[0][511:480] <= 32'hC0934800;
            reg_val_2_80002000[1][31:0] <= 32'h53C8D4F1;
            reg_val_2_80002000[1][63:32] <= 32'h400921FB;
            reg_val_2_80002000[1][95:64] <= 32'hE2308C3A;
            reg_val_2_80002000[1][127:96] <= 32'h3E45798E;
            reg_val_2_80002000[1][159:128] <= 32'h00000000;
            reg_val_2_80002000[1][191:160] <= 32'h00000000;
            reg_val_2_80002000[1][223:192] <= 32'h55206DDF;
            reg_val_2_80002000[1][255:224] <= 32'h400921FB;
            reg_val_2_80002000[1][287:256] <= 32'h00000000;
            reg_val_2_80002000[1][319:288] <= 32'h40040000;
            reg_val_2_80002000[1][351:320] <= 32'h00000000;
            reg_val_2_80002000[1][383:352] <= 32'h3FF00000;
            reg_val_2_80002000[1][415:384] <= 32'h00000000;
            reg_val_2_80002000[1][447:416] <= 32'h00000000;
            reg_val_2_80002000[1][479:448] <= 32'h00000000;
            reg_val_2_80002000[1][511:480] <= 32'h3FF80000;
            reg_val_2_80002000[2][31:0] <= 32'h66666666;
            reg_val_2_80002000[2][63:32] <= 32'hC0934C66;
            reg_val_2_80002000[2][95:64] <= 32'h9999999A;
            reg_val_2_80002000[2][127:96] <= 32'hBFF19999;
            reg_val_2_80002000[2][159:128] <= 32'h00000000;
            reg_val_2_80002000[2][191:160] <= 32'h00000000;
            reg_val_2_80002000[2][223:192] <= 32'h00000000;
            reg_val_2_80002000[2][255:224] <= 32'hC0934800;
            reg_val_2_80002000[2][287:256] <= 32'h53C8D4F1;
            reg_val_2_80002000[2][319:288] <= 32'h400921FB;
            reg_val_2_80002000[2][351:320] <= 32'hE2308C3A;
            reg_val_2_80002000[2][383:352] <= 32'h3E45798E;
            reg_val_2_80002000[2][415:384] <= 32'h00000000;
            reg_val_2_80002000[2][447:416] <= 32'h00000000;
            reg_val_2_80002000[2][479:448] <= 32'h52713C03;
            reg_val_2_80002000[2][511:480] <= 32'h400921FB;
            reg_val_2_80002000[3][31:0] <= 32'h00000000;
            reg_val_2_80002000[3][63:32] <= 32'h40040000;
            reg_val_2_80002000[3][95:64] <= 32'h00000000;
            reg_val_2_80002000[3][127:96] <= 32'h3FF00000;
            reg_val_2_80002000[3][159:128] <= 32'h00000000;
            reg_val_2_80002000[3][191:160] <= 32'h00000000;
            reg_val_2_80002000[3][223:192] <= 32'h00000000;
            reg_val_2_80002000[3][255:224] <= 32'h40040000;
            reg_val_2_80002000[3][287:256] <= 32'h66666666;
            reg_val_2_80002000[3][319:288] <= 32'hC0934C66;
            reg_val_2_80002000[3][351:320] <= 32'h9999999A;
            reg_val_2_80002000[3][383:352] <= 32'hBFF19999;
            reg_val_2_80002000[3][415:384] <= 32'h00000000;
            reg_val_2_80002000[3][447:416] <= 32'h00000000;
            reg_val_2_80002000[3][479:448] <= 32'hA3D70A3D;
            reg_val_2_80002000[3][511:480] <= 32'h40953A70;
            reg_val_2_80002000[4][31:0] <= 32'h53C8D4F1;
            reg_val_2_80002000[4][63:32] <= 32'h400921FB;
            reg_val_2_80002000[4][95:64] <= 32'hE2308C3A;
            reg_val_2_80002000[4][127:96] <= 32'h3E45798E;
            reg_val_2_80002000[4][159:128] <= 32'h00000000;
            reg_val_2_80002000[4][191:160] <= 32'h00000000;
            reg_val_2_80002000[4][223:192] <= 32'hA5C1FF09;
            reg_val_2_80002000[4][255:224] <= 32'h3E60DDC5;
            reg_val_2_80002000[4][287:256] <= 32'h00000000;
            reg_val_2_80002000[4][319:288] <= 32'h7FF00000;
            reg_val_2_80002000[4][351:320] <= 32'h00000000;
            reg_val_2_80002000[4][383:352] <= 32'h7FF00000;
            reg_val_2_80002000[4][415:384] <= 32'h00000000;
            reg_val_2_80002000[4][447:416] <= 32'h00000000;
            reg_val_2_80002000[4][479:448] <= 32'h00000000;
            reg_val_2_80002000[4][511:480] <= 32'h7FF80000;
            // fill-in reset values:
            reg_val_2_80002000[5][31:0] <= 32'h00000000;
            reg_val_2_80002000[5][63:32] <= 32'h00000000;
            reg_val_2_80002000[5][95:64] <= 32'h00000000;
            reg_val_2_80002000[5][127:96] <= 32'h00000000;
            reg_val_2_80002000[5][159:128] <= 32'h00000000;
            reg_val_2_80002000[5][191:160] <= 32'h00000000;
            reg_val_2_80002000[5][223:192] <= 32'h00000000;
            reg_val_2_80002000[5][255:224] <= 32'h00000000;
            reg_val_2_80002000[5][287:256] <= 32'h00000000;
            reg_val_2_80002000[5][319:288] <= 32'h00000000;
            reg_val_2_80002000[5][351:320] <= 32'h00000000;
            reg_val_2_80002000[5][383:352] <= 32'h00000000;
            reg_val_2_80002000[5][415:384] <= 32'h00000000;
            reg_val_2_80002000[5][447:416] <= 32'h00000000;
            reg_val_2_80002000[5][479:448] <= 32'h00000000;
            reg_val_2_80002000[5][511:480] <= 32'h00000000;
            reg_val_2_80002000[6][31:0] <= 32'h00000000;
            reg_val_2_80002000[6][63:32] <= 32'h00000000;
            reg_val_2_80002000[6][95:64] <= 32'h00000000;
            reg_val_2_80002000[6][127:96] <= 32'h00000000;
            reg_val_2_80002000[6][159:128] <= 32'h00000000;
            reg_val_2_80002000[6][191:160] <= 32'h00000000;
            reg_val_2_80002000[6][223:192] <= 32'h00000000;
            reg_val_2_80002000[6][255:224] <= 32'h00000000;
            reg_val_2_80002000[6][287:256] <= 32'h00000000;
            reg_val_2_80002000[6][319:288] <= 32'h00000000;
            reg_val_2_80002000[6][351:320] <= 32'h00000000;
            reg_val_2_80002000[6][383:352] <= 32'h00000000;
            reg_val_2_80002000[6][415:384] <= 32'h00000000;
            reg_val_2_80002000[6][447:416] <= 32'h00000000;
            reg_val_2_80002000[6][479:448] <= 32'h00000000;
            reg_val_2_80002000[6][511:480] <= 32'h00000000;
            reg_val_2_80002000[7][31:0] <= 32'h00000000;
            reg_val_2_80002000[7][63:32] <= 32'h00000000;
            reg_val_2_80002000[7][95:64] <= 32'h00000000;
            reg_val_2_80002000[7][127:96] <= 32'h00000000;
            reg_val_2_80002000[7][159:128] <= 32'h00000000;
            reg_val_2_80002000[7][191:160] <= 32'h00000000;
            reg_val_2_80002000[7][223:192] <= 32'h00000000;
            reg_val_2_80002000[7][255:224] <= 32'h00000000;
            reg_val_2_80002000[7][287:256] <= 32'h00000000;
            reg_val_2_80002000[7][319:288] <= 32'h00000000;
            reg_val_2_80002000[7][351:320] <= 32'h00000000;
            reg_val_2_80002000[7][383:352] <= 32'h00000000;
            reg_val_2_80002000[7][415:384] <= 32'h00000000;
            reg_val_2_80002000[7][447:416] <= 32'h00000000;
            reg_val_2_80002000[7][479:448] <= 32'h00000000;
            reg_val_2_80002000[7][511:480] <= 32'h00000000;
        end
        else
        begin
            reg_val_2_80002000 <= next_reg_val_2_80002000;
        end
    end
    
    always_comb begin : WRITE_LOGIC_2_80002000
        // hold reg val by default
        for (int i = 0; i < 8; i++)
        begin
            next_reg_val_2_80002000[i] = reg_val_2_80002000[i];
        end
        // update reg val if wen
        if (wen_2_80002000)
        begin
            // check for this byte enabled
            if (mem_req_byteen[0])  next_reg_val_2_80002000[wsel_2_80002000][7:0] = wdata_2_80002000[7:0];
            if (mem_req_byteen[1])  next_reg_val_2_80002000[wsel_2_80002000][15:8] = wdata_2_80002000[15:8];
            if (mem_req_byteen[2])  next_reg_val_2_80002000[wsel_2_80002000][23:16] = wdata_2_80002000[23:16];
            if (mem_req_byteen[3])  next_reg_val_2_80002000[wsel_2_80002000][31:24] = wdata_2_80002000[31:24];
            if (mem_req_byteen[4])  next_reg_val_2_80002000[wsel_2_80002000][39:32] = wdata_2_80002000[39:32];
            if (mem_req_byteen[5])  next_reg_val_2_80002000[wsel_2_80002000][47:40] = wdata_2_80002000[47:40];
            if (mem_req_byteen[6])  next_reg_val_2_80002000[wsel_2_80002000][55:48] = wdata_2_80002000[55:48];
            if (mem_req_byteen[7])  next_reg_val_2_80002000[wsel_2_80002000][63:56] = wdata_2_80002000[63:56];
            if (mem_req_byteen[8])  next_reg_val_2_80002000[wsel_2_80002000][71:64] = wdata_2_80002000[71:64];
            if (mem_req_byteen[9])  next_reg_val_2_80002000[wsel_2_80002000][79:72] = wdata_2_80002000[79:72];
            if (mem_req_byteen[10])  next_reg_val_2_80002000[wsel_2_80002000][87:80] = wdata_2_80002000[87:80];
            if (mem_req_byteen[11])  next_reg_val_2_80002000[wsel_2_80002000][95:88] = wdata_2_80002000[95:88];
            if (mem_req_byteen[12])  next_reg_val_2_80002000[wsel_2_80002000][103:96] = wdata_2_80002000[103:96];
            if (mem_req_byteen[13])  next_reg_val_2_80002000[wsel_2_80002000][111:104] = wdata_2_80002000[111:104];
            if (mem_req_byteen[14])  next_reg_val_2_80002000[wsel_2_80002000][119:112] = wdata_2_80002000[119:112];
            if (mem_req_byteen[15])  next_reg_val_2_80002000[wsel_2_80002000][127:120] = wdata_2_80002000[127:120];
            if (mem_req_byteen[16])  next_reg_val_2_80002000[wsel_2_80002000][135:128] = wdata_2_80002000[135:128];
            if (mem_req_byteen[17])  next_reg_val_2_80002000[wsel_2_80002000][143:136] = wdata_2_80002000[143:136];
            if (mem_req_byteen[18])  next_reg_val_2_80002000[wsel_2_80002000][151:144] = wdata_2_80002000[151:144];
            if (mem_req_byteen[19])  next_reg_val_2_80002000[wsel_2_80002000][159:152] = wdata_2_80002000[159:152];
            if (mem_req_byteen[20])  next_reg_val_2_80002000[wsel_2_80002000][167:160] = wdata_2_80002000[167:160];
            if (mem_req_byteen[21])  next_reg_val_2_80002000[wsel_2_80002000][175:168] = wdata_2_80002000[175:168];
            if (mem_req_byteen[22])  next_reg_val_2_80002000[wsel_2_80002000][183:176] = wdata_2_80002000[183:176];
            if (mem_req_byteen[23])  next_reg_val_2_80002000[wsel_2_80002000][191:184] = wdata_2_80002000[191:184];
            if (mem_req_byteen[24])  next_reg_val_2_80002000[wsel_2_80002000][199:192] = wdata_2_80002000[199:192];
            if (mem_req_byteen[25])  next_reg_val_2_80002000[wsel_2_80002000][207:200] = wdata_2_80002000[207:200];
            if (mem_req_byteen[26])  next_reg_val_2_80002000[wsel_2_80002000][215:208] = wdata_2_80002000[215:208];
            if (mem_req_byteen[27])  next_reg_val_2_80002000[wsel_2_80002000][223:216] = wdata_2_80002000[223:216];
            if (mem_req_byteen[28])  next_reg_val_2_80002000[wsel_2_80002000][231:224] = wdata_2_80002000[231:224];
            if (mem_req_byteen[29])  next_reg_val_2_80002000[wsel_2_80002000][239:232] = wdata_2_80002000[239:232];
            if (mem_req_byteen[30])  next_reg_val_2_80002000[wsel_2_80002000][247:240] = wdata_2_80002000[247:240];
            if (mem_req_byteen[31])  next_reg_val_2_80002000[wsel_2_80002000][255:248] = wdata_2_80002000[255:248];
            if (mem_req_byteen[32])  next_reg_val_2_80002000[wsel_2_80002000][263:256] = wdata_2_80002000[263:256];
            if (mem_req_byteen[33])  next_reg_val_2_80002000[wsel_2_80002000][271:264] = wdata_2_80002000[271:264];
            if (mem_req_byteen[34])  next_reg_val_2_80002000[wsel_2_80002000][279:272] = wdata_2_80002000[279:272];
            if (mem_req_byteen[35])  next_reg_val_2_80002000[wsel_2_80002000][287:280] = wdata_2_80002000[287:280];
            if (mem_req_byteen[36])  next_reg_val_2_80002000[wsel_2_80002000][295:288] = wdata_2_80002000[295:288];
            if (mem_req_byteen[37])  next_reg_val_2_80002000[wsel_2_80002000][303:296] = wdata_2_80002000[303:296];
            if (mem_req_byteen[38])  next_reg_val_2_80002000[wsel_2_80002000][311:304] = wdata_2_80002000[311:304];
            if (mem_req_byteen[39])  next_reg_val_2_80002000[wsel_2_80002000][319:312] = wdata_2_80002000[319:312];
            if (mem_req_byteen[40])  next_reg_val_2_80002000[wsel_2_80002000][327:320] = wdata_2_80002000[327:320];
            if (mem_req_byteen[41])  next_reg_val_2_80002000[wsel_2_80002000][335:328] = wdata_2_80002000[335:328];
            if (mem_req_byteen[42])  next_reg_val_2_80002000[wsel_2_80002000][343:336] = wdata_2_80002000[343:336];
            if (mem_req_byteen[43])  next_reg_val_2_80002000[wsel_2_80002000][351:344] = wdata_2_80002000[351:344];
            if (mem_req_byteen[44])  next_reg_val_2_80002000[wsel_2_80002000][359:352] = wdata_2_80002000[359:352];
            if (mem_req_byteen[45])  next_reg_val_2_80002000[wsel_2_80002000][367:360] = wdata_2_80002000[367:360];
            if (mem_req_byteen[46])  next_reg_val_2_80002000[wsel_2_80002000][375:368] = wdata_2_80002000[375:368];
            if (mem_req_byteen[47])  next_reg_val_2_80002000[wsel_2_80002000][383:376] = wdata_2_80002000[383:376];
            if (mem_req_byteen[48])  next_reg_val_2_80002000[wsel_2_80002000][391:384] = wdata_2_80002000[391:384];
            if (mem_req_byteen[49])  next_reg_val_2_80002000[wsel_2_80002000][399:392] = wdata_2_80002000[399:392];
            if (mem_req_byteen[50])  next_reg_val_2_80002000[wsel_2_80002000][407:400] = wdata_2_80002000[407:400];
            if (mem_req_byteen[51])  next_reg_val_2_80002000[wsel_2_80002000][415:408] = wdata_2_80002000[415:408];
            if (mem_req_byteen[52])  next_reg_val_2_80002000[wsel_2_80002000][423:416] = wdata_2_80002000[423:416];
            if (mem_req_byteen[53])  next_reg_val_2_80002000[wsel_2_80002000][431:424] = wdata_2_80002000[431:424];
            if (mem_req_byteen[54])  next_reg_val_2_80002000[wsel_2_80002000][439:432] = wdata_2_80002000[439:432];
            if (mem_req_byteen[55])  next_reg_val_2_80002000[wsel_2_80002000][447:440] = wdata_2_80002000[447:440];
            if (mem_req_byteen[56])  next_reg_val_2_80002000[wsel_2_80002000][455:448] = wdata_2_80002000[455:448];
            if (mem_req_byteen[57])  next_reg_val_2_80002000[wsel_2_80002000][463:456] = wdata_2_80002000[463:456];
            if (mem_req_byteen[58])  next_reg_val_2_80002000[wsel_2_80002000][471:464] = wdata_2_80002000[471:464];
            if (mem_req_byteen[59])  next_reg_val_2_80002000[wsel_2_80002000][479:472] = wdata_2_80002000[479:472];
            if (mem_req_byteen[60])  next_reg_val_2_80002000[wsel_2_80002000][487:480] = wdata_2_80002000[487:480];
            if (mem_req_byteen[61])  next_reg_val_2_80002000[wsel_2_80002000][495:488] = wdata_2_80002000[495:488];
            if (mem_req_byteen[62])  next_reg_val_2_80002000[wsel_2_80002000][503:496] = wdata_2_80002000[503:496];
            if (mem_req_byteen[63])  next_reg_val_2_80002000[wsel_2_80002000][511:504] = wdata_2_80002000[511:504];
        end
    end
    
    always_comb begin : READ_LOGIC_2_80002000
        // read val at rsel
        // multi block version (need select line)
        rdata_2_80002000 = reg_val_2_80002000[rsel_2_80002000];
    end
    
    // need reg file/chunk selection signal
    logic [2-1:0] chunk_sel;

    // addr hashing logic
    always_comb begin : ADDR_HASHING_LOGIC
        // default as address not out of bounds
        tb_addr_out_of_bounds = 1'b0;
        
        // bad address assertion:
        assert (
            (26'b10000000000000000000000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000000000000 + 32) ||
            (26'b10000000000000000001000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000001000000 + 2) ||
            (26'b10000000000000000010000000 <= mem_req_addr && mem_req_addr < 26'b10000000000000000010000000 + 8)
        ) else begin
            $display("mem request at address 0x%h = 0b%b not available in chunks", mem_req_addr, mem_req_addr);
            tb_addr_out_of_bounds = 1'b1;
        end
        
        // bit = 1 branch
        if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 19] == 1'b1)
        begin
            // select chunk @ 0x80002000
            chunk_sel = 2;
        end
        // bit = 0 branch
        else if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 19] == 1'b0)
        begin
            if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 20] == 1'b0)
            begin
                // select chunk @ 0x80000000
                chunk_sel = 0;
            end
            else if (mem_req_addr[`VX_MEM_ADDR_WIDTH - 20] == 1'b1)
            begin
                // select chunk @ 0x80001000
                chunk_sel = 1;
            end
        end
        else
        begin
            $display("error: got to else in high-level branch");
            tb_addr_out_of_bounds = 1'b1;
        end
        
        // hardlogicd outputs:
        
        // hardwiring for chunk 0 with multiple blocks
        wsel_0_80000000 = mem_req_addr[5-1 : 0];
        wdata_0_80000000 = mem_req_data;
        rsel_0_80000000 = mem_req_addr[5-1 : 0];
        
        // hardwiring for chunk 1 with multiple blocks
        wsel_1_80001000 = mem_req_addr[1-1 : 0];
        wdata_1_80001000 = mem_req_data;
        rsel_1_80001000 = mem_req_addr[1-1 : 0];
        
        // hardwiring for chunk 2 with multiple blocks
        wsel_2_80002000 = mem_req_addr[3-1 : 0];
        wdata_2_80002000 = mem_req_data;
        rsel_2_80002000 = mem_req_addr[3-1 : 0];
        
        // default outputs:
        mem_rsp_data = {16{32'hdeadbeef}};
        // chunk wen's:
        wen_0_80000000 = 1'b0;
        wen_1_80001000 = 1'b0;
        wen_2_80002000 = 1'b0;
        
        // case for routing to diff reg file chunks
        casez (chunk_sel)
        
            // select chunk 0 @ 0x80000000
            0:
            begin
                // write routing
                wen_0_80000000 = mem_req_rw & mem_req_valid;
                // read routing
                mem_rsp_data = rdata_0_80000000;
            end
        
            // select chunk 1 @ 0x80001000
            1:
            begin
                // write routing
                wen_1_80001000 = mem_req_rw & mem_req_valid;
                // read routing
                mem_rsp_data = rdata_1_80001000;
            end
        
            // select chunk 2 @ 0x80002000
            2:
            begin
                // write routing
                wen_2_80002000 = mem_req_rw & mem_req_valid;
                // read routing
                mem_rsp_data = rdata_2_80002000;
            end
        
            // shouldn't get here
            default:
            begin
                $display("error: got to default in chunk_sel case");
                mem_rsp_data = {16{32'hdeadbeef}};
                tb_addr_out_of_bounds = 1'b1;
            end
        endcase
    end

    // other combinational logic for memory interface
    always_comb begin : OTHER_MEM_COMB_LOGIC

        // mem_req_ready = 1'b1;           // always ready for request
        mem_rsp_valid = mem_req_valid;  // read ready immediately
            // update to buffer to later clock cycle
                // along with data read value

        mem_rsp_tag = mem_req_tag;      // match req immediately
    end

    // delayed mem_req_ready signals
    parameter MEM_REQ_READY_DELAY = 0;
    logic [MEM_REQ_READY_DELAY-1:0] mem_req_ready_reg, next_mem_req_ready_reg; 

    // delayed mem_req_ready reg logic
    always_ff @ (posedge clk) begin : MEM_REQ_READY_REG_LOGIC
    
        if (reset)
        begin
            mem_req_ready_reg = '0;
        end
        else
        begin
            mem_req_ready_reg = next_mem_req_ready_reg;
        end
    end

    // delayed mem_req_ready delay next state logic
    always_comb begin : MEM_REQ_READY_DELAY_NEXT_STATE_LOGIC

        next_mem_req_ready_reg = {mem_req_ready_reg[MEM_REQ_READY_DELAY-2:0], 1'b1};    // shift 1 left
        mem_req_ready = mem_req_ready_reg[MEM_REQ_READY_DELAY-1];                       // msb of shifter
    end

    // NOTES:
    // don't know what to do with: 
        // busy

endmodule

